magic
tech sky130A
magscale 1 2
timestamp 1647889164
<< viali >>
rect 9965 37417 9999 37451
rect 37841 37417 37875 37451
rect 49065 37417 49099 37451
rect 12357 37349 12391 37383
rect 23857 37349 23891 37383
rect 4445 37281 4479 37315
rect 9321 37281 9355 37315
rect 11897 37281 11931 37315
rect 14289 37281 14323 37315
rect 16129 37281 16163 37315
rect 28733 37281 28767 37315
rect 29929 37281 29963 37315
rect 30665 37281 30699 37315
rect 43269 37281 43303 37315
rect 48053 37281 48087 37315
rect 52193 37281 52227 37315
rect 1685 37213 1719 37247
rect 2421 37213 2455 37247
rect 2881 37213 2915 37247
rect 4261 37213 4295 37247
rect 6377 37213 6411 37247
rect 7389 37213 7423 37247
rect 7849 37213 7883 37247
rect 9873 37213 9907 37247
rect 12541 37213 12575 37247
rect 14565 37213 14599 37247
rect 16681 37213 16715 37247
rect 18429 37213 18463 37247
rect 19625 37213 19659 37247
rect 20177 37213 20211 37247
rect 24409 37213 24443 37247
rect 25421 37213 25455 37247
rect 25881 37213 25915 37247
rect 27997 37213 28031 37247
rect 28549 37213 28583 37247
rect 30481 37213 30515 37247
rect 32597 37213 32631 37247
rect 33517 37213 33551 37247
rect 33977 37213 34011 37247
rect 35909 37213 35943 37247
rect 37749 37213 37783 37247
rect 39037 37213 39071 37247
rect 39129 37213 39163 37247
rect 40141 37213 40175 37247
rect 40877 37213 40911 37247
rect 41705 37213 41739 37247
rect 42625 37213 42659 37247
rect 42717 37213 42751 37247
rect 46489 37213 46523 37247
rect 48973 37213 49007 37247
rect 50629 37213 50663 37247
rect 52745 37213 52779 37247
rect 54217 37213 54251 37247
rect 55689 37213 55723 37247
rect 56241 37213 56275 37247
rect 57897 37213 57931 37247
rect 20545 37145 20579 37179
rect 22385 37145 22419 37179
rect 22937 37145 22971 37179
rect 34805 37145 34839 37179
rect 34989 37145 35023 37179
rect 35633 37145 35667 37179
rect 36093 37145 36127 37179
rect 46213 37145 46247 37179
rect 46673 37145 46707 37179
rect 48329 37145 48363 37179
rect 56701 37145 56735 37179
rect 1501 37077 1535 37111
rect 2237 37077 2271 37111
rect 6561 37077 6595 37111
rect 8033 37077 8067 37111
rect 16865 37077 16899 37111
rect 18245 37077 18279 37111
rect 22293 37077 22327 37111
rect 24593 37077 24627 37111
rect 26065 37077 26099 37111
rect 32413 37077 32447 37111
rect 34161 37077 34195 37111
rect 35173 37077 35207 37111
rect 35725 37077 35759 37111
rect 38853 37077 38887 37111
rect 39957 37077 39991 37111
rect 40693 37077 40727 37111
rect 41889 37077 41923 37111
rect 42441 37077 42475 37111
rect 46305 37077 46339 37111
rect 50721 37077 50755 37111
rect 52929 37077 52963 37111
rect 54401 37077 54435 37111
rect 58081 37077 58115 37111
rect 1501 36873 1535 36907
rect 3985 36873 4019 36907
rect 26341 36873 26375 36907
rect 37473 36873 37507 36907
rect 47593 36873 47627 36907
rect 48421 36873 48455 36907
rect 48973 36873 49007 36907
rect 50353 36873 50387 36907
rect 57345 36873 57379 36907
rect 8493 36805 8527 36839
rect 14197 36805 14231 36839
rect 20821 36805 20855 36839
rect 28089 36805 28123 36839
rect 38393 36805 38427 36839
rect 41797 36805 41831 36839
rect 43913 36805 43947 36839
rect 56793 36805 56827 36839
rect 58081 36805 58115 36839
rect 1685 36737 1719 36771
rect 5457 36737 5491 36771
rect 7481 36737 7515 36771
rect 8309 36737 8343 36771
rect 8585 36737 8619 36771
rect 9045 36737 9079 36771
rect 20177 36737 20211 36771
rect 22477 36737 22511 36771
rect 24133 36737 24167 36771
rect 24961 36737 24995 36771
rect 26157 36737 26191 36771
rect 28733 36737 28767 36771
rect 32321 36737 32355 36771
rect 34713 36737 34747 36771
rect 34897 36737 34931 36771
rect 35541 36737 35575 36771
rect 38301 36737 38335 36771
rect 38577 36737 38611 36771
rect 39313 36737 39347 36771
rect 40325 36737 40359 36771
rect 40509 36737 40543 36771
rect 41613 36737 41647 36771
rect 41889 36737 41923 36771
rect 42533 36737 42567 36771
rect 43545 36737 43579 36771
rect 43729 36737 43763 36771
rect 46121 36737 46155 36771
rect 46581 36737 46615 36771
rect 47777 36737 47811 36771
rect 5549 36669 5583 36703
rect 5825 36669 5859 36703
rect 7113 36669 7147 36703
rect 7573 36669 7607 36703
rect 8125 36669 8159 36703
rect 19901 36669 19935 36703
rect 22385 36669 22419 36703
rect 24041 36669 24075 36703
rect 25697 36669 25731 36703
rect 26065 36669 26099 36703
rect 27261 36669 27295 36703
rect 28641 36669 28675 36703
rect 32413 36669 32447 36703
rect 47961 36669 47995 36703
rect 22845 36601 22879 36635
rect 40693 36601 40727 36635
rect 57897 36601 57931 36635
rect 6469 36533 6503 36567
rect 29101 36533 29135 36567
rect 30205 36533 30239 36567
rect 32689 36533 32723 36567
rect 35081 36533 35115 36567
rect 35817 36533 35851 36567
rect 36001 36533 36035 36567
rect 38761 36533 38795 36567
rect 39405 36533 39439 36567
rect 39773 36533 39807 36567
rect 41429 36533 41463 36567
rect 42625 36533 42659 36567
rect 42993 36533 43027 36567
rect 8953 36329 8987 36363
rect 19441 36329 19475 36363
rect 21741 36329 21775 36363
rect 23857 36329 23891 36363
rect 24409 36329 24443 36363
rect 24777 36329 24811 36363
rect 26433 36329 26467 36363
rect 28641 36329 28675 36363
rect 31585 36329 31619 36363
rect 33425 36329 33459 36363
rect 38485 36329 38519 36363
rect 48697 36329 48731 36363
rect 7113 36261 7147 36295
rect 32781 36261 32815 36295
rect 9321 36193 9355 36227
rect 19717 36193 19751 36227
rect 22201 36193 22235 36227
rect 30757 36193 30791 36227
rect 32505 36193 32539 36227
rect 38117 36193 38151 36227
rect 41429 36193 41463 36227
rect 49065 36193 49099 36227
rect 1685 36125 1719 36159
rect 8217 36125 8251 36159
rect 8401 36125 8435 36159
rect 9137 36125 9171 36159
rect 9781 36125 9815 36159
rect 19257 36125 19291 36159
rect 19441 36125 19475 36159
rect 21281 36125 21315 36159
rect 21373 36125 21407 36159
rect 21557 36125 21591 36159
rect 22385 36125 22419 36159
rect 23673 36125 23707 36159
rect 23857 36125 23891 36159
rect 24409 36125 24443 36159
rect 24501 36125 24535 36159
rect 26249 36125 26283 36159
rect 26433 36125 26467 36159
rect 28457 36125 28491 36159
rect 28641 36125 28675 36159
rect 29561 36125 29595 36159
rect 29837 36125 29871 36159
rect 30665 36125 30699 36159
rect 30849 36125 30883 36159
rect 31309 36125 31343 36159
rect 32413 36125 32447 36159
rect 36461 36125 36495 36159
rect 37197 36125 37231 36159
rect 38209 36125 38243 36159
rect 39957 36125 39991 36159
rect 40325 36125 40359 36159
rect 42625 36125 42659 36159
rect 42993 36125 43027 36159
rect 47133 36125 47167 36159
rect 47685 36125 47719 36159
rect 48973 36125 49007 36159
rect 58173 36125 58207 36159
rect 7757 36057 7791 36091
rect 22569 36057 22603 36091
rect 30021 36057 30055 36091
rect 33609 36057 33643 36091
rect 35541 36057 35575 36091
rect 44465 36057 44499 36091
rect 57897 36057 57931 36091
rect 1501 35989 1535 36023
rect 8309 35989 8343 36023
rect 29653 35989 29687 36023
rect 31769 35989 31803 36023
rect 33241 35989 33275 36023
rect 33409 35989 33443 36023
rect 39129 35989 39163 36023
rect 6653 35785 6687 35819
rect 6745 35785 6779 35819
rect 8861 35785 8895 35819
rect 28483 35785 28517 35819
rect 29101 35785 29135 35819
rect 32781 35785 32815 35819
rect 40141 35785 40175 35819
rect 46121 35785 46155 35819
rect 49249 35785 49283 35819
rect 58173 35785 58207 35819
rect 6561 35717 6595 35751
rect 8033 35717 8067 35751
rect 9965 35717 9999 35751
rect 19165 35717 19199 35751
rect 23213 35717 23247 35751
rect 23397 35717 23431 35751
rect 28273 35717 28307 35751
rect 6929 35649 6963 35683
rect 7941 35649 7975 35683
rect 8125 35649 8159 35683
rect 8309 35649 8343 35683
rect 8769 35649 8803 35683
rect 8953 35649 8987 35683
rect 11713 35649 11747 35683
rect 11897 35649 11931 35683
rect 18797 35649 18831 35683
rect 19625 35649 19659 35683
rect 19717 35649 19751 35683
rect 23029 35649 23063 35683
rect 29469 35649 29503 35683
rect 32321 35649 32355 35683
rect 32505 35649 32539 35683
rect 32873 35649 32907 35683
rect 45293 35649 45327 35683
rect 49249 35649 49283 35683
rect 49433 35649 49467 35683
rect 18705 35581 18739 35615
rect 29377 35581 29411 35615
rect 45201 35581 45235 35615
rect 6377 35513 6411 35547
rect 11989 35513 12023 35547
rect 19073 35513 19107 35547
rect 19993 35513 20027 35547
rect 28641 35513 28675 35547
rect 7757 35445 7791 35479
rect 9413 35445 9447 35479
rect 12541 35445 12575 35479
rect 19809 35445 19843 35479
rect 28457 35445 28491 35479
rect 30205 35445 30239 35479
rect 41061 35445 41095 35479
rect 6745 35241 6779 35275
rect 7757 35241 7791 35275
rect 9045 35241 9079 35275
rect 9597 35241 9631 35275
rect 11713 35241 11747 35275
rect 16589 35241 16623 35275
rect 18521 35241 18555 35275
rect 18705 35241 18739 35275
rect 22293 35241 22327 35275
rect 25237 35241 25271 35275
rect 28641 35241 28675 35275
rect 37473 35241 37507 35275
rect 43637 35241 43671 35275
rect 22385 35173 22419 35207
rect 34713 35173 34747 35207
rect 53573 35173 53607 35207
rect 7021 35105 7055 35139
rect 8217 35105 8251 35139
rect 10885 35105 10919 35139
rect 11345 35105 11379 35139
rect 35173 35105 35207 35139
rect 37565 35105 37599 35139
rect 43269 35105 43303 35139
rect 47593 35105 47627 35139
rect 53113 35105 53147 35139
rect 57897 35105 57931 35139
rect 7113 35037 7147 35071
rect 7941 35037 7975 35071
rect 8125 35037 8159 35071
rect 11529 35037 11563 35071
rect 12173 35037 12207 35071
rect 12541 35037 12575 35071
rect 12725 35037 12759 35071
rect 13277 35037 13311 35071
rect 16037 35037 16071 35071
rect 17141 35037 17175 35071
rect 21097 35037 21131 35071
rect 21557 35037 21591 35071
rect 23489 35037 23523 35071
rect 23673 35037 23707 35071
rect 25145 35037 25179 35071
rect 25421 35037 25455 35071
rect 25605 35037 25639 35071
rect 28365 35037 28399 35071
rect 28641 35037 28675 35071
rect 35081 35037 35115 35071
rect 37473 35037 37507 35071
rect 43361 35037 43395 35071
rect 48605 35037 48639 35071
rect 49157 35037 49191 35071
rect 49341 35037 49375 35071
rect 53205 35037 53239 35071
rect 58173 35037 58207 35071
rect 15669 34969 15703 35003
rect 15853 34969 15887 35003
rect 18337 34969 18371 35003
rect 20729 34969 20763 35003
rect 22753 34969 22787 35003
rect 23857 34969 23891 35003
rect 50169 34969 50203 35003
rect 12541 34901 12575 34935
rect 18537 34901 18571 34935
rect 28457 34901 28491 34935
rect 37841 34901 37875 34935
rect 49341 34901 49375 34935
rect 8493 34697 8527 34731
rect 16865 34697 16899 34731
rect 18251 34697 18285 34731
rect 20269 34697 20303 34731
rect 21097 34697 21131 34731
rect 48789 34697 48823 34731
rect 52193 34697 52227 34731
rect 53573 34697 53607 34731
rect 58173 34697 58207 34731
rect 10793 34629 10827 34663
rect 11713 34629 11747 34663
rect 20729 34629 20763 34663
rect 20945 34629 20979 34663
rect 25053 34629 25087 34663
rect 27905 34629 27939 34663
rect 35173 34629 35207 34663
rect 35357 34629 35391 34663
rect 39129 34629 39163 34663
rect 53021 34629 53055 34663
rect 54125 34629 54159 34663
rect 7849 34561 7883 34595
rect 8033 34561 8067 34595
rect 10609 34561 10643 34595
rect 12357 34561 12391 34595
rect 12725 34561 12759 34595
rect 15485 34561 15519 34595
rect 16681 34561 16715 34595
rect 16865 34561 16899 34595
rect 18153 34561 18187 34595
rect 18337 34561 18371 34595
rect 18429 34561 18463 34595
rect 20085 34561 20119 34595
rect 20269 34561 20303 34595
rect 24961 34561 24995 34595
rect 25237 34561 25271 34595
rect 25421 34561 25455 34595
rect 27721 34561 27755 34595
rect 27997 34561 28031 34595
rect 32413 34561 32447 34595
rect 32781 34561 32815 34595
rect 34989 34561 35023 34595
rect 35817 34561 35851 34595
rect 36001 34561 36035 34595
rect 37841 34561 37875 34595
rect 38669 34561 38703 34595
rect 38945 34561 38979 34595
rect 40049 34561 40083 34595
rect 42993 34561 43027 34595
rect 43177 34561 43211 34595
rect 48513 34561 48547 34595
rect 49709 34561 49743 34595
rect 49985 34561 50019 34595
rect 50353 34561 50387 34595
rect 52009 34561 52043 34595
rect 52193 34561 52227 34595
rect 52745 34561 52779 34595
rect 52837 34561 52871 34595
rect 53481 34561 53515 34595
rect 53665 34561 53699 34595
rect 7205 34493 7239 34527
rect 9045 34493 9079 34527
rect 10977 34493 11011 34527
rect 15209 34493 15243 34527
rect 16129 34493 16163 34527
rect 27261 34493 27295 34527
rect 37933 34493 37967 34527
rect 39681 34493 39715 34527
rect 40141 34493 40175 34527
rect 48789 34493 48823 34527
rect 49433 34493 49467 34527
rect 11529 34425 11563 34459
rect 27997 34425 28031 34459
rect 33609 34425 33643 34459
rect 35909 34425 35943 34459
rect 38761 34425 38795 34459
rect 43177 34425 43211 34459
rect 48605 34425 48639 34459
rect 50721 34425 50755 34459
rect 53021 34425 53055 34459
rect 7665 34357 7699 34391
rect 14197 34357 14231 34391
rect 20913 34357 20947 34391
rect 28457 34357 28491 34391
rect 38117 34357 38151 34391
rect 10885 34153 10919 34187
rect 15209 34153 15243 34187
rect 16037 34153 16071 34187
rect 19257 34153 19291 34187
rect 25145 34153 25179 34187
rect 27905 34153 27939 34187
rect 28549 34153 28583 34187
rect 32781 34153 32815 34187
rect 33149 34153 33183 34187
rect 38393 34153 38427 34187
rect 40049 34153 40083 34187
rect 43821 34153 43855 34187
rect 48697 34153 48731 34187
rect 49525 34153 49559 34187
rect 24961 34085 24995 34119
rect 28917 34085 28951 34119
rect 38301 34085 38335 34119
rect 42257 34085 42291 34119
rect 44189 34085 44223 34119
rect 50721 34085 50755 34119
rect 11529 34017 11563 34051
rect 11713 34017 11747 34051
rect 22661 34017 22695 34051
rect 23397 34017 23431 34051
rect 32229 34017 32263 34051
rect 35909 34017 35943 34051
rect 37289 34017 37323 34051
rect 37933 34017 37967 34051
rect 41797 34017 41831 34051
rect 43913 34017 43947 34051
rect 53481 34017 53515 34051
rect 8125 33949 8159 33983
rect 8401 33949 8435 33983
rect 9321 33949 9355 33983
rect 10885 33949 10919 33983
rect 11069 33949 11103 33983
rect 12449 33949 12483 33983
rect 12633 33949 12667 33983
rect 12909 33949 12943 33983
rect 15025 33949 15059 33983
rect 15209 33949 15243 33983
rect 15669 33949 15703 33983
rect 15853 33949 15887 33983
rect 18429 33949 18463 33983
rect 18705 33949 18739 33983
rect 19441 33949 19475 33983
rect 19717 33949 19751 33983
rect 23213 33949 23247 33983
rect 28549 33949 28583 33983
rect 28641 33949 28675 33983
rect 31217 33949 31251 33983
rect 31401 33949 31435 33983
rect 32689 33949 32723 33983
rect 37197 33949 37231 33983
rect 37381 33949 37415 33983
rect 39957 33949 39991 33983
rect 40141 33949 40175 33983
rect 40785 33949 40819 33983
rect 40969 33949 41003 33983
rect 41889 33949 41923 33983
rect 42901 33949 42935 33983
rect 42993 33949 43027 33983
rect 43177 33949 43211 33983
rect 43821 33949 43855 33983
rect 45017 33949 45051 33983
rect 45109 33949 45143 33983
rect 45293 33949 45327 33983
rect 49433 33949 49467 33983
rect 51273 33949 51307 33983
rect 51549 33949 51583 33983
rect 52193 33949 52227 33983
rect 52561 33949 52595 33983
rect 52929 33949 52963 33983
rect 9505 33881 9539 33915
rect 12081 33881 12115 33915
rect 18521 33881 18555 33915
rect 24685 33881 24719 33915
rect 27721 33881 27755 33915
rect 27921 33881 27955 33915
rect 35357 33881 35391 33915
rect 40877 33881 40911 33915
rect 49249 33881 49283 33915
rect 51733 33881 51767 33915
rect 53573 33881 53607 33915
rect 18429 33813 18463 33847
rect 19625 33813 19659 33847
rect 28089 33813 28123 33847
rect 43361 33813 43395 33847
rect 45477 33813 45511 33847
rect 51365 33813 51399 33847
rect 11805 33609 11839 33643
rect 17969 33609 18003 33643
rect 27629 33609 27663 33643
rect 31033 33609 31067 33643
rect 57989 33609 58023 33643
rect 8493 33541 8527 33575
rect 9137 33541 9171 33575
rect 9689 33541 9723 33575
rect 17141 33541 17175 33575
rect 23305 33541 23339 33575
rect 29101 33541 29135 33575
rect 42533 33541 42567 33575
rect 48421 33541 48455 33575
rect 52193 33541 52227 33575
rect 52745 33541 52779 33575
rect 52945 33541 52979 33575
rect 1869 33473 1903 33507
rect 6745 33473 6779 33507
rect 6929 33473 6963 33507
rect 7573 33473 7607 33507
rect 8401 33473 8435 33507
rect 8585 33473 8619 33507
rect 11989 33473 12023 33507
rect 23029 33473 23063 33507
rect 23213 33473 23247 33507
rect 24869 33473 24903 33507
rect 27537 33473 27571 33507
rect 27813 33473 27847 33507
rect 28641 33473 28675 33507
rect 30941 33473 30975 33507
rect 31217 33473 31251 33507
rect 31401 33473 31435 33507
rect 35725 33473 35759 33507
rect 42441 33473 42475 33507
rect 42625 33473 42659 33507
rect 44649 33473 44683 33507
rect 44925 33473 44959 33507
rect 45109 33473 45143 33507
rect 45477 33473 45511 33507
rect 48973 33473 49007 33507
rect 49341 33473 49375 33507
rect 58173 33473 58207 33507
rect 7481 33405 7515 33439
rect 12173 33405 12207 33439
rect 17417 33405 17451 33439
rect 24961 33405 24995 33439
rect 27077 33405 27111 33439
rect 28549 33405 28583 33439
rect 36185 33405 36219 33439
rect 45385 33405 45419 33439
rect 47961 33405 47995 33439
rect 6653 33337 6687 33371
rect 7941 33337 7975 33371
rect 25237 33337 25271 33371
rect 44741 33337 44775 33371
rect 53113 33337 53147 33371
rect 1961 33269 1995 33303
rect 22845 33269 22879 33303
rect 27813 33269 27847 33303
rect 35909 33269 35943 33303
rect 52929 33269 52963 33303
rect 1593 33065 1627 33099
rect 8953 33065 8987 33099
rect 18521 33065 18555 33099
rect 28089 33065 28123 33099
rect 28181 33065 28215 33099
rect 48881 33065 48915 33099
rect 58173 33065 58207 33099
rect 16681 32997 16715 33031
rect 19257 32997 19291 33031
rect 27537 32997 27571 33031
rect 38761 32997 38795 33031
rect 7665 32929 7699 32963
rect 19533 32929 19567 32963
rect 22845 32929 22879 32963
rect 26341 32929 26375 32963
rect 28273 32929 28307 32963
rect 30481 32929 30515 32963
rect 31309 32929 31343 32963
rect 35817 32929 35851 32963
rect 49433 32929 49467 32963
rect 7113 32861 7147 32895
rect 7297 32861 7331 32895
rect 8125 32861 8159 32895
rect 11621 32861 11655 32895
rect 11989 32861 12023 32895
rect 16497 32861 16531 32895
rect 16773 32861 16807 32895
rect 18429 32861 18463 32895
rect 18521 32861 18555 32895
rect 19625 32861 19659 32895
rect 22017 32861 22051 32895
rect 22293 32861 22327 32895
rect 26433 32861 26467 32895
rect 27261 32861 27295 32895
rect 27997 32861 28031 32895
rect 34805 32861 34839 32895
rect 35173 32861 35207 32895
rect 37933 32861 37967 32895
rect 45017 32861 45051 32895
rect 45201 32861 45235 32895
rect 45845 32861 45879 32895
rect 46213 32861 46247 32895
rect 48789 32861 48823 32895
rect 48973 32861 49007 32895
rect 18245 32793 18279 32827
rect 27537 32793 27571 32827
rect 38485 32793 38519 32827
rect 47685 32793 47719 32827
rect 7297 32725 7331 32759
rect 8309 32725 8343 32759
rect 12633 32725 12667 32759
rect 16313 32725 16347 32759
rect 17325 32725 17359 32759
rect 20361 32725 20395 32759
rect 26801 32725 26835 32759
rect 27353 32725 27387 32759
rect 38945 32725 38979 32759
rect 45109 32725 45143 32759
rect 38301 32521 38335 32555
rect 40049 32521 40083 32555
rect 45569 32521 45603 32555
rect 49525 32521 49559 32555
rect 9505 32453 9539 32487
rect 15301 32453 15335 32487
rect 18705 32453 18739 32487
rect 24409 32453 24443 32487
rect 24593 32453 24627 32487
rect 30573 32453 30607 32487
rect 33885 32453 33919 32487
rect 34621 32453 34655 32487
rect 7389 32385 7423 32419
rect 8125 32385 8159 32419
rect 10425 32385 10459 32419
rect 13277 32385 13311 32419
rect 13921 32385 13955 32419
rect 15209 32385 15243 32419
rect 15393 32385 15427 32419
rect 16681 32385 16715 32419
rect 18245 32385 18279 32419
rect 18337 32385 18371 32419
rect 18521 32385 18555 32419
rect 24225 32385 24259 32419
rect 30481 32385 30515 32419
rect 30665 32385 30699 32419
rect 33793 32385 33827 32419
rect 33977 32385 34011 32419
rect 34529 32385 34563 32419
rect 34805 32385 34839 32419
rect 37289 32385 37323 32419
rect 38209 32385 38243 32419
rect 38393 32385 38427 32419
rect 39037 32385 39071 32419
rect 39221 32385 39255 32419
rect 41337 32385 41371 32419
rect 43361 32385 43395 32419
rect 45293 32385 45327 32419
rect 45661 32385 45695 32419
rect 48697 32385 48731 32419
rect 49157 32385 49191 32419
rect 52929 32385 52963 32419
rect 9045 32317 9079 32351
rect 10701 32317 10735 32351
rect 17141 32317 17175 32351
rect 22017 32317 22051 32351
rect 22477 32317 22511 32351
rect 37473 32317 37507 32351
rect 41245 32317 41279 32351
rect 41705 32317 41739 32351
rect 43453 32317 43487 32351
rect 45109 32317 45143 32351
rect 53113 32317 53147 32351
rect 22293 32249 22327 32283
rect 34989 32249 35023 32283
rect 43729 32249 43763 32283
rect 10517 32181 10551 32215
rect 10609 32181 10643 32215
rect 14381 32181 14415 32215
rect 16773 32181 16807 32215
rect 17601 32181 17635 32215
rect 27077 32181 27111 32215
rect 27721 32181 27755 32215
rect 52745 32181 52779 32215
rect 2513 31977 2547 32011
rect 8401 31977 8435 32011
rect 9321 31977 9355 32011
rect 10609 31977 10643 32011
rect 13277 31977 13311 32011
rect 15669 31977 15703 32011
rect 16313 31977 16347 32011
rect 16497 31977 16531 32011
rect 17049 31977 17083 32011
rect 18429 31977 18463 32011
rect 22569 31977 22603 32011
rect 23305 31977 23339 32011
rect 26801 31977 26835 32011
rect 32597 31977 32631 32011
rect 34161 31977 34195 32011
rect 41797 31977 41831 32011
rect 47961 31977 47995 32011
rect 49065 31977 49099 32011
rect 10149 31909 10183 31943
rect 10977 31909 11011 31943
rect 20177 31909 20211 31943
rect 22753 31909 22787 31943
rect 32413 31909 32447 31943
rect 57897 31909 57931 31943
rect 9413 31841 9447 31875
rect 9873 31841 9907 31875
rect 10701 31841 10735 31875
rect 21833 31841 21867 31875
rect 24501 31841 24535 31875
rect 24961 31841 24995 31875
rect 30665 31841 30699 31875
rect 35725 31841 35759 31875
rect 38117 31841 38151 31875
rect 38669 31841 38703 31875
rect 39129 31841 39163 31875
rect 48605 31841 48639 31875
rect 2053 31773 2087 31807
rect 2697 31773 2731 31807
rect 3157 31773 3191 31807
rect 7113 31773 7147 31807
rect 7573 31773 7607 31807
rect 9137 31773 9171 31807
rect 10057 31773 10091 31807
rect 10149 31773 10183 31807
rect 10609 31773 10643 31807
rect 13553 31773 13587 31807
rect 15209 31773 15243 31807
rect 15485 31773 15519 31807
rect 17969 31773 18003 31807
rect 18245 31773 18279 31807
rect 20821 31773 20855 31807
rect 22293 31773 22327 31807
rect 24593 31773 24627 31807
rect 26985 31773 27019 31807
rect 27261 31773 27295 31807
rect 27445 31773 27479 31807
rect 29653 31773 29687 31807
rect 33977 31773 34011 31807
rect 34161 31773 34195 31807
rect 34805 31773 34839 31807
rect 38025 31773 38059 31807
rect 38209 31773 38243 31807
rect 39037 31773 39071 31807
rect 39313 31773 39347 31807
rect 41705 31773 41739 31807
rect 41889 31773 41923 31807
rect 45109 31773 45143 31807
rect 45569 31773 45603 31807
rect 45753 31773 45787 31807
rect 47869 31773 47903 31807
rect 48053 31773 48087 31807
rect 48697 31773 48731 31807
rect 52929 31773 52963 31807
rect 53297 31773 53331 31807
rect 55321 31773 55355 31807
rect 56333 31773 56367 31807
rect 57437 31773 57471 31807
rect 58081 31773 58115 31807
rect 1869 31705 1903 31739
rect 13277 31705 13311 31739
rect 15301 31705 15335 31739
rect 16129 31705 16163 31739
rect 16329 31705 16363 31739
rect 32137 31705 32171 31739
rect 45385 31705 45419 31739
rect 8953 31637 8987 31671
rect 13461 31637 13495 31671
rect 18061 31637 18095 31671
rect 29009 31637 29043 31671
rect 10057 31433 10091 31467
rect 13737 31433 13771 31467
rect 32597 31433 32631 31467
rect 37841 31433 37875 31467
rect 48881 31433 48915 31467
rect 49801 31433 49835 31467
rect 1593 31365 1627 31399
rect 7297 31365 7331 31399
rect 7665 31365 7699 31399
rect 13369 31365 13403 31399
rect 13569 31365 13603 31399
rect 22845 31365 22879 31399
rect 27077 31365 27111 31399
rect 32137 31365 32171 31399
rect 54953 31365 54987 31399
rect 7205 31297 7239 31331
rect 10149 31297 10183 31331
rect 18061 31297 18095 31331
rect 18245 31297 18279 31331
rect 18521 31297 18555 31331
rect 21833 31297 21867 31331
rect 22201 31297 22235 31331
rect 27537 31297 27571 31331
rect 28273 31297 28307 31331
rect 28641 31297 28675 31331
rect 29653 31297 29687 31331
rect 37473 31297 37507 31331
rect 40785 31297 40819 31331
rect 45477 31297 45511 31331
rect 45753 31297 45787 31331
rect 48421 31297 48455 31331
rect 48513 31297 48547 31331
rect 49341 31297 49375 31331
rect 51917 31297 51951 31331
rect 52101 31297 52135 31331
rect 52193 31297 52227 31331
rect 55413 31297 55447 31331
rect 7389 31229 7423 31263
rect 9781 31229 9815 31263
rect 18429 31229 18463 31263
rect 22109 31229 22143 31263
rect 27169 31229 27203 31263
rect 30113 31229 30147 31263
rect 37381 31229 37415 31263
rect 40693 31229 40727 31263
rect 41153 31229 41187 31263
rect 44465 31229 44499 31263
rect 48605 31229 48639 31263
rect 48697 31229 48731 31263
rect 55505 31229 55539 31263
rect 7849 31161 7883 31195
rect 22201 31161 22235 31195
rect 28089 31161 28123 31195
rect 32413 31161 32447 31195
rect 44833 31161 44867 31195
rect 44925 31161 44959 31195
rect 45569 31161 45603 31195
rect 45661 31161 45695 31195
rect 45937 31161 45971 31195
rect 9873 31093 9907 31127
rect 9965 31093 9999 31127
rect 13553 31093 13587 31127
rect 21189 31093 21223 31127
rect 28365 31093 28399 31127
rect 29101 31093 29135 31127
rect 29745 31093 29779 31127
rect 49433 31093 49467 31127
rect 51733 31093 51767 31127
rect 10057 30889 10091 30923
rect 13001 30889 13035 30923
rect 19349 30889 19383 30923
rect 22661 30889 22695 30923
rect 27813 30889 27847 30923
rect 37381 30889 37415 30923
rect 45109 30889 45143 30923
rect 45661 30889 45695 30923
rect 55505 30889 55539 30923
rect 10333 30821 10367 30855
rect 18061 30821 18095 30855
rect 30941 30821 30975 30855
rect 48973 30821 49007 30855
rect 18337 30753 18371 30787
rect 26893 30753 26927 30787
rect 30481 30753 30515 30787
rect 31401 30753 31435 30787
rect 45017 30753 45051 30787
rect 55321 30753 55355 30787
rect 7297 30685 7331 30719
rect 10241 30685 10275 30719
rect 10425 30685 10459 30719
rect 10517 30685 10551 30719
rect 13001 30685 13035 30719
rect 13093 30685 13127 30719
rect 14381 30685 14415 30719
rect 14565 30685 14599 30719
rect 17509 30685 17543 30719
rect 18429 30685 18463 30719
rect 22845 30685 22879 30719
rect 23121 30685 23155 30719
rect 26985 30685 27019 30719
rect 27997 30685 28031 30719
rect 28181 30685 28215 30719
rect 30573 30685 30607 30719
rect 37197 30685 37231 30719
rect 37381 30685 37415 30719
rect 45480 30685 45514 30719
rect 48329 30685 48363 30719
rect 48421 30685 48455 30719
rect 48605 30685 48639 30719
rect 48789 30685 48823 30719
rect 50905 30685 50939 30719
rect 52285 30685 52319 30719
rect 52745 30685 52779 30719
rect 55781 30685 55815 30719
rect 7389 30617 7423 30651
rect 16037 30617 16071 30651
rect 48697 30617 48731 30651
rect 51089 30617 51123 30651
rect 13369 30549 13403 30583
rect 19901 30549 19935 30583
rect 22201 30549 22235 30583
rect 23029 30549 23063 30583
rect 24501 30549 24535 30583
rect 27353 30549 27387 30583
rect 28733 30549 28767 30583
rect 45477 30549 45511 30583
rect 51273 30549 51307 30583
rect 55689 30549 55723 30583
rect 56241 30549 56275 30583
rect 23121 30345 23155 30379
rect 24501 30345 24535 30379
rect 27537 30345 27571 30379
rect 40141 30345 40175 30379
rect 44373 30345 44407 30379
rect 45109 30345 45143 30379
rect 48605 30345 48639 30379
rect 55965 30345 55999 30379
rect 7021 30277 7055 30311
rect 9597 30277 9631 30311
rect 13185 30277 13219 30311
rect 16681 30277 16715 30311
rect 22477 30277 22511 30311
rect 33701 30277 33735 30311
rect 42625 30277 42659 30311
rect 55137 30277 55171 30311
rect 6837 30209 6871 30243
rect 7481 30209 7515 30243
rect 7665 30209 7699 30243
rect 9873 30209 9907 30243
rect 12909 30209 12943 30243
rect 13001 30209 13035 30243
rect 15393 30209 15427 30243
rect 15577 30209 15611 30243
rect 15853 30209 15887 30243
rect 16129 30209 16163 30243
rect 16957 30209 16991 30243
rect 18429 30209 18463 30243
rect 19901 30209 19935 30243
rect 20729 30209 20763 30243
rect 23029 30209 23063 30243
rect 23213 30209 23247 30243
rect 24133 30209 24167 30243
rect 32873 30209 32907 30243
rect 35173 30209 35207 30243
rect 36001 30209 36035 30243
rect 37289 30209 37323 30243
rect 37565 30209 37599 30243
rect 37841 30209 37875 30243
rect 37933 30209 37967 30243
rect 39773 30209 39807 30243
rect 42441 30209 42475 30243
rect 42717 30209 42751 30243
rect 43177 30209 43211 30243
rect 43361 30209 43395 30243
rect 44281 30209 44315 30243
rect 44465 30209 44499 30243
rect 44925 30209 44959 30243
rect 45293 30209 45327 30243
rect 48145 30209 48179 30243
rect 51273 30209 51307 30243
rect 51641 30209 51675 30243
rect 52745 30209 52779 30243
rect 55321 30209 55355 30243
rect 55505 30209 55539 30243
rect 55965 30209 55999 30243
rect 56149 30209 56183 30243
rect 9781 30141 9815 30175
rect 9965 30141 9999 30175
rect 13185 30141 13219 30175
rect 16773 30141 16807 30175
rect 18705 30141 18739 30175
rect 19809 30141 19843 30175
rect 24225 30141 24259 30175
rect 32781 30141 32815 30175
rect 35081 30141 35115 30175
rect 36461 30141 36495 30175
rect 39681 30141 39715 30175
rect 41061 30141 41095 30175
rect 52101 30141 52135 30175
rect 16129 30073 16163 30107
rect 20269 30073 20303 30107
rect 30389 30073 30423 30107
rect 35541 30073 35575 30107
rect 37657 30073 37691 30107
rect 40693 30073 40727 30107
rect 42441 30073 42475 30107
rect 43545 30073 43579 30107
rect 51181 30073 51215 30107
rect 7665 30005 7699 30039
rect 10609 30005 10643 30039
rect 16681 30005 16715 30039
rect 17141 30005 17175 30039
rect 20913 30005 20947 30039
rect 24133 30005 24167 30039
rect 24961 30005 24995 30039
rect 36093 30005 36127 30039
rect 40601 30005 40635 30039
rect 45293 30005 45327 30039
rect 48329 30005 48363 30039
rect 52837 30005 52871 30039
rect 53205 30005 53239 30039
rect 57069 30005 57103 30039
rect 2237 29801 2271 29835
rect 9689 29801 9723 29835
rect 9873 29801 9907 29835
rect 10701 29801 10735 29835
rect 10885 29801 10919 29835
rect 13001 29801 13035 29835
rect 14473 29801 14507 29835
rect 15393 29801 15427 29835
rect 15853 29801 15887 29835
rect 19349 29801 19383 29835
rect 22937 29801 22971 29835
rect 27537 29801 27571 29835
rect 30297 29801 30331 29835
rect 32965 29801 32999 29835
rect 36829 29801 36863 29835
rect 37473 29801 37507 29835
rect 42809 29801 42843 29835
rect 45385 29801 45419 29835
rect 48329 29801 48363 29835
rect 9321 29733 9355 29767
rect 19901 29733 19935 29767
rect 23673 29733 23707 29767
rect 23765 29733 23799 29767
rect 42993 29733 43027 29767
rect 47869 29733 47903 29767
rect 48697 29733 48731 29767
rect 3893 29665 3927 29699
rect 5733 29665 5767 29699
rect 6009 29665 6043 29699
rect 7665 29665 7699 29699
rect 21649 29665 21683 29699
rect 23581 29665 23615 29699
rect 30941 29665 30975 29699
rect 32689 29665 32723 29699
rect 32781 29665 32815 29699
rect 56057 29665 56091 29699
rect 57345 29665 57379 29699
rect 1685 29597 1719 29631
rect 3985 29597 4019 29631
rect 5641 29597 5675 29631
rect 7389 29597 7423 29631
rect 10333 29597 10367 29631
rect 12449 29597 12483 29631
rect 12817 29597 12851 29631
rect 15025 29597 15059 29631
rect 15209 29597 15243 29631
rect 16037 29597 16071 29631
rect 16221 29597 16255 29631
rect 19257 29597 19291 29631
rect 23489 29597 23523 29631
rect 23857 29597 23891 29631
rect 24409 29597 24443 29631
rect 24593 29597 24627 29631
rect 24685 29597 24719 29631
rect 24777 29597 24811 29631
rect 27721 29597 27755 29631
rect 27997 29597 28031 29631
rect 28181 29597 28215 29631
rect 31033 29597 31067 29631
rect 31861 29597 31895 29631
rect 36461 29597 36495 29631
rect 36645 29597 36679 29631
rect 37289 29597 37323 29631
rect 37473 29597 37507 29631
rect 40417 29597 40451 29631
rect 40693 29597 40727 29631
rect 45017 29597 45051 29631
rect 45201 29597 45235 29631
rect 47685 29597 47719 29631
rect 47869 29597 47903 29631
rect 48513 29597 48547 29631
rect 48789 29597 48823 29631
rect 52101 29597 52135 29631
rect 53021 29597 53055 29631
rect 55321 29597 55355 29631
rect 55689 29597 55723 29631
rect 56333 29597 56367 29631
rect 56793 29597 56827 29631
rect 57253 29597 57287 29631
rect 57529 29597 57563 29631
rect 57805 29597 57839 29631
rect 57989 29597 58023 29631
rect 12633 29529 12667 29563
rect 12725 29529 12759 29563
rect 21465 29529 21499 29563
rect 42625 29529 42659 29563
rect 51549 29529 51583 29563
rect 1501 29461 1535 29495
rect 4353 29461 4387 29495
rect 4905 29461 4939 29495
rect 9689 29461 9723 29495
rect 10701 29461 10735 29495
rect 18613 29461 18647 29495
rect 22201 29461 22235 29495
rect 25053 29461 25087 29495
rect 32321 29461 32355 29495
rect 40509 29461 40543 29495
rect 40877 29461 40911 29495
rect 42825 29461 42859 29495
rect 5641 29257 5675 29291
rect 7297 29257 7331 29291
rect 10977 29257 11011 29291
rect 15025 29257 15059 29291
rect 20545 29257 20579 29291
rect 21189 29257 21223 29291
rect 23581 29257 23615 29291
rect 30757 29257 30791 29291
rect 32321 29257 32355 29291
rect 34437 29257 34471 29291
rect 49617 29257 49651 29291
rect 51733 29257 51767 29291
rect 54953 29257 54987 29291
rect 56885 29257 56919 29291
rect 6929 29189 6963 29223
rect 7113 29189 7147 29223
rect 19165 29189 19199 29223
rect 19901 29189 19935 29223
rect 5273 29121 5307 29155
rect 9321 29121 9355 29155
rect 10425 29121 10459 29155
rect 10609 29121 10643 29155
rect 10701 29121 10735 29155
rect 10793 29121 10827 29155
rect 13376 29121 13410 29155
rect 13517 29121 13551 29155
rect 13645 29121 13679 29155
rect 13737 29121 13771 29155
rect 13875 29121 13909 29155
rect 14473 29121 14507 29155
rect 14657 29121 14691 29155
rect 14749 29121 14783 29155
rect 14887 29121 14921 29155
rect 15485 29121 15519 29155
rect 17509 29121 17543 29155
rect 17785 29121 17819 29155
rect 23489 29121 23523 29155
rect 23673 29121 23707 29155
rect 26985 29121 27019 29155
rect 27169 29121 27203 29155
rect 27905 29121 27939 29155
rect 28181 29121 28215 29155
rect 28825 29121 28859 29155
rect 30389 29121 30423 29155
rect 32229 29121 32263 29155
rect 34069 29121 34103 29155
rect 34897 29121 34931 29155
rect 43085 29121 43119 29155
rect 45109 29121 45143 29155
rect 48421 29121 48455 29155
rect 49433 29121 49467 29155
rect 51917 29121 51951 29155
rect 52101 29121 52135 29155
rect 55689 29121 55723 29155
rect 57345 29121 57379 29155
rect 58173 29121 58207 29155
rect 5365 29053 5399 29087
rect 12081 29053 12115 29087
rect 12357 29053 12391 29087
rect 20085 29053 20119 29087
rect 24133 29053 24167 29087
rect 24409 29053 24443 29087
rect 26433 29053 26467 29087
rect 28641 29053 28675 29087
rect 29009 29053 29043 29087
rect 30297 29053 30331 29087
rect 33977 29053 34011 29087
rect 42901 29053 42935 29087
rect 44741 29053 44775 29087
rect 45017 29053 45051 29087
rect 48513 29053 48547 29087
rect 49249 29053 49283 29087
rect 55873 29053 55907 29087
rect 9505 28985 9539 29019
rect 14013 28985 14047 29019
rect 18061 28985 18095 29019
rect 19349 28985 19383 29019
rect 27169 28985 27203 29019
rect 29469 28985 29503 29019
rect 43269 28985 43303 29019
rect 48789 28985 48823 29019
rect 57989 28985 58023 29019
rect 7113 28917 7147 28951
rect 22201 28917 22235 28951
rect 22661 28917 22695 28951
rect 27629 28917 27663 28951
rect 28089 28917 28123 28951
rect 57069 28917 57103 28951
rect 9137 28713 9171 28747
rect 18613 28713 18647 28747
rect 23765 28713 23799 28747
rect 25237 28713 25271 28747
rect 42533 28713 42567 28747
rect 48513 28713 48547 28747
rect 51365 28713 51399 28747
rect 57621 28713 57655 28747
rect 58173 28713 58207 28747
rect 24593 28645 24627 28679
rect 27445 28645 27479 28679
rect 31585 28645 31619 28679
rect 35265 28645 35299 28679
rect 39221 28645 39255 28679
rect 11989 28577 12023 28611
rect 21557 28577 21591 28611
rect 21833 28577 21867 28611
rect 22569 28577 22603 28611
rect 27721 28577 27755 28611
rect 34805 28577 34839 28611
rect 37565 28577 37599 28611
rect 37933 28577 37967 28611
rect 38761 28577 38795 28611
rect 42257 28577 42291 28611
rect 8953 28509 8987 28543
rect 9137 28509 9171 28543
rect 9689 28509 9723 28543
rect 9873 28509 9907 28543
rect 11161 28509 11195 28543
rect 12265 28509 12299 28543
rect 14657 28509 14691 28543
rect 18521 28509 18555 28543
rect 18705 28509 18739 28543
rect 20269 28509 20303 28543
rect 21465 28509 21499 28543
rect 22477 28509 22511 28543
rect 23673 28509 23707 28543
rect 23857 28509 23891 28543
rect 24409 28509 24443 28543
rect 28181 28509 28215 28543
rect 28365 28509 28399 28543
rect 34897 28509 34931 28543
rect 37749 28509 37783 28543
rect 38853 28509 38887 28543
rect 42349 28509 42383 28543
rect 45477 28509 45511 28543
rect 45661 28509 45695 28543
rect 48053 28509 48087 28543
rect 48329 28509 48363 28543
rect 49433 28509 49467 28543
rect 49617 28509 49651 28543
rect 51549 28509 51583 28543
rect 57161 28509 57195 28543
rect 57437 28509 57471 28543
rect 9965 28441 9999 28475
rect 10977 28441 11011 28475
rect 19533 28441 19567 28475
rect 31217 28441 31251 28475
rect 31401 28441 31435 28475
rect 45569 28441 45603 28475
rect 48145 28441 48179 28475
rect 51273 28441 51307 28475
rect 51457 28441 51491 28475
rect 7021 28373 7055 28407
rect 7665 28373 7699 28407
rect 14565 28373 14599 28407
rect 22845 28373 22879 28407
rect 27261 28373 27295 28407
rect 28549 28373 28583 28407
rect 30665 28373 30699 28407
rect 41889 28373 41923 28407
rect 49617 28373 49651 28407
rect 56149 28373 56183 28407
rect 57253 28373 57287 28407
rect 6729 28169 6763 28203
rect 9781 28169 9815 28203
rect 14381 28169 14415 28203
rect 25421 28169 25455 28203
rect 31401 28169 31435 28203
rect 36737 28169 36771 28203
rect 42901 28169 42935 28203
rect 55321 28169 55355 28203
rect 56977 28169 57011 28203
rect 6929 28101 6963 28135
rect 7573 28101 7607 28135
rect 8401 28101 8435 28135
rect 15025 28101 15059 28135
rect 41613 28101 41647 28135
rect 51457 28101 51491 28135
rect 57145 28101 57179 28135
rect 57345 28101 57379 28135
rect 3709 28033 3743 28067
rect 9597 28033 9631 28067
rect 13921 28033 13955 28067
rect 14657 28033 14691 28067
rect 14933 28033 14967 28067
rect 16957 28033 16991 28067
rect 17233 28033 17267 28067
rect 22477 28033 22511 28067
rect 24685 28033 24719 28067
rect 24869 28033 24903 28067
rect 25329 28033 25363 28067
rect 25513 28033 25547 28067
rect 31033 28033 31067 28067
rect 36369 28033 36403 28067
rect 36553 28033 36587 28067
rect 39129 28033 39163 28067
rect 39313 28033 39347 28067
rect 41061 28033 41095 28067
rect 41153 28033 41187 28067
rect 41337 28033 41371 28067
rect 41429 28033 41463 28067
rect 42533 28033 42567 28067
rect 42625 28033 42659 28067
rect 42717 28033 42751 28067
rect 44741 28033 44775 28067
rect 51089 28033 51123 28067
rect 51237 28033 51271 28067
rect 51365 28033 51399 28067
rect 51595 28033 51629 28067
rect 55505 28033 55539 28067
rect 55597 28033 55631 28067
rect 55965 28033 55999 28067
rect 2789 27965 2823 27999
rect 3065 27965 3099 27999
rect 3617 27965 3651 27999
rect 4077 27965 4111 27999
rect 9413 27965 9447 27999
rect 13645 27965 13679 27999
rect 14565 27965 14599 27999
rect 20729 27965 20763 27999
rect 22017 27965 22051 27999
rect 22753 27965 22787 27999
rect 25973 27965 26007 27999
rect 30941 27965 30975 27999
rect 39221 27965 39255 27999
rect 45017 27965 45051 27999
rect 55689 27965 55723 27999
rect 55781 27965 55815 27999
rect 4629 27897 4663 27931
rect 8217 27897 8251 27931
rect 44833 27897 44867 27931
rect 6561 27829 6595 27863
rect 6745 27829 6779 27863
rect 7481 27829 7515 27863
rect 15577 27829 15611 27863
rect 18245 27829 18279 27863
rect 24225 27829 24259 27863
rect 24777 27829 24811 27863
rect 29653 27829 29687 27863
rect 30389 27829 30423 27863
rect 44925 27829 44959 27863
rect 51733 27829 51767 27863
rect 57161 27829 57195 27863
rect 3249 27625 3283 27659
rect 45477 27625 45511 27659
rect 48697 27625 48731 27659
rect 51457 27625 51491 27659
rect 2053 27557 2087 27591
rect 5641 27557 5675 27591
rect 14749 27557 14783 27591
rect 15301 27557 15335 27591
rect 16865 27557 16899 27591
rect 17049 27557 17083 27591
rect 17601 27557 17635 27591
rect 22753 27557 22787 27591
rect 30941 27557 30975 27591
rect 33057 27557 33091 27591
rect 38577 27557 38611 27591
rect 41521 27557 41555 27591
rect 47777 27557 47811 27591
rect 48513 27557 48547 27591
rect 52377 27557 52411 27591
rect 56977 27557 57011 27591
rect 57989 27557 58023 27591
rect 2513 27489 2547 27523
rect 6929 27489 6963 27523
rect 13185 27489 13219 27523
rect 16589 27489 16623 27523
rect 21005 27489 21039 27523
rect 22385 27489 22419 27523
rect 25053 27489 25087 27523
rect 25513 27489 25547 27523
rect 32597 27489 32631 27523
rect 33609 27489 33643 27523
rect 38117 27489 38151 27523
rect 41245 27489 41279 27523
rect 45109 27489 45143 27523
rect 47317 27489 47351 27523
rect 56517 27489 56551 27523
rect 2421 27421 2455 27455
rect 5917 27421 5951 27455
rect 6377 27421 6411 27455
rect 6469 27421 6503 27455
rect 6653 27421 6687 27455
rect 6745 27421 6779 27455
rect 8401 27421 8435 27455
rect 13093 27421 13127 27455
rect 13277 27421 13311 27455
rect 14105 27421 14139 27455
rect 14289 27421 14323 27455
rect 14381 27421 14415 27455
rect 14473 27421 14507 27455
rect 23397 27421 23431 27455
rect 23673 27421 23707 27455
rect 25145 27421 25179 27455
rect 26157 27421 26191 27455
rect 26341 27421 26375 27455
rect 26801 27421 26835 27455
rect 26985 27421 27019 27455
rect 27169 27421 27203 27455
rect 27905 27421 27939 27455
rect 28089 27421 28123 27455
rect 28365 27421 28399 27455
rect 29837 27421 29871 27455
rect 30113 27421 30147 27455
rect 30757 27421 30791 27455
rect 32689 27421 32723 27455
rect 36277 27421 36311 27455
rect 36461 27421 36495 27455
rect 38209 27421 38243 27455
rect 41337 27421 41371 27455
rect 41613 27421 41647 27455
rect 45201 27421 45235 27455
rect 47409 27421 47443 27455
rect 49157 27421 49191 27455
rect 49341 27421 49375 27455
rect 50997 27421 51031 27455
rect 51273 27421 51307 27455
rect 52193 27421 52227 27455
rect 54125 27421 54159 27455
rect 54677 27421 54711 27455
rect 55321 27421 55355 27455
rect 55505 27421 55539 27455
rect 55781 27421 55815 27455
rect 56609 27421 56643 27455
rect 58173 27421 58207 27455
rect 5641 27353 5675 27387
rect 7665 27353 7699 27387
rect 8309 27353 8343 27387
rect 10517 27353 10551 27387
rect 10701 27353 10735 27387
rect 48237 27353 48271 27387
rect 5825 27285 5859 27319
rect 7573 27285 7607 27319
rect 8953 27285 8987 27319
rect 18153 27285 18187 27319
rect 22845 27285 22879 27319
rect 23397 27285 23431 27319
rect 26249 27285 26283 27319
rect 28549 27285 28583 27319
rect 36461 27285 36495 27319
rect 41245 27285 41279 27319
rect 49249 27285 49283 27319
rect 51089 27285 51123 27319
rect 55965 27285 55999 27319
rect 5825 27081 5859 27115
rect 7389 27081 7423 27115
rect 7849 27081 7883 27115
rect 13093 27081 13127 27115
rect 15117 27081 15151 27115
rect 17969 27081 18003 27115
rect 19073 27081 19107 27115
rect 35357 27081 35391 27115
rect 38945 27081 38979 27115
rect 41337 27081 41371 27115
rect 44649 27081 44683 27115
rect 45109 27081 45143 27115
rect 50813 27081 50847 27115
rect 55873 27081 55907 27115
rect 58173 27081 58207 27115
rect 1869 27013 1903 27047
rect 5181 27013 5215 27047
rect 8017 27013 8051 27047
rect 8217 27013 8251 27047
rect 10057 27013 10091 27047
rect 10257 27013 10291 27047
rect 12081 27013 12115 27047
rect 13737 27013 13771 27047
rect 14013 27013 14047 27047
rect 15853 27013 15887 27047
rect 27261 27013 27295 27047
rect 27445 27013 27479 27047
rect 29101 27013 29135 27047
rect 38761 27013 38795 27047
rect 40325 27013 40359 27047
rect 40969 27013 41003 27047
rect 41169 27013 41203 27047
rect 53757 27013 53791 27047
rect 5641 26945 5675 26979
rect 6837 26945 6871 26979
rect 6929 26945 6963 26979
rect 7113 26945 7147 26979
rect 7205 26945 7239 26979
rect 13609 26945 13643 26979
rect 13829 26945 13863 26979
rect 14473 26945 14507 26979
rect 14566 26945 14600 26979
rect 14749 26945 14783 26979
rect 14841 26945 14875 26979
rect 14979 26945 15013 26979
rect 15669 26945 15703 26979
rect 20269 26945 20303 26979
rect 22753 26945 22787 26979
rect 22937 26945 22971 26979
rect 28089 26945 28123 26979
rect 34989 26945 35023 26979
rect 38577 26945 38611 26979
rect 40233 26945 40267 26979
rect 40509 26945 40543 26979
rect 44281 26945 44315 26979
rect 45109 26945 45143 26979
rect 45293 26945 45327 26979
rect 50721 26945 50755 26979
rect 50905 26945 50939 26979
rect 53389 26945 53423 26979
rect 53573 26945 53607 26979
rect 55689 26945 55723 26979
rect 55965 26945 55999 26979
rect 56977 26945 57011 26979
rect 13921 26877 13955 26911
rect 20361 26877 20395 26911
rect 28365 26877 28399 26911
rect 34897 26877 34931 26911
rect 44189 26877 44223 26911
rect 56885 26877 56919 26911
rect 2053 26809 2087 26843
rect 11897 26809 11931 26843
rect 28641 26809 28675 26843
rect 29377 26809 29411 26843
rect 40509 26809 40543 26843
rect 55689 26809 55723 26843
rect 8033 26741 8067 26775
rect 10241 26741 10275 26775
rect 10425 26741 10459 26775
rect 20637 26741 20671 26775
rect 21097 26741 21131 26775
rect 22845 26741 22879 26775
rect 27629 26741 27663 26775
rect 28181 26741 28215 26775
rect 29561 26741 29595 26775
rect 41153 26741 41187 26775
rect 57345 26741 57379 26775
rect 1685 26537 1719 26571
rect 3893 26537 3927 26571
rect 6469 26537 6503 26571
rect 10701 26537 10735 26571
rect 14105 26537 14139 26571
rect 18705 26537 18739 26571
rect 19901 26537 19935 26571
rect 24501 26537 24535 26571
rect 34161 26537 34195 26571
rect 34805 26537 34839 26571
rect 35173 26537 35207 26571
rect 41429 26537 41463 26571
rect 50721 26537 50755 26571
rect 53113 26537 53147 26571
rect 55965 26537 55999 26571
rect 17601 26469 17635 26503
rect 21189 26469 21223 26503
rect 6929 26401 6963 26435
rect 15025 26401 15059 26435
rect 21465 26401 21499 26435
rect 22385 26401 22419 26435
rect 23213 26401 23247 26435
rect 33701 26401 33735 26435
rect 38485 26401 38519 26435
rect 41245 26401 41279 26435
rect 50261 26401 50295 26435
rect 6193 26333 6227 26367
rect 6285 26333 6319 26367
rect 6469 26333 6503 26367
rect 7205 26333 7239 26367
rect 10149 26333 10183 26367
rect 10241 26333 10275 26367
rect 10425 26333 10459 26367
rect 10517 26333 10551 26367
rect 17049 26333 17083 26367
rect 17325 26333 17359 26367
rect 17417 26333 17451 26367
rect 18061 26333 18095 26367
rect 18154 26333 18188 26367
rect 18429 26333 18463 26367
rect 18567 26333 18601 26367
rect 19257 26333 19291 26367
rect 19350 26333 19384 26367
rect 19763 26333 19797 26367
rect 22201 26333 22235 26367
rect 23305 26333 23339 26367
rect 23581 26333 23615 26367
rect 23673 26333 23707 26367
rect 24409 26333 24443 26367
rect 24593 26333 24627 26367
rect 27905 26333 27939 26367
rect 30573 26333 30607 26367
rect 30757 26333 30791 26367
rect 33793 26333 33827 26367
rect 34713 26333 34747 26367
rect 37197 26333 37231 26367
rect 37381 26333 37415 26367
rect 37749 26333 37783 26367
rect 38393 26333 38427 26367
rect 38577 26333 38611 26367
rect 41153 26333 41187 26367
rect 50353 26333 50387 26367
rect 51181 26333 51215 26367
rect 51365 26333 51399 26367
rect 52837 26333 52871 26367
rect 55965 26333 55999 26367
rect 56149 26333 56183 26367
rect 11253 26265 11287 26299
rect 11437 26265 11471 26299
rect 14841 26265 14875 26299
rect 17233 26265 17267 26299
rect 18337 26265 18371 26299
rect 19533 26265 19567 26299
rect 19625 26265 19659 26299
rect 25053 26265 25087 26299
rect 31585 26265 31619 26299
rect 37657 26265 37691 26299
rect 51549 26265 51583 26299
rect 52377 26265 52411 26299
rect 53113 26265 53147 26299
rect 53573 26265 53607 26299
rect 21005 26197 21039 26231
rect 22017 26197 22051 26231
rect 23857 26197 23891 26231
rect 27997 26197 28031 26231
rect 40785 26197 40819 26231
rect 52929 26197 52963 26231
rect 2789 25993 2823 26027
rect 6469 25993 6503 26027
rect 9965 25993 9999 26027
rect 13829 25993 13863 26027
rect 17785 25993 17819 26027
rect 18337 25993 18371 26027
rect 22017 25993 22051 26027
rect 27905 25993 27939 26027
rect 38761 25993 38795 26027
rect 44005 25993 44039 26027
rect 47961 25993 47995 26027
rect 50077 25993 50111 26027
rect 53205 25993 53239 26027
rect 53865 25993 53899 26027
rect 54033 25993 54067 26027
rect 56241 25993 56275 26027
rect 4261 25925 4295 25959
rect 13553 25925 13587 25959
rect 17509 25925 17543 25959
rect 18981 25925 19015 25959
rect 21097 25925 21131 25959
rect 24317 25925 24351 25959
rect 24409 25925 24443 25959
rect 47777 25925 47811 25959
rect 48697 25925 48731 25959
rect 53665 25925 53699 25959
rect 3157 25857 3191 25891
rect 5825 25857 5859 25891
rect 6653 25857 6687 25891
rect 8125 25857 8159 25891
rect 9229 25857 9263 25891
rect 9413 25857 9447 25891
rect 9505 25857 9539 25891
rect 10149 25857 10183 25891
rect 10241 25857 10275 25891
rect 10425 25857 10459 25891
rect 10517 25857 10551 25891
rect 11529 25857 11563 25891
rect 11713 25857 11747 25891
rect 11805 25857 11839 25891
rect 13277 25857 13311 25891
rect 13461 25857 13495 25891
rect 13645 25857 13679 25891
rect 14289 25857 14323 25891
rect 17233 25857 17267 25891
rect 17417 25857 17451 25891
rect 17601 25857 17635 25891
rect 22201 25857 22235 25891
rect 22293 25857 22327 25891
rect 24041 25857 24075 25891
rect 24189 25857 24223 25891
rect 24506 25857 24540 25891
rect 28089 25857 28123 25891
rect 30481 25857 30515 25891
rect 37473 25857 37507 25891
rect 43637 25857 43671 25891
rect 46857 25857 46891 25891
rect 47041 25857 47075 25891
rect 47593 25857 47627 25891
rect 49985 25857 50019 25891
rect 50169 25857 50203 25891
rect 52745 25857 52779 25891
rect 52837 25857 52871 25891
rect 53021 25857 53055 25891
rect 55873 25857 55907 25891
rect 3065 25789 3099 25823
rect 7849 25789 7883 25823
rect 28273 25789 28307 25823
rect 30389 25789 30423 25823
rect 37381 25789 37415 25823
rect 37841 25789 37875 25823
rect 38301 25789 38335 25823
rect 43729 25789 43763 25823
rect 46949 25789 46983 25823
rect 49249 25789 49283 25823
rect 55781 25789 55815 25823
rect 3985 25721 4019 25755
rect 9229 25721 9263 25755
rect 11529 25721 11563 25755
rect 14473 25721 14507 25755
rect 19165 25721 19199 25755
rect 21281 25721 21315 25755
rect 24685 25721 24719 25755
rect 38577 25721 38611 25755
rect 3801 25653 3835 25687
rect 23121 25653 23155 25687
rect 30757 25653 30791 25687
rect 53849 25653 53883 25687
rect 6561 25449 6595 25483
rect 10149 25449 10183 25483
rect 10333 25449 10367 25483
rect 18521 25449 18555 25483
rect 21741 25449 21775 25483
rect 43821 25449 43855 25483
rect 46489 25449 46523 25483
rect 50169 25449 50203 25483
rect 52837 25449 52871 25483
rect 54677 25449 54711 25483
rect 55965 25449 55999 25483
rect 4353 25381 4387 25415
rect 17233 25381 17267 25415
rect 20545 25381 20579 25415
rect 30665 25381 30699 25415
rect 31769 25381 31803 25415
rect 35265 25381 35299 25415
rect 38025 25381 38059 25415
rect 38117 25381 38151 25415
rect 7757 25313 7791 25347
rect 23673 25313 23707 25347
rect 28917 25313 28951 25347
rect 31309 25313 31343 25347
rect 34805 25313 34839 25347
rect 40509 25313 40543 25347
rect 50261 25313 50295 25347
rect 52837 25313 52871 25347
rect 52929 25313 52963 25347
rect 53113 25313 53147 25347
rect 55597 25313 55631 25347
rect 55781 25313 55815 25347
rect 2053 25245 2087 25279
rect 2697 25245 2731 25279
rect 2973 25245 3007 25279
rect 3065 25245 3099 25279
rect 3801 25245 3835 25279
rect 4169 25245 4203 25279
rect 4813 25245 4847 25279
rect 4997 25245 5031 25279
rect 8033 25245 8067 25279
rect 13001 25245 13035 25279
rect 13369 25245 13403 25279
rect 14105 25245 14139 25279
rect 14253 25245 14287 25279
rect 14611 25245 14645 25279
rect 16681 25245 16715 25279
rect 17049 25245 17083 25279
rect 17877 25245 17911 25279
rect 17970 25245 18004 25279
rect 18245 25245 18279 25279
rect 18342 25245 18376 25279
rect 21649 25245 21683 25279
rect 22937 25245 22971 25279
rect 23581 25245 23615 25279
rect 23765 25245 23799 25279
rect 24409 25245 24443 25279
rect 24557 25245 24591 25279
rect 24874 25245 24908 25279
rect 27629 25245 27663 25279
rect 27813 25245 27847 25279
rect 28365 25245 28399 25279
rect 28733 25245 28767 25279
rect 31401 25245 31435 25279
rect 34897 25245 34931 25279
rect 35725 25245 35759 25279
rect 40141 25245 40175 25279
rect 40969 25245 41003 25279
rect 41153 25245 41187 25279
rect 41337 25245 41371 25279
rect 41981 25245 42015 25279
rect 42165 25245 42199 25279
rect 42625 25245 42659 25279
rect 42809 25245 42843 25279
rect 42993 25245 43027 25279
rect 43729 25245 43763 25279
rect 45845 25245 45879 25279
rect 46029 25245 46063 25279
rect 46121 25245 46155 25279
rect 46259 25245 46293 25279
rect 50169 25245 50203 25279
rect 53205 25245 53239 25279
rect 54585 25245 54619 25279
rect 55505 25245 55539 25279
rect 55689 25245 55723 25279
rect 57897 25245 57931 25279
rect 1869 25177 1903 25211
rect 2881 25177 2915 25211
rect 3985 25177 4019 25211
rect 4077 25177 4111 25211
rect 4905 25177 4939 25211
rect 6377 25177 6411 25211
rect 6577 25177 6611 25211
rect 9965 25177 9999 25211
rect 10181 25177 10215 25211
rect 13185 25177 13219 25211
rect 13277 25177 13311 25211
rect 14381 25177 14415 25211
rect 14473 25177 14507 25211
rect 16865 25177 16899 25211
rect 16957 25177 16991 25211
rect 18153 25177 18187 25211
rect 22753 25177 22787 25211
rect 24685 25177 24719 25211
rect 24777 25177 24811 25211
rect 37657 25177 37691 25211
rect 40325 25177 40359 25211
rect 41797 25177 41831 25211
rect 3249 25109 3283 25143
rect 6745 25109 6779 25143
rect 13553 25109 13587 25143
rect 14749 25109 14783 25143
rect 25053 25109 25087 25143
rect 27537 25109 27571 25143
rect 34069 25109 34103 25143
rect 44189 25109 44223 25143
rect 50537 25109 50571 25143
rect 58081 25109 58115 25143
rect 1685 24905 1719 24939
rect 3249 24905 3283 24939
rect 4077 24905 4111 24939
rect 27997 24905 28031 24939
rect 34989 24905 35023 24939
rect 40233 24905 40267 24939
rect 50077 24905 50111 24939
rect 57989 24905 58023 24939
rect 8217 24837 8251 24871
rect 17877 24837 17911 24871
rect 45017 24837 45051 24871
rect 46213 24837 46247 24871
rect 55689 24837 55723 24871
rect 55781 24837 55815 24871
rect 2513 24769 2547 24803
rect 2697 24769 2731 24803
rect 3157 24769 3191 24803
rect 3433 24769 3467 24803
rect 6929 24769 6963 24803
rect 7021 24769 7055 24803
rect 7205 24769 7239 24803
rect 7297 24769 7331 24803
rect 7481 24769 7515 24803
rect 8033 24769 8067 24803
rect 8318 24791 8352 24825
rect 9689 24769 9723 24803
rect 10241 24769 10275 24803
rect 13461 24769 13495 24803
rect 17141 24769 17175 24803
rect 20085 24769 20119 24803
rect 20729 24769 20763 24803
rect 20913 24769 20947 24803
rect 23489 24769 23523 24803
rect 24409 24769 24443 24803
rect 25697 24769 25731 24803
rect 26157 24769 26191 24803
rect 27905 24769 27939 24803
rect 28089 24769 28123 24803
rect 30573 24769 30607 24803
rect 33977 24769 34011 24803
rect 34897 24769 34931 24803
rect 37749 24769 37783 24803
rect 40049 24769 40083 24803
rect 40233 24769 40267 24803
rect 41613 24769 41647 24803
rect 41797 24769 41831 24803
rect 44281 24769 44315 24803
rect 44557 24769 44591 24803
rect 44925 24769 44959 24803
rect 45753 24769 45787 24803
rect 45845 24769 45879 24803
rect 46029 24769 46063 24803
rect 50721 24769 50755 24803
rect 51089 24769 51123 24803
rect 55413 24769 55447 24803
rect 55505 24769 55539 24803
rect 55873 24769 55907 24803
rect 56885 24769 56919 24803
rect 56977 24769 57011 24803
rect 57161 24769 57195 24803
rect 57345 24769 57379 24803
rect 57897 24769 57931 24803
rect 57989 24769 58023 24803
rect 58173 24769 58207 24803
rect 2329 24701 2363 24735
rect 13277 24701 13311 24735
rect 25329 24701 25363 24735
rect 30297 24701 30331 24735
rect 31125 24701 31159 24735
rect 33885 24701 33919 24735
rect 37841 24701 37875 24735
rect 41705 24701 41739 24735
rect 45109 24701 45143 24735
rect 46121 24701 46155 24735
rect 8033 24633 8067 24667
rect 9505 24633 9539 24667
rect 13645 24633 13679 24667
rect 17325 24633 17359 24667
rect 18061 24633 18095 24667
rect 20269 24633 20303 24667
rect 24225 24633 24259 24667
rect 34345 24633 34379 24667
rect 56057 24633 56091 24667
rect 3617 24565 3651 24599
rect 10425 24565 10459 24599
rect 14105 24565 14139 24599
rect 20729 24565 20763 24599
rect 28549 24565 28583 24599
rect 33241 24565 33275 24599
rect 37749 24565 37783 24599
rect 38117 24565 38151 24599
rect 49525 24565 49559 24599
rect 3893 24361 3927 24395
rect 7757 24361 7791 24395
rect 10701 24361 10735 24395
rect 13093 24361 13127 24395
rect 17969 24361 18003 24395
rect 21465 24361 21499 24395
rect 25145 24361 25179 24395
rect 27721 24361 27755 24395
rect 27905 24361 27939 24395
rect 28549 24361 28583 24395
rect 31125 24361 31159 24395
rect 33977 24361 34011 24395
rect 38209 24361 38243 24395
rect 38577 24361 38611 24395
rect 39129 24361 39163 24395
rect 39221 24361 39255 24395
rect 42257 24361 42291 24395
rect 45661 24361 45695 24395
rect 56333 24361 56367 24395
rect 13277 24293 13311 24327
rect 14749 24293 14783 24327
rect 20361 24293 20395 24327
rect 27169 24293 27203 24327
rect 37657 24293 37691 24327
rect 41429 24293 41463 24327
rect 43913 24293 43947 24327
rect 18613 24225 18647 24259
rect 37381 24225 37415 24259
rect 39313 24225 39347 24259
rect 40969 24225 41003 24259
rect 48881 24225 48915 24259
rect 53113 24225 53147 24259
rect 7573 24157 7607 24191
rect 8309 24157 8343 24191
rect 10149 24157 10183 24191
rect 10241 24157 10275 24191
rect 10425 24157 10459 24191
rect 10517 24157 10551 24191
rect 11529 24157 11563 24191
rect 14105 24157 14139 24191
rect 14198 24157 14232 24191
rect 14473 24157 14507 24191
rect 14570 24157 14604 24191
rect 16313 24157 16347 24191
rect 16589 24157 16623 24191
rect 16681 24157 16715 24191
rect 17325 24157 17359 24191
rect 17418 24157 17452 24191
rect 17790 24157 17824 24191
rect 19809 24157 19843 24191
rect 20085 24157 20119 24191
rect 20177 24157 20211 24191
rect 20821 24157 20855 24191
rect 20969 24157 21003 24191
rect 21327 24157 21361 24191
rect 23489 24157 23523 24191
rect 24501 24157 24535 24191
rect 24594 24157 24628 24191
rect 24869 24157 24903 24191
rect 25007 24157 25041 24191
rect 28549 24157 28583 24191
rect 28825 24157 28859 24191
rect 30389 24157 30423 24191
rect 33425 24157 33459 24191
rect 33885 24157 33919 24191
rect 34713 24157 34747 24191
rect 37289 24157 37323 24191
rect 38117 24157 38151 24191
rect 39037 24157 39071 24191
rect 41061 24157 41095 24191
rect 42073 24157 42107 24191
rect 43637 24157 43671 24191
rect 45017 24157 45051 24191
rect 45201 24157 45235 24191
rect 45293 24157 45327 24191
rect 45385 24157 45419 24191
rect 47869 24157 47903 24191
rect 48053 24157 48087 24191
rect 52653 24157 52687 24191
rect 52929 24157 52963 24191
rect 53297 24157 53331 24191
rect 55321 24157 55355 24191
rect 55413 24157 55447 24191
rect 55597 24157 55631 24191
rect 55689 24157 55723 24191
rect 58173 24157 58207 24191
rect 9413 24089 9447 24123
rect 9597 24089 9631 24123
rect 11345 24089 11379 24123
rect 13553 24089 13587 24123
rect 14381 24089 14415 24123
rect 16497 24089 16531 24123
rect 17601 24089 17635 24123
rect 17693 24089 17727 24123
rect 19993 24089 20027 24123
rect 21097 24089 21131 24123
rect 21189 24089 21223 24123
rect 24777 24089 24811 24123
rect 27873 24089 27907 24123
rect 28089 24089 28123 24123
rect 30941 24089 30975 24123
rect 34989 24089 35023 24123
rect 41889 24089 41923 24123
rect 43913 24089 43947 24123
rect 56517 24089 56551 24123
rect 56701 24089 56735 24123
rect 57897 24089 57931 24123
rect 16865 24021 16899 24055
rect 22017 24021 22051 24055
rect 23581 24021 23615 24055
rect 28733 24021 28767 24055
rect 29837 24021 29871 24055
rect 31125 24021 31159 24055
rect 31309 24021 31343 24055
rect 43729 24021 43763 24055
rect 55873 24021 55907 24055
rect 7021 23817 7055 23851
rect 9413 23817 9447 23851
rect 10333 23817 10367 23851
rect 10793 23817 10827 23851
rect 13829 23817 13863 23851
rect 17233 23817 17267 23851
rect 18061 23817 18095 23851
rect 19717 23817 19751 23851
rect 23029 23817 23063 23851
rect 46949 23817 46983 23851
rect 48053 23817 48087 23851
rect 53205 23817 53239 23851
rect 56057 23817 56091 23851
rect 3893 23749 3927 23783
rect 9965 23749 9999 23783
rect 16865 23749 16899 23783
rect 23489 23749 23523 23783
rect 24961 23749 24995 23783
rect 25789 23749 25823 23783
rect 25973 23749 26007 23783
rect 34805 23749 34839 23783
rect 37933 23749 37967 23783
rect 43729 23749 43763 23783
rect 43945 23749 43979 23783
rect 46305 23749 46339 23783
rect 10195 23715 10229 23749
rect 2237 23681 2271 23715
rect 2513 23681 2547 23715
rect 5457 23681 5491 23715
rect 6837 23681 6871 23715
rect 7573 23681 7607 23715
rect 7757 23681 7791 23715
rect 8769 23681 8803 23715
rect 9229 23681 9263 23715
rect 9505 23681 9539 23715
rect 12449 23681 12483 23715
rect 12633 23681 12667 23715
rect 12721 23681 12755 23715
rect 12817 23681 12851 23715
rect 13645 23681 13679 23715
rect 16681 23681 16715 23715
rect 16957 23681 16991 23715
rect 17049 23681 17083 23715
rect 17969 23681 18003 23715
rect 18889 23681 18923 23715
rect 19625 23681 19659 23715
rect 19809 23681 19843 23715
rect 20443 23703 20477 23737
rect 20545 23681 20579 23715
rect 20656 23681 20690 23715
rect 20821 23681 20855 23715
rect 23857 23681 23891 23715
rect 23949 23681 23983 23715
rect 24600 23681 24634 23715
rect 24686 23681 24720 23715
rect 24869 23681 24903 23715
rect 25058 23681 25092 23715
rect 30941 23681 30975 23715
rect 34621 23681 34655 23715
rect 34897 23681 34931 23715
rect 37289 23681 37323 23715
rect 37473 23681 37507 23715
rect 37749 23681 37783 23715
rect 40141 23681 40175 23715
rect 46857 23681 46891 23715
rect 47041 23681 47075 23715
rect 50353 23681 50387 23715
rect 50537 23681 50571 23715
rect 50997 23681 51031 23715
rect 51181 23681 51215 23715
rect 51641 23681 51675 23715
rect 53021 23681 53055 23715
rect 55965 23681 55999 23715
rect 56149 23681 56183 23715
rect 5365 23613 5399 23647
rect 5825 23613 5859 23647
rect 7941 23613 7975 23647
rect 13461 23613 13495 23647
rect 23581 23613 23615 23647
rect 30757 23613 30791 23647
rect 31309 23613 31343 23647
rect 39405 23613 39439 23647
rect 40049 23613 40083 23647
rect 47593 23613 47627 23647
rect 52745 23613 52779 23647
rect 9229 23545 9263 23579
rect 13001 23545 13035 23579
rect 21005 23545 21039 23579
rect 24133 23545 24167 23579
rect 30205 23545 30239 23579
rect 31217 23545 31251 23579
rect 44097 23545 44131 23579
rect 47869 23545 47903 23579
rect 50445 23545 50479 23579
rect 4813 23477 4847 23511
rect 10149 23477 10183 23511
rect 14289 23477 14323 23511
rect 19073 23477 19107 23511
rect 25237 23477 25271 23511
rect 28365 23477 28399 23511
rect 29653 23477 29687 23511
rect 34621 23477 34655 23511
rect 36737 23477 36771 23511
rect 40417 23477 40451 23511
rect 43913 23477 43947 23511
rect 51089 23477 51123 23511
rect 52837 23477 52871 23511
rect 58081 23477 58115 23511
rect 4353 23273 4387 23307
rect 13001 23273 13035 23307
rect 14289 23273 14323 23307
rect 23857 23273 23891 23307
rect 30389 23273 30423 23307
rect 34989 23273 35023 23307
rect 54769 23273 54803 23307
rect 55505 23273 55539 23307
rect 6469 23205 6503 23239
rect 7389 23205 7423 23239
rect 8217 23205 8251 23239
rect 23213 23205 23247 23239
rect 35173 23205 35207 23239
rect 53481 23205 53515 23239
rect 6193 23137 6227 23171
rect 7021 23137 7055 23171
rect 7481 23137 7515 23171
rect 16589 23137 16623 23171
rect 26709 23137 26743 23171
rect 29561 23137 29595 23171
rect 32413 23137 32447 23171
rect 44005 23137 44039 23171
rect 44189 23137 44223 23171
rect 46489 23137 46523 23171
rect 51181 23137 51215 23171
rect 52101 23137 52135 23171
rect 1869 23069 1903 23103
rect 4261 23069 4295 23103
rect 6101 23069 6135 23103
rect 8033 23069 8067 23103
rect 9873 23069 9907 23103
rect 10149 23069 10183 23103
rect 17325 23069 17359 23103
rect 17509 23069 17543 23103
rect 17693 23069 17727 23103
rect 23029 23069 23063 23103
rect 23673 23069 23707 23103
rect 23857 23069 23891 23103
rect 24869 23069 24903 23103
rect 26801 23069 26835 23103
rect 27629 23069 27663 23103
rect 28825 23069 28859 23103
rect 29009 23069 29043 23103
rect 29745 23069 29779 23103
rect 29929 23069 29963 23103
rect 30573 23069 30607 23103
rect 30849 23069 30883 23103
rect 31401 23069 31435 23103
rect 43913 23069 43947 23103
rect 46029 23069 46063 23103
rect 46305 23069 46339 23103
rect 47317 23069 47351 23103
rect 47409 23069 47443 23103
rect 47593 23069 47627 23103
rect 47777 23069 47811 23103
rect 50261 23069 50295 23103
rect 52469 23069 52503 23103
rect 53113 23069 53147 23103
rect 54493 23069 54527 23103
rect 54585 23069 54619 23103
rect 56517 23069 56551 23103
rect 57069 23069 57103 23103
rect 2053 23001 2087 23035
rect 5365 23001 5399 23035
rect 14105 23001 14139 23035
rect 14305 23001 14339 23035
rect 15025 23001 15059 23035
rect 15209 23001 15243 23035
rect 16773 23001 16807 23035
rect 17601 23001 17635 23035
rect 20453 23001 20487 23035
rect 30757 23001 30791 23035
rect 34805 23001 34839 23035
rect 35005 23001 35039 23035
rect 54769 23001 54803 23035
rect 55321 23001 55355 23035
rect 13461 22933 13495 22967
rect 14473 22933 14507 22967
rect 17877 22933 17911 22967
rect 24961 22933 24995 22967
rect 27169 22933 27203 22967
rect 27813 22933 27847 22967
rect 28917 22933 28951 22967
rect 33517 22933 33551 22967
rect 34161 22933 34195 22967
rect 35633 22933 35667 22967
rect 43545 22933 43579 22967
rect 46121 22933 46155 22967
rect 55521 22933 55555 22967
rect 55689 22933 55723 22967
rect 1685 22729 1719 22763
rect 5089 22729 5123 22763
rect 6653 22729 6687 22763
rect 9413 22729 9447 22763
rect 11713 22729 11747 22763
rect 15209 22729 15243 22763
rect 17233 22729 17267 22763
rect 19809 22729 19843 22763
rect 23397 22729 23431 22763
rect 28457 22729 28491 22763
rect 30297 22729 30331 22763
rect 34069 22729 34103 22763
rect 34989 22729 35023 22763
rect 35449 22729 35483 22763
rect 37841 22729 37875 22763
rect 43085 22729 43119 22763
rect 46505 22729 46539 22763
rect 46673 22729 46707 22763
rect 53389 22729 53423 22763
rect 57069 22729 57103 22763
rect 8769 22661 8803 22695
rect 8953 22661 8987 22695
rect 13093 22661 13127 22695
rect 18705 22661 18739 22695
rect 19441 22661 19475 22695
rect 21189 22661 21223 22695
rect 24593 22661 24627 22695
rect 35725 22661 35759 22695
rect 46305 22661 46339 22695
rect 50353 22661 50387 22695
rect 54493 22661 54527 22695
rect 56517 22661 56551 22695
rect 3525 22593 3559 22627
rect 3801 22593 3835 22627
rect 7665 22593 7699 22627
rect 7849 22593 7883 22627
rect 11529 22593 11563 22627
rect 12817 22593 12851 22627
rect 13001 22593 13035 22627
rect 13185 22593 13219 22627
rect 13829 22593 13863 22627
rect 13977 22593 14011 22627
rect 14105 22593 14139 22627
rect 14197 22593 14231 22627
rect 14335 22593 14369 22627
rect 15117 22593 15151 22627
rect 16681 22593 16715 22627
rect 16773 22593 16807 22627
rect 16957 22593 16991 22627
rect 17049 22593 17083 22627
rect 19165 22593 19199 22627
rect 19313 22593 19347 22627
rect 19533 22593 19567 22627
rect 19671 22593 19705 22627
rect 21833 22593 21867 22627
rect 21925 22593 21959 22627
rect 22109 22593 22143 22627
rect 22201 22593 22235 22627
rect 23857 22593 23891 22627
rect 23949 22593 23983 22627
rect 24133 22593 24167 22627
rect 25145 22593 25179 22627
rect 28089 22593 28123 22627
rect 30205 22593 30239 22627
rect 30389 22593 30423 22627
rect 33057 22593 33091 22627
rect 33701 22593 33735 22627
rect 34529 22593 34563 22627
rect 34621 22593 34655 22627
rect 34805 22593 34839 22627
rect 35449 22593 35483 22627
rect 35541 22593 35575 22627
rect 37473 22593 37507 22627
rect 40233 22593 40267 22627
rect 42533 22593 42567 22627
rect 42901 22593 42935 22627
rect 49341 22593 49375 22627
rect 52745 22593 52779 22627
rect 52929 22593 52963 22627
rect 53021 22593 53055 22627
rect 53159 22593 53193 22627
rect 54769 22593 54803 22627
rect 55137 22593 55171 22627
rect 55229 22593 55263 22627
rect 56241 22593 56275 22627
rect 56333 22593 56367 22627
rect 56977 22593 57011 22627
rect 57161 22593 57195 22627
rect 12357 22525 12391 22559
rect 22385 22525 22419 22559
rect 27997 22525 28031 22559
rect 33609 22525 33643 22559
rect 37381 22525 37415 22559
rect 40141 22525 40175 22559
rect 40601 22525 40635 22559
rect 13369 22457 13403 22491
rect 14473 22457 14507 22491
rect 16037 22457 16071 22491
rect 36645 22457 36679 22491
rect 55321 22457 55355 22491
rect 4629 22389 4663 22423
rect 10241 22389 10275 22423
rect 21097 22389 21131 22423
rect 24133 22389 24167 22423
rect 42901 22389 42935 22423
rect 46489 22389 46523 22423
rect 9321 22185 9355 22219
rect 15761 22185 15795 22219
rect 16589 22185 16623 22219
rect 20729 22185 20763 22219
rect 21741 22185 21775 22219
rect 23673 22185 23707 22219
rect 24961 22185 24995 22219
rect 34897 22185 34931 22219
rect 37197 22185 37231 22219
rect 42533 22185 42567 22219
rect 42809 22185 42843 22219
rect 46121 22185 46155 22219
rect 46581 22185 46615 22219
rect 7481 22117 7515 22151
rect 8401 22117 8435 22151
rect 23857 22117 23891 22151
rect 39313 22117 39347 22151
rect 40601 22117 40635 22151
rect 56977 22117 57011 22151
rect 7297 22049 7331 22083
rect 12817 22049 12851 22083
rect 14657 22049 14691 22083
rect 30573 22049 30607 22083
rect 36829 22049 36863 22083
rect 38853 22049 38887 22083
rect 40785 22049 40819 22083
rect 1869 21981 1903 22015
rect 2329 21981 2363 22015
rect 2513 21981 2547 22015
rect 3065 21981 3099 22015
rect 3249 21981 3283 22015
rect 4353 21981 4387 22015
rect 4629 21981 4663 22015
rect 5089 21981 5123 22015
rect 5273 21981 5307 22015
rect 7481 21981 7515 22015
rect 7849 21981 7883 22015
rect 9965 21981 9999 22015
rect 10057 21981 10091 22015
rect 10241 21981 10275 22015
rect 10333 21981 10367 22015
rect 11069 21981 11103 22015
rect 13461 21981 13495 22015
rect 14105 21981 14139 22015
rect 14473 21981 14507 22015
rect 16313 21981 16347 22015
rect 20085 21981 20119 22015
rect 20545 21981 20579 22015
rect 20729 21981 20763 22015
rect 21189 21981 21223 22015
rect 21465 21981 21499 22015
rect 21557 21981 21591 22015
rect 24409 21981 24443 22015
rect 24501 21981 24535 22015
rect 24685 21981 24719 22015
rect 24777 21981 24811 22015
rect 25697 21981 25731 22015
rect 34161 21981 34195 22015
rect 34713 21981 34747 22015
rect 36921 21981 36955 22015
rect 38945 21981 38979 22015
rect 42809 21981 42843 22015
rect 42993 21981 43027 22015
rect 45661 21981 45695 22015
rect 45937 21981 45971 22015
rect 46581 21981 46615 22015
rect 46857 21981 46891 22015
rect 56701 21981 56735 22015
rect 56977 21981 57011 22015
rect 9137 21913 9171 21947
rect 16405 21913 16439 21947
rect 16589 21913 16623 21947
rect 21373 21913 21407 21947
rect 23489 21913 23523 21947
rect 26157 21913 26191 21947
rect 40325 21913 40359 21947
rect 46673 21913 46707 21947
rect 2513 21845 2547 21879
rect 3157 21845 3191 21879
rect 4169 21845 4203 21879
rect 4537 21845 4571 21879
rect 5365 21845 5399 21879
rect 9337 21845 9371 21879
rect 9505 21845 9539 21879
rect 10517 21845 10551 21879
rect 11253 21845 11287 21879
rect 13369 21845 13403 21879
rect 14473 21845 14507 21879
rect 19349 21845 19383 21879
rect 22937 21845 22971 21879
rect 23689 21845 23723 21879
rect 25513 21845 25547 21879
rect 26801 21845 26835 21879
rect 33333 21845 33367 21879
rect 35449 21845 35483 21879
rect 38209 21845 38243 21879
rect 45753 21845 45787 21879
rect 56793 21845 56827 21879
rect 2237 21641 2271 21675
rect 9603 21641 9637 21675
rect 11529 21641 11563 21675
rect 13553 21641 13587 21675
rect 16037 21641 16071 21675
rect 19717 21641 19751 21675
rect 23121 21641 23155 21675
rect 23673 21641 23707 21675
rect 25605 21641 25639 21675
rect 31585 21641 31619 21675
rect 32781 21641 32815 21675
rect 34437 21641 34471 21675
rect 46397 21641 46431 21675
rect 49065 21641 49099 21675
rect 52193 21641 52227 21675
rect 53297 21641 53331 21675
rect 54401 21641 54435 21675
rect 56517 21641 56551 21675
rect 57069 21641 57103 21675
rect 57989 21641 58023 21675
rect 3157 21573 3191 21607
rect 9505 21573 9539 21607
rect 9689 21573 9723 21607
rect 17141 21573 17175 21607
rect 19441 21573 19475 21607
rect 20361 21573 20395 21607
rect 24225 21573 24259 21607
rect 24425 21573 24459 21607
rect 26249 21573 26283 21607
rect 1409 21505 1443 21539
rect 2145 21505 2179 21539
rect 2973 21505 3007 21539
rect 4169 21505 4203 21539
rect 4629 21505 4663 21539
rect 7113 21505 7147 21539
rect 7665 21505 7699 21539
rect 9781 21505 9815 21539
rect 10333 21505 10367 21539
rect 10517 21505 10551 21539
rect 13001 21505 13035 21539
rect 13185 21505 13219 21539
rect 13277 21505 13311 21539
rect 13369 21505 13403 21539
rect 14381 21505 14415 21539
rect 19073 21505 19107 21539
rect 19166 21505 19200 21539
rect 19349 21505 19383 21539
rect 19579 21505 19613 21539
rect 25053 21505 25087 21539
rect 25145 21505 25179 21539
rect 25329 21505 25363 21539
rect 25421 21505 25455 21539
rect 27445 21505 27479 21539
rect 27629 21505 27663 21539
rect 30573 21505 30607 21539
rect 30941 21505 30975 21539
rect 33241 21505 33275 21539
rect 35449 21505 35483 21539
rect 46397 21505 46431 21539
rect 48421 21505 48455 21539
rect 49709 21505 49743 21539
rect 49893 21505 49927 21539
rect 52009 21505 52043 21539
rect 52745 21505 52779 21539
rect 53021 21505 53055 21539
rect 53849 21505 53883 21539
rect 53941 21505 53975 21539
rect 54125 21505 54159 21539
rect 54217 21505 54251 21539
rect 56333 21505 56367 21539
rect 56977 21505 57011 21539
rect 57161 21505 57195 21539
rect 57897 21505 57931 21539
rect 2789 21437 2823 21471
rect 33333 21437 33367 21471
rect 45845 21437 45879 21471
rect 46489 21437 46523 21471
rect 48329 21437 48363 21471
rect 51733 21437 51767 21471
rect 53205 21437 53239 21471
rect 56149 21437 56183 21471
rect 27537 21369 27571 21403
rect 1593 21301 1627 21335
rect 5825 21301 5859 21335
rect 14197 21301 14231 21335
rect 17233 21301 17267 21335
rect 18521 21301 18555 21335
rect 20453 21301 20487 21335
rect 21097 21301 21131 21335
rect 24409 21301 24443 21335
rect 24593 21301 24627 21335
rect 26157 21301 26191 21335
rect 30021 21301 30055 21335
rect 35633 21301 35667 21335
rect 43361 21301 43395 21335
rect 49801 21301 49835 21335
rect 51825 21301 51859 21335
rect 1409 21097 1443 21131
rect 4353 21097 4387 21131
rect 9505 21097 9539 21131
rect 10149 21097 10183 21131
rect 14105 21097 14139 21131
rect 25973 21097 26007 21131
rect 27813 21097 27847 21131
rect 30757 21097 30791 21131
rect 32781 21097 32815 21131
rect 34989 21097 35023 21131
rect 45477 21097 45511 21131
rect 48421 21097 48455 21131
rect 49617 21097 49651 21131
rect 53941 21097 53975 21131
rect 15393 21029 15427 21063
rect 17049 21029 17083 21063
rect 22201 21029 22235 21063
rect 23765 21029 23799 21063
rect 28273 21029 28307 21063
rect 28917 21029 28951 21063
rect 30113 21029 30147 21063
rect 32045 21029 32079 21063
rect 32965 21029 32999 21063
rect 52377 21029 52411 21063
rect 2881 20961 2915 20995
rect 6745 20961 6779 20995
rect 7113 20961 7147 20995
rect 18061 20961 18095 20995
rect 36921 20961 36955 20995
rect 42993 20961 43027 20995
rect 48789 20961 48823 20995
rect 51089 20961 51123 20995
rect 54125 20961 54159 20995
rect 57897 20961 57931 20995
rect 2513 20893 2547 20927
rect 2697 20893 2731 20927
rect 4261 20893 4295 20927
rect 4445 20893 4479 20927
rect 4813 20893 4847 20927
rect 6653 20893 6687 20927
rect 9965 20893 9999 20927
rect 10793 20893 10827 20927
rect 13277 20893 13311 20927
rect 14841 20893 14875 20927
rect 15209 20893 15243 20927
rect 15853 20893 15887 20927
rect 15946 20893 15980 20927
rect 16221 20893 16255 20927
rect 16318 20893 16352 20927
rect 18429 20893 18463 20927
rect 18521 20893 18555 20927
rect 19257 20893 19291 20927
rect 19405 20893 19439 20927
rect 19722 20893 19756 20927
rect 20545 20893 20579 20927
rect 20729 20893 20763 20927
rect 20913 20893 20947 20927
rect 21557 20893 21591 20927
rect 21677 20893 21711 20927
rect 21833 20893 21867 20927
rect 22022 20893 22056 20927
rect 24409 20893 24443 20927
rect 24685 20893 24719 20927
rect 25697 20893 25731 20927
rect 26617 20893 26651 20927
rect 27261 20893 27295 20927
rect 27537 20893 27571 20927
rect 27629 20893 27663 20927
rect 29561 20893 29595 20927
rect 29653 20893 29687 20927
rect 29837 20893 29871 20927
rect 29929 20893 29963 20927
rect 30757 20893 30791 20927
rect 30849 20893 30883 20927
rect 31585 20893 31619 20927
rect 31769 20893 31803 20927
rect 32137 20893 32171 20927
rect 34989 20893 35023 20927
rect 37013 20893 37047 20927
rect 40325 20893 40359 20927
rect 41981 20893 42015 20927
rect 42165 20893 42199 20927
rect 43453 20893 43487 20927
rect 43637 20893 43671 20927
rect 43913 20893 43947 20927
rect 45017 20893 45051 20927
rect 45293 20893 45327 20927
rect 48329 20893 48363 20927
rect 49249 20893 49283 20927
rect 49433 20893 49467 20927
rect 51365 20893 51399 20927
rect 52009 20893 52043 20927
rect 53849 20893 53883 20927
rect 54217 20893 54251 20927
rect 55689 20893 55723 20927
rect 56379 20893 56413 20927
rect 56517 20893 56551 20927
rect 56792 20893 56826 20927
rect 56885 20893 56919 20927
rect 58173 20893 58207 20927
rect 13093 20825 13127 20859
rect 15025 20825 15059 20859
rect 15117 20825 15151 20859
rect 16129 20825 16163 20859
rect 18153 20825 18187 20859
rect 19533 20825 19567 20859
rect 19625 20825 19659 20859
rect 20821 20825 20855 20859
rect 21925 20825 21959 20859
rect 25973 20825 26007 20859
rect 27445 20825 27479 20859
rect 32597 20825 32631 20859
rect 34713 20825 34747 20859
rect 34897 20825 34931 20859
rect 40509 20825 40543 20859
rect 44005 20825 44039 20859
rect 54309 20825 54343 20859
rect 55505 20825 55539 20859
rect 56609 20825 56643 20859
rect 4629 20757 4663 20791
rect 6469 20757 6503 20791
rect 10885 20757 10919 20791
rect 16497 20757 16531 20791
rect 18705 20757 18739 20791
rect 19901 20757 19935 20791
rect 21097 20757 21131 20791
rect 25789 20757 25823 20791
rect 26709 20757 26743 20791
rect 31125 20757 31159 20791
rect 32781 20757 32815 20791
rect 37381 20757 37415 20791
rect 45109 20757 45143 20791
rect 56241 20757 56275 20791
rect 3065 20553 3099 20587
rect 5273 20553 5307 20587
rect 7941 20553 7975 20587
rect 14657 20553 14691 20587
rect 18061 20553 18095 20587
rect 18613 20553 18647 20587
rect 21833 20553 21867 20587
rect 24133 20553 24167 20587
rect 26985 20553 27019 20587
rect 29193 20553 29227 20587
rect 31217 20553 31251 20587
rect 33977 20553 34011 20587
rect 34529 20553 34563 20587
rect 40877 20553 40911 20587
rect 43729 20553 43763 20587
rect 51825 20553 51859 20587
rect 57161 20553 57195 20587
rect 2329 20485 2363 20519
rect 10425 20485 10459 20519
rect 13461 20485 13495 20519
rect 25329 20485 25363 20519
rect 26065 20485 26099 20519
rect 27721 20485 27755 20519
rect 28825 20485 28859 20519
rect 29025 20485 29059 20519
rect 32965 20485 32999 20519
rect 33609 20485 33643 20519
rect 39221 20485 39255 20519
rect 42441 20485 42475 20519
rect 44925 20485 44959 20519
rect 57253 20485 57287 20519
rect 58173 20485 58207 20519
rect 2145 20417 2179 20451
rect 2513 20417 2547 20451
rect 4077 20417 4111 20451
rect 4261 20417 4295 20451
rect 7849 20417 7883 20451
rect 8125 20417 8159 20451
rect 9689 20417 9723 20451
rect 9965 20417 9999 20451
rect 13277 20417 13311 20451
rect 13369 20417 13403 20451
rect 13579 20417 13613 20451
rect 13737 20417 13771 20451
rect 18521 20417 18555 20451
rect 18705 20417 18739 20451
rect 19533 20417 19567 20451
rect 20269 20417 20303 20451
rect 29653 20417 29687 20451
rect 29837 20417 29871 20451
rect 29929 20417 29963 20451
rect 30941 20417 30975 20451
rect 33517 20417 33551 20451
rect 33793 20417 33827 20451
rect 34437 20417 34471 20451
rect 34713 20417 34747 20451
rect 38393 20417 38427 20451
rect 40509 20417 40543 20451
rect 43361 20417 43395 20451
rect 44189 20417 44223 20451
rect 45109 20417 45143 20451
rect 45201 20417 45235 20451
rect 51181 20417 51215 20451
rect 51365 20417 51399 20451
rect 51457 20417 51491 20451
rect 51549 20417 51583 20451
rect 56977 20417 57011 20451
rect 3985 20349 4019 20383
rect 4169 20349 4203 20383
rect 30389 20349 30423 20383
rect 31217 20349 31251 20383
rect 38485 20349 38519 20383
rect 40417 20349 40451 20383
rect 43453 20349 43487 20383
rect 8125 20281 8159 20315
rect 9781 20281 9815 20315
rect 13093 20281 13127 20315
rect 19349 20281 19383 20315
rect 29653 20281 29687 20315
rect 34897 20281 34931 20315
rect 42717 20281 42751 20315
rect 45201 20281 45235 20315
rect 4445 20213 4479 20247
rect 15761 20213 15795 20247
rect 20085 20213 20119 20247
rect 25973 20213 26007 20247
rect 27813 20213 27847 20247
rect 29009 20213 29043 20247
rect 31033 20213 31067 20247
rect 39773 20213 39807 20247
rect 42901 20213 42935 20247
rect 43545 20213 43579 20247
rect 56793 20213 56827 20247
rect 4721 20009 4755 20043
rect 5365 20009 5399 20043
rect 8217 20009 8251 20043
rect 13553 20009 13587 20043
rect 15393 20009 15427 20043
rect 26617 20009 26651 20043
rect 34161 20009 34195 20043
rect 43177 20009 43211 20043
rect 53941 20009 53975 20043
rect 54401 20009 54435 20043
rect 7205 19941 7239 19975
rect 11437 19941 11471 19975
rect 16313 19941 16347 19975
rect 27445 19941 27479 19975
rect 5733 19873 5767 19907
rect 11161 19873 11195 19907
rect 11989 19873 12023 19907
rect 16497 19873 16531 19907
rect 19349 19873 19383 19907
rect 30849 19873 30883 19907
rect 38301 19873 38335 19907
rect 38669 19873 38703 19907
rect 46765 19873 46799 19907
rect 47593 19873 47627 19907
rect 56793 19873 56827 19907
rect 3249 19805 3283 19839
rect 4445 19805 4479 19839
rect 5549 19805 5583 19839
rect 7113 19805 7147 19839
rect 7389 19805 7423 19839
rect 9689 19805 9723 19839
rect 11069 19805 11103 19839
rect 14105 19805 14139 19839
rect 14289 19805 14323 19839
rect 17049 19805 17083 19839
rect 19625 19805 19659 19839
rect 27169 19805 27203 19839
rect 28089 19805 28123 19839
rect 28273 19805 28307 19839
rect 28457 19805 28491 19839
rect 28917 19805 28951 19839
rect 33885 19805 33919 19839
rect 34161 19805 34195 19839
rect 34989 19805 35023 19839
rect 36001 19805 36035 19839
rect 36185 19805 36219 19839
rect 37013 19805 37047 19839
rect 38485 19805 38519 19839
rect 50169 19805 50203 19839
rect 50537 19805 50571 19839
rect 50721 19805 50755 19839
rect 53481 19805 53515 19839
rect 53757 19805 53791 19839
rect 54401 19805 54435 19839
rect 56701 19805 56735 19839
rect 56885 19805 56919 19839
rect 56977 19805 57011 19839
rect 2881 19737 2915 19771
rect 3065 19737 3099 19771
rect 8033 19737 8067 19771
rect 8233 19737 8267 19771
rect 9505 19737 9539 19771
rect 10057 19737 10091 19771
rect 16037 19737 16071 19771
rect 17233 19737 17267 19771
rect 23305 19737 23339 19771
rect 27261 19737 27295 19771
rect 27445 19737 27479 19771
rect 28181 19737 28215 19771
rect 32229 19737 32263 19771
rect 32413 19737 32447 19771
rect 34069 19737 34103 19771
rect 42993 19737 43027 19771
rect 54493 19737 54527 19771
rect 54677 19737 54711 19771
rect 4905 19669 4939 19703
rect 6285 19669 6319 19703
rect 7573 19669 7607 19703
rect 8401 19669 8435 19703
rect 14197 19669 14231 19703
rect 14841 19669 14875 19703
rect 21649 19669 21683 19703
rect 23213 19669 23247 19703
rect 27905 19669 27939 19703
rect 34805 19669 34839 19703
rect 42441 19669 42475 19703
rect 43193 19669 43227 19703
rect 43361 19669 43395 19703
rect 50537 19669 50571 19703
rect 53573 19669 53607 19703
rect 56517 19669 56551 19703
rect 4997 19465 5031 19499
rect 13369 19465 13403 19499
rect 17785 19465 17819 19499
rect 18797 19465 18831 19499
rect 19901 19465 19935 19499
rect 22477 19465 22511 19499
rect 24041 19465 24075 19499
rect 32689 19465 32723 19499
rect 35081 19465 35115 19499
rect 44189 19465 44223 19499
rect 50813 19465 50847 19499
rect 51549 19465 51583 19499
rect 12541 19397 12575 19431
rect 15945 19397 15979 19431
rect 18521 19397 18555 19431
rect 22109 19397 22143 19431
rect 24317 19397 24351 19431
rect 43269 19397 43303 19431
rect 47961 19397 47995 19431
rect 51365 19397 51399 19431
rect 56977 19397 57011 19431
rect 1501 19329 1535 19363
rect 3341 19329 3375 19363
rect 3709 19329 3743 19363
rect 5089 19329 5123 19363
rect 5733 19329 5767 19363
rect 7205 19329 7239 19363
rect 7481 19329 7515 19363
rect 7941 19329 7975 19363
rect 13645 19329 13679 19363
rect 13921 19329 13955 19363
rect 14657 19329 14691 19363
rect 14841 19329 14875 19363
rect 15117 19329 15151 19363
rect 15209 19329 15243 19363
rect 15485 19329 15519 19363
rect 17601 19329 17635 19363
rect 17785 19329 17819 19363
rect 18245 19329 18279 19363
rect 18429 19329 18463 19363
rect 18613 19329 18647 19363
rect 19257 19329 19291 19363
rect 19350 19329 19384 19363
rect 19533 19329 19567 19363
rect 19625 19329 19659 19363
rect 19722 19329 19756 19363
rect 21097 19329 21131 19363
rect 21839 19329 21873 19363
rect 21926 19329 21960 19363
rect 22201 19329 22235 19363
rect 22298 19329 22332 19363
rect 23213 19329 23247 19363
rect 23305 19329 23339 19363
rect 23489 19329 23523 19363
rect 23581 19329 23615 19363
rect 24225 19329 24259 19363
rect 24409 19329 24443 19363
rect 24593 19329 24627 19363
rect 28273 19329 28307 19363
rect 31401 19329 31435 19363
rect 32413 19329 32447 19363
rect 34345 19329 34379 19363
rect 38117 19329 38151 19363
rect 42993 19329 43027 19363
rect 43821 19329 43855 19363
rect 44005 19329 44039 19363
rect 45569 19329 45603 19363
rect 46581 19329 46615 19363
rect 47593 19329 47627 19363
rect 47777 19329 47811 19363
rect 48789 19329 48823 19363
rect 48973 19329 49007 19363
rect 49433 19329 49467 19363
rect 49525 19329 49559 19363
rect 49709 19329 49743 19363
rect 49801 19329 49835 19363
rect 50445 19329 50479 19363
rect 50813 19329 50847 19363
rect 54033 19329 54067 19363
rect 56793 19329 56827 19363
rect 7757 19261 7791 19295
rect 10793 19261 10827 19295
rect 13553 19261 13587 19295
rect 14013 19261 14047 19295
rect 16773 19261 16807 19295
rect 20453 19261 20487 19295
rect 27445 19261 27479 19295
rect 27997 19261 28031 19295
rect 32229 19261 32263 19295
rect 32321 19261 32355 19295
rect 32505 19261 32539 19295
rect 38025 19261 38059 19295
rect 42809 19261 42843 19295
rect 43361 19261 43395 19295
rect 50537 19261 50571 19295
rect 50721 19261 50755 19295
rect 53573 19261 53607 19295
rect 53941 19261 53975 19295
rect 7849 19193 7883 19227
rect 23029 19193 23063 19227
rect 34529 19193 34563 19227
rect 48789 19193 48823 19227
rect 49985 19193 50019 19227
rect 1777 19125 1811 19159
rect 4077 19125 4111 19159
rect 12817 19125 12851 19159
rect 21189 19125 21223 19159
rect 31493 19125 31527 19159
rect 38393 19125 38427 19159
rect 41797 19125 41831 19159
rect 51549 19125 51583 19159
rect 51733 19125 51767 19159
rect 54217 19125 54251 19159
rect 57161 19125 57195 19159
rect 1409 18921 1443 18955
rect 7481 18921 7515 18955
rect 10241 18921 10275 18955
rect 11161 18921 11195 18955
rect 18061 18921 18095 18955
rect 19625 18921 19659 18955
rect 22201 18921 22235 18955
rect 24409 18921 24443 18955
rect 29009 18921 29043 18955
rect 31033 18921 31067 18955
rect 32873 18921 32907 18955
rect 34161 18921 34195 18955
rect 42717 18921 42751 18955
rect 46029 18921 46063 18955
rect 52377 18921 52411 18955
rect 53757 18921 53791 18955
rect 5733 18853 5767 18887
rect 17417 18853 17451 18887
rect 20177 18853 20211 18887
rect 27629 18853 27663 18887
rect 36277 18853 36311 18887
rect 41797 18853 41831 18887
rect 7665 18785 7699 18819
rect 10977 18785 11011 18819
rect 11713 18785 11747 18819
rect 13553 18785 13587 18819
rect 15209 18785 15243 18819
rect 40325 18785 40359 18819
rect 40785 18785 40819 18819
rect 50813 18785 50847 18819
rect 56793 18785 56827 18819
rect 57345 18785 57379 18819
rect 2329 18717 2363 18751
rect 4261 18717 4295 18751
rect 4905 18717 4939 18751
rect 7205 18717 7239 18751
rect 7389 18717 7423 18751
rect 7573 18717 7607 18751
rect 10885 18717 10919 18751
rect 14381 18717 14415 18751
rect 14933 18717 14967 18751
rect 15301 18717 15335 18751
rect 15853 18717 15887 18751
rect 16221 18717 16255 18751
rect 18061 18717 18095 18751
rect 18245 18717 18279 18751
rect 19257 18717 19291 18751
rect 19441 18717 19475 18751
rect 21649 18717 21683 18751
rect 21925 18717 21959 18751
rect 22017 18717 22051 18751
rect 24409 18717 24443 18751
rect 24593 18717 24627 18751
rect 25053 18717 25087 18751
rect 25697 18717 25731 18751
rect 26065 18717 26099 18751
rect 28089 18717 28123 18751
rect 29745 18717 29779 18751
rect 29929 18717 29963 18751
rect 30113 18717 30147 18751
rect 31033 18717 31067 18751
rect 31217 18717 31251 18751
rect 31861 18717 31895 18751
rect 33609 18717 33643 18751
rect 33701 18717 33735 18751
rect 33885 18717 33919 18751
rect 33977 18717 34011 18751
rect 36001 18717 36035 18751
rect 40417 18717 40451 18751
rect 41705 18717 41739 18751
rect 41889 18717 41923 18751
rect 42533 18717 42567 18751
rect 45845 18717 45879 18751
rect 46029 18717 46063 18751
rect 50169 18717 50203 18751
rect 50353 18717 50387 18751
rect 50445 18717 50479 18751
rect 50537 18717 50571 18751
rect 52285 18717 52319 18751
rect 52561 18717 52595 18751
rect 52653 18717 52687 18751
rect 53205 18717 53239 18751
rect 53297 18717 53331 18751
rect 53481 18717 53515 18751
rect 53573 18717 53607 18751
rect 56609 18717 56643 18751
rect 57897 18717 57931 18751
rect 58081 18717 58115 18751
rect 2513 18649 2547 18683
rect 17141 18649 17175 18683
rect 21833 18649 21867 18683
rect 26709 18649 26743 18683
rect 28273 18649 28307 18683
rect 29837 18649 29871 18683
rect 32689 18649 32723 18683
rect 36277 18649 36311 18683
rect 42349 18649 42383 18683
rect 7941 18581 7975 18615
rect 17601 18581 17635 18615
rect 23857 18581 23891 18615
rect 29561 18581 29595 18615
rect 31769 18581 31803 18615
rect 32889 18581 32923 18615
rect 33057 18581 33091 18615
rect 36093 18581 36127 18615
rect 52745 18581 52779 18615
rect 57989 18581 58023 18615
rect 2789 18377 2823 18411
rect 6929 18377 6963 18411
rect 15669 18377 15703 18411
rect 26341 18377 26375 18411
rect 29193 18377 29227 18411
rect 32137 18377 32171 18411
rect 34529 18377 34563 18411
rect 40693 18377 40727 18411
rect 49341 18377 49375 18411
rect 53389 18377 53423 18411
rect 56701 18377 56735 18411
rect 57989 18377 58023 18411
rect 1869 18309 1903 18343
rect 14657 18309 14691 18343
rect 22937 18309 22971 18343
rect 24593 18309 24627 18343
rect 29377 18309 29411 18343
rect 39405 18309 39439 18343
rect 45753 18309 45787 18343
rect 2053 18241 2087 18275
rect 2789 18241 2823 18275
rect 3065 18241 3099 18275
rect 7021 18241 7055 18275
rect 7665 18241 7699 18275
rect 7849 18241 7883 18275
rect 8309 18241 8343 18275
rect 10977 18241 11011 18275
rect 11621 18241 11655 18275
rect 14473 18241 14507 18275
rect 14749 18241 14783 18275
rect 14841 18241 14875 18275
rect 15485 18241 15519 18275
rect 17785 18241 17819 18275
rect 19257 18241 19291 18275
rect 23673 18241 23707 18275
rect 24455 18241 24489 18275
rect 24685 18241 24719 18275
rect 24868 18241 24902 18275
rect 24961 18241 24995 18275
rect 27813 18241 27847 18275
rect 29101 18241 29135 18275
rect 30665 18241 30699 18275
rect 31401 18241 31435 18275
rect 32965 18241 32999 18275
rect 34345 18241 34379 18275
rect 34621 18241 34655 18275
rect 36001 18241 36035 18275
rect 36093 18241 36127 18275
rect 36277 18241 36311 18275
rect 36369 18241 36403 18275
rect 37289 18241 37323 18275
rect 38761 18241 38795 18275
rect 40509 18241 40543 18275
rect 40693 18241 40727 18275
rect 48881 18241 48915 18275
rect 48973 18241 49007 18275
rect 49157 18241 49191 18275
rect 53481 18241 53515 18275
rect 53665 18241 53699 18275
rect 56609 18241 56643 18275
rect 56793 18241 56827 18275
rect 57897 18241 57931 18275
rect 58081 18241 58115 18275
rect 8585 18173 8619 18207
rect 12633 18173 12667 18207
rect 17601 18173 17635 18207
rect 18981 18173 19015 18207
rect 19717 18173 19751 18207
rect 19993 18173 20027 18207
rect 25421 18173 25455 18207
rect 27537 18173 27571 18207
rect 29929 18173 29963 18207
rect 30389 18173 30423 18207
rect 30849 18173 30883 18207
rect 38485 18173 38519 18207
rect 44925 18173 44959 18207
rect 17969 18105 18003 18139
rect 29377 18105 29411 18139
rect 34345 18105 34379 18139
rect 36553 18105 36587 18139
rect 2237 18037 2271 18071
rect 13093 18037 13127 18071
rect 15025 18037 15059 18071
rect 23581 18037 23615 18071
rect 24317 18037 24351 18071
rect 26985 18037 27019 18071
rect 30481 18037 30515 18071
rect 31493 18037 31527 18071
rect 37473 18037 37507 18071
rect 53205 18037 53239 18071
rect 2697 17833 2731 17867
rect 7021 17833 7055 17867
rect 7665 17833 7699 17867
rect 8033 17833 8067 17867
rect 21925 17833 21959 17867
rect 24961 17833 24995 17867
rect 27629 17833 27663 17867
rect 31861 17833 31895 17867
rect 33057 17833 33091 17867
rect 33425 17833 33459 17867
rect 36185 17833 36219 17867
rect 45109 17833 45143 17867
rect 48421 17833 48455 17867
rect 53573 17833 53607 17867
rect 56977 17833 57011 17867
rect 7205 17765 7239 17799
rect 36369 17765 36403 17799
rect 41337 17765 41371 17799
rect 6193 17697 6227 17731
rect 12449 17697 12483 17731
rect 17601 17697 17635 17731
rect 19717 17697 19751 17731
rect 26985 17697 27019 17731
rect 40877 17697 40911 17731
rect 44281 17697 44315 17731
rect 44465 17697 44499 17731
rect 45477 17697 45511 17731
rect 53665 17697 53699 17731
rect 57069 17697 57103 17731
rect 4997 17629 5031 17663
rect 5181 17629 5215 17663
rect 5825 17629 5859 17663
rect 6009 17629 6043 17663
rect 7665 17629 7699 17663
rect 7849 17629 7883 17663
rect 8953 17629 8987 17663
rect 9137 17629 9171 17663
rect 12633 17629 12667 17663
rect 14289 17629 14323 17663
rect 15209 17629 15243 17663
rect 17785 17629 17819 17663
rect 19533 17629 19567 17663
rect 20177 17629 20211 17663
rect 20270 17629 20304 17663
rect 20642 17629 20676 17663
rect 22661 17629 22695 17663
rect 23305 17629 23339 17663
rect 23673 17629 23707 17663
rect 24409 17629 24443 17663
rect 24777 17629 24811 17663
rect 25881 17629 25915 17663
rect 27169 17629 27203 17663
rect 28181 17629 28215 17663
rect 28825 17629 28859 17663
rect 30021 17629 30055 17663
rect 30665 17629 30699 17663
rect 32321 17629 32355 17663
rect 33057 17629 33091 17663
rect 33241 17629 33275 17663
rect 40969 17629 41003 17663
rect 44189 17629 44223 17663
rect 45017 17629 45051 17663
rect 48237 17629 48271 17663
rect 49341 17629 49375 17663
rect 49433 17629 49467 17663
rect 53941 17629 53975 17663
rect 56793 17629 56827 17663
rect 56885 17629 56919 17663
rect 58081 17629 58115 17663
rect 2421 17561 2455 17595
rect 5365 17561 5399 17595
rect 6837 17561 6871 17595
rect 7053 17561 7087 17595
rect 15025 17561 15059 17595
rect 15577 17561 15611 17595
rect 20453 17561 20487 17595
rect 20545 17561 20579 17595
rect 22017 17561 22051 17595
rect 23489 17561 23523 17595
rect 23581 17561 23615 17595
rect 24593 17561 24627 17595
rect 24685 17561 24719 17595
rect 27261 17561 27295 17595
rect 30205 17561 30239 17595
rect 33885 17561 33919 17595
rect 36001 17561 36035 17595
rect 36217 17561 36251 17595
rect 36921 17561 36955 17595
rect 44465 17561 44499 17595
rect 48329 17561 48363 17595
rect 48513 17561 48547 17595
rect 57713 17561 57747 17595
rect 8953 17493 8987 17527
rect 12817 17493 12851 17527
rect 14473 17493 14507 17527
rect 18337 17493 18371 17527
rect 20821 17493 20855 17527
rect 22753 17493 22787 17527
rect 23857 17493 23891 17527
rect 26341 17493 26375 17527
rect 28273 17493 28307 17527
rect 30849 17493 30883 17527
rect 32505 17493 32539 17527
rect 40233 17493 40267 17527
rect 48973 17493 49007 17527
rect 49617 17493 49651 17527
rect 53389 17493 53423 17527
rect 3341 17289 3375 17323
rect 8335 17289 8369 17323
rect 20085 17289 20119 17323
rect 45661 17289 45695 17323
rect 52929 17289 52963 17323
rect 58081 17289 58115 17323
rect 7481 17221 7515 17255
rect 7665 17221 7699 17255
rect 8125 17221 8159 17255
rect 9045 17221 9079 17255
rect 14289 17221 14323 17255
rect 21189 17221 21223 17255
rect 23765 17221 23799 17255
rect 24685 17221 24719 17255
rect 25973 17221 26007 17255
rect 28641 17221 28675 17255
rect 31217 17221 31251 17255
rect 31309 17221 31343 17255
rect 33425 17221 33459 17255
rect 36553 17221 36587 17255
rect 37749 17221 37783 17255
rect 57069 17221 57103 17255
rect 8953 17153 8987 17187
rect 9137 17153 9171 17187
rect 9965 17153 9999 17187
rect 10241 17153 10275 17187
rect 10793 17153 10827 17187
rect 14105 17153 14139 17187
rect 14381 17153 14415 17187
rect 14473 17153 14507 17187
rect 15117 17153 15151 17187
rect 15301 17153 15335 17187
rect 15393 17153 15427 17187
rect 15485 17153 15519 17187
rect 18245 17153 18279 17187
rect 19533 17153 19567 17187
rect 19717 17153 19751 17187
rect 19809 17153 19843 17187
rect 19901 17153 19935 17187
rect 20545 17153 20579 17187
rect 20729 17153 20763 17187
rect 28365 17153 28399 17187
rect 28549 17153 28583 17187
rect 28733 17153 28767 17187
rect 31033 17153 31067 17187
rect 31401 17153 31435 17187
rect 32505 17153 32539 17187
rect 33241 17153 33275 17187
rect 33517 17153 33551 17187
rect 33609 17153 33643 17187
rect 34345 17153 34379 17187
rect 36001 17153 36035 17187
rect 37473 17153 37507 17187
rect 37841 17153 37875 17187
rect 40785 17153 40819 17187
rect 45293 17153 45327 17187
rect 45385 17153 45419 17187
rect 48145 17153 48179 17187
rect 49157 17153 49191 17187
rect 49341 17153 49375 17187
rect 50445 17153 50479 17187
rect 50813 17153 50847 17187
rect 51273 17153 51307 17187
rect 52745 17153 52779 17187
rect 53021 17153 53055 17187
rect 53665 17153 53699 17187
rect 54033 17153 54067 17187
rect 2881 17085 2915 17119
rect 7297 17085 7331 17119
rect 13645 17085 13679 17119
rect 37289 17085 37323 17119
rect 40693 17085 40727 17119
rect 48053 17085 48087 17119
rect 48513 17085 48547 17119
rect 48973 17085 49007 17119
rect 50261 17085 50295 17119
rect 51365 17085 51399 17119
rect 53481 17085 53515 17119
rect 56517 17085 56551 17119
rect 3249 17017 3283 17051
rect 10885 17017 10919 17051
rect 18061 17017 18095 17051
rect 23581 17017 23615 17051
rect 26157 17017 26191 17051
rect 41153 17017 41187 17051
rect 52745 17017 52779 17051
rect 53941 17017 53975 17051
rect 1685 16949 1719 16983
rect 8309 16949 8343 16983
rect 8493 16949 8527 16983
rect 14657 16949 14691 16983
rect 15669 16949 15703 16983
rect 20545 16949 20579 16983
rect 24593 16949 24627 16983
rect 28917 16949 28951 16983
rect 30021 16949 30055 16983
rect 31585 16949 31619 16983
rect 32689 16949 32723 16983
rect 33793 16949 33827 16983
rect 36645 16949 36679 16983
rect 40049 16949 40083 16983
rect 45293 16949 45327 16983
rect 50721 16949 50755 16983
rect 51273 16949 51307 16983
rect 51641 16949 51675 16983
rect 1961 16745 1995 16779
rect 7849 16745 7883 16779
rect 10425 16745 10459 16779
rect 12909 16745 12943 16779
rect 13461 16745 13495 16779
rect 15577 16745 15611 16779
rect 46305 16745 46339 16779
rect 50169 16745 50203 16779
rect 51089 16745 51123 16779
rect 52193 16745 52227 16779
rect 53665 16745 53699 16779
rect 54125 16745 54159 16779
rect 54309 16745 54343 16779
rect 2881 16677 2915 16711
rect 5825 16677 5859 16711
rect 9505 16677 9539 16711
rect 11989 16677 12023 16711
rect 12817 16677 12851 16711
rect 20729 16677 20763 16711
rect 23857 16677 23891 16711
rect 24869 16677 24903 16711
rect 27077 16677 27111 16711
rect 39037 16677 39071 16711
rect 44005 16677 44039 16711
rect 47133 16677 47167 16711
rect 3249 16609 3283 16643
rect 16865 16609 16899 16643
rect 19717 16609 19751 16643
rect 28365 16609 28399 16643
rect 30849 16609 30883 16643
rect 31401 16609 31435 16643
rect 33241 16609 33275 16643
rect 34713 16609 34747 16643
rect 35265 16609 35299 16643
rect 36185 16609 36219 16643
rect 37105 16609 37139 16643
rect 38761 16609 38795 16643
rect 46029 16609 46063 16643
rect 57161 16609 57195 16643
rect 4169 16541 4203 16575
rect 4629 16541 4663 16575
rect 7757 16541 7791 16575
rect 7941 16541 7975 16575
rect 9413 16541 9447 16575
rect 9505 16541 9539 16575
rect 14197 16541 14231 16575
rect 14565 16541 14599 16575
rect 15485 16541 15519 16575
rect 19901 16541 19935 16575
rect 19993 16541 20027 16575
rect 20177 16541 20211 16575
rect 20269 16541 20303 16575
rect 20913 16541 20947 16575
rect 21281 16541 21315 16575
rect 23581 16541 23615 16575
rect 23857 16541 23891 16575
rect 24409 16541 24443 16575
rect 24501 16541 24535 16575
rect 24685 16541 24719 16575
rect 26433 16541 26467 16575
rect 26526 16541 26560 16575
rect 26801 16541 26835 16575
rect 26939 16541 26973 16575
rect 28089 16541 28123 16575
rect 31033 16541 31067 16575
rect 32965 16541 32999 16575
rect 35081 16541 35115 16575
rect 36277 16541 36311 16575
rect 38669 16541 38703 16575
rect 43177 16541 43211 16575
rect 43729 16541 43763 16575
rect 44005 16541 44039 16575
rect 45937 16541 45971 16575
rect 46765 16541 46799 16575
rect 46949 16541 46983 16575
rect 51825 16541 51859 16575
rect 52009 16541 52043 16575
rect 53205 16541 53239 16575
rect 53481 16541 53515 16575
rect 56241 16541 56275 16575
rect 56425 16541 56459 16575
rect 58173 16541 58207 16575
rect 1869 16473 1903 16507
rect 7297 16473 7331 16507
rect 9229 16473 9263 16507
rect 10241 16473 10275 16507
rect 10425 16473 10459 16507
rect 12449 16473 12483 16507
rect 14381 16473 14415 16507
rect 14473 16473 14507 16507
rect 15301 16473 15335 16507
rect 21005 16473 21039 16507
rect 21097 16473 21131 16507
rect 26709 16473 26743 16507
rect 31309 16473 31343 16507
rect 42901 16473 42935 16507
rect 43085 16473 43119 16507
rect 54493 16473 54527 16507
rect 57897 16473 57931 16507
rect 2789 16405 2823 16439
rect 10609 16405 10643 16439
rect 14749 16405 14783 16439
rect 16313 16405 16347 16439
rect 23673 16405 23707 16439
rect 25881 16405 25915 16439
rect 29745 16405 29779 16439
rect 31861 16405 31895 16439
rect 35081 16405 35115 16439
rect 42349 16405 42383 16439
rect 43177 16405 43211 16439
rect 43821 16405 43855 16439
rect 53297 16405 53331 16439
rect 54283 16405 54317 16439
rect 1777 16201 1811 16235
rect 3709 16201 3743 16235
rect 8217 16201 8251 16235
rect 9137 16201 9171 16235
rect 13553 16201 13587 16235
rect 23673 16201 23707 16235
rect 27169 16201 27203 16235
rect 32505 16201 32539 16235
rect 34621 16201 34655 16235
rect 36645 16201 36679 16235
rect 53021 16201 53055 16235
rect 58173 16201 58207 16235
rect 3341 16133 3375 16167
rect 9505 16133 9539 16167
rect 13001 16133 13035 16167
rect 14289 16133 14323 16167
rect 19901 16133 19935 16167
rect 26341 16133 26375 16167
rect 27537 16133 27571 16167
rect 28457 16133 28491 16167
rect 29193 16133 29227 16167
rect 36277 16133 36311 16167
rect 2421 16065 2455 16099
rect 3249 16065 3283 16099
rect 3525 16065 3559 16099
rect 7205 16065 7239 16099
rect 7573 16065 7607 16099
rect 8033 16065 8067 16099
rect 9045 16065 9079 16099
rect 9321 16065 9355 16099
rect 9965 16065 9999 16099
rect 10517 16065 10551 16099
rect 12899 16065 12933 16099
rect 13093 16065 13127 16099
rect 15945 16065 15979 16099
rect 16129 16065 16163 16099
rect 17141 16065 17175 16099
rect 19625 16065 19659 16099
rect 19718 16065 19752 16099
rect 19993 16065 20027 16099
rect 20131 16065 20165 16099
rect 23029 16065 23063 16099
rect 23122 16065 23156 16099
rect 23305 16065 23339 16099
rect 23397 16065 23431 16099
rect 23494 16065 23528 16099
rect 24225 16065 24259 16099
rect 27353 16065 27387 16099
rect 27445 16065 27479 16099
rect 27721 16065 27755 16099
rect 28273 16065 28307 16099
rect 28917 16065 28951 16099
rect 29009 16065 29043 16099
rect 30021 16065 30055 16099
rect 30297 16065 30331 16099
rect 33149 16065 33183 16099
rect 36093 16065 36127 16099
rect 36369 16065 36403 16099
rect 36507 16065 36541 16099
rect 38669 16065 38703 16099
rect 42809 16065 42843 16099
rect 43085 16065 43119 16099
rect 44281 16065 44315 16099
rect 44373 16065 44407 16099
rect 52745 16065 52779 16099
rect 56241 16065 56275 16099
rect 56517 16065 56551 16099
rect 56609 16065 56643 16099
rect 2513 15997 2547 16031
rect 10333 15997 10367 16031
rect 14473 15997 14507 16031
rect 30481 15997 30515 16031
rect 34161 15997 34195 16031
rect 38577 15997 38611 16031
rect 39497 15997 39531 16031
rect 44189 15997 44223 16031
rect 44465 15997 44499 16031
rect 53021 15997 53055 16031
rect 2789 15929 2823 15963
rect 20269 15929 20303 15963
rect 22477 15929 22511 15963
rect 25789 15929 25823 15963
rect 29193 15929 29227 15963
rect 15209 15861 15243 15895
rect 16129 15861 16163 15895
rect 17233 15861 17267 15895
rect 19073 15861 19107 15895
rect 24777 15861 24811 15895
rect 30113 15861 30147 15895
rect 44649 15861 44683 15895
rect 52837 15861 52871 15895
rect 56333 15861 56367 15895
rect 56793 15861 56827 15895
rect 3065 15657 3099 15691
rect 10057 15657 10091 15691
rect 14473 15657 14507 15691
rect 19809 15657 19843 15691
rect 22845 15657 22879 15691
rect 26801 15657 26835 15691
rect 29837 15657 29871 15691
rect 31033 15657 31067 15691
rect 39865 15657 39899 15691
rect 44097 15657 44131 15691
rect 46581 15657 46615 15691
rect 46765 15657 46799 15691
rect 52929 15657 52963 15691
rect 53113 15657 53147 15691
rect 7849 15589 7883 15623
rect 13553 15589 13587 15623
rect 24409 15589 24443 15623
rect 40969 15589 41003 15623
rect 50445 15589 50479 15623
rect 11345 15521 11379 15555
rect 11897 15521 11931 15555
rect 40509 15521 40543 15555
rect 47317 15521 47351 15555
rect 47777 15521 47811 15555
rect 53573 15521 53607 15555
rect 56793 15521 56827 15555
rect 57713 15521 57747 15555
rect 3801 15453 3835 15487
rect 3985 15453 4019 15487
rect 6929 15453 6963 15487
rect 7389 15453 7423 15487
rect 7757 15453 7791 15487
rect 9505 15453 9539 15487
rect 9597 15453 9631 15487
rect 9781 15453 9815 15487
rect 9873 15453 9907 15487
rect 10609 15453 10643 15487
rect 10793 15453 10827 15487
rect 14197 15453 14231 15487
rect 14289 15453 14323 15487
rect 15117 15453 15151 15487
rect 15393 15453 15427 15487
rect 16405 15453 16439 15487
rect 16553 15453 16587 15487
rect 16911 15453 16945 15487
rect 19257 15453 19291 15487
rect 19441 15453 19475 15487
rect 19625 15453 19659 15487
rect 20453 15453 20487 15487
rect 21373 15453 21407 15487
rect 23029 15453 23063 15487
rect 23397 15453 23431 15487
rect 24593 15453 24627 15487
rect 24777 15453 24811 15487
rect 24961 15453 24995 15487
rect 26065 15453 26099 15487
rect 32137 15453 32171 15487
rect 32505 15453 32539 15487
rect 40601 15453 40635 15487
rect 41981 15453 42015 15487
rect 42533 15453 42567 15487
rect 42809 15453 42843 15487
rect 46305 15453 46339 15487
rect 47409 15453 47443 15487
rect 50169 15453 50203 15487
rect 52745 15453 52779 15487
rect 52929 15453 52963 15487
rect 57069 15453 57103 15487
rect 16681 15385 16715 15419
rect 16773 15385 16807 15419
rect 19533 15385 19567 15419
rect 23121 15385 23155 15419
rect 23213 15385 23247 15419
rect 24685 15385 24719 15419
rect 26249 15385 26283 15419
rect 34069 15385 34103 15419
rect 42625 15385 42659 15419
rect 43913 15385 43947 15419
rect 50445 15385 50479 15419
rect 3893 15317 3927 15351
rect 8953 15317 8987 15351
rect 10701 15317 10735 15351
rect 17049 15317 17083 15351
rect 20361 15317 20395 15351
rect 21281 15317 21315 15351
rect 25881 15317 25915 15351
rect 31585 15317 31619 15351
rect 32137 15317 32171 15351
rect 32321 15317 32355 15351
rect 32413 15317 32447 15351
rect 32965 15317 32999 15351
rect 33517 15317 33551 15351
rect 42993 15317 43027 15351
rect 44113 15317 44147 15351
rect 44281 15317 44315 15351
rect 50261 15317 50295 15351
rect 2605 15113 2639 15147
rect 7573 15113 7607 15147
rect 9229 15113 9263 15147
rect 10885 15113 10919 15147
rect 14631 15113 14665 15147
rect 20729 15113 20763 15147
rect 29929 15113 29963 15147
rect 38393 15113 38427 15147
rect 38945 15113 38979 15147
rect 50721 15113 50755 15147
rect 56885 15113 56919 15147
rect 2145 15045 2179 15079
rect 2881 15045 2915 15079
rect 2973 15045 3007 15079
rect 3801 15045 3835 15079
rect 10057 15045 10091 15079
rect 11529 15045 11563 15079
rect 11745 15045 11779 15079
rect 14841 15045 14875 15079
rect 15761 15045 15795 15079
rect 15853 15045 15887 15079
rect 20361 15045 20395 15079
rect 24409 15045 24443 15079
rect 24501 15045 24535 15079
rect 28733 15045 28767 15079
rect 30941 15045 30975 15079
rect 49525 15045 49559 15079
rect 49893 15045 49927 15079
rect 50353 15045 50387 15079
rect 50553 15045 50587 15079
rect 54309 15045 54343 15079
rect 2789 14977 2823 15011
rect 3157 14977 3191 15011
rect 3617 14977 3651 15011
rect 3893 14977 3927 15011
rect 3990 14977 4024 15011
rect 5825 14977 5859 15011
rect 6561 14977 6595 15011
rect 7389 14977 7423 15011
rect 7665 14977 7699 15011
rect 7849 14977 7883 15011
rect 9229 14977 9263 15011
rect 9413 14977 9447 15011
rect 9873 14977 9907 15011
rect 10241 14977 10275 15011
rect 10701 14977 10735 15011
rect 12357 14977 12391 15011
rect 12449 14977 12483 15011
rect 12633 14977 12667 15011
rect 13277 14977 13311 15011
rect 13553 14977 13587 15011
rect 14013 14977 14047 15011
rect 15577 14977 15611 15011
rect 15969 14977 16003 15011
rect 17141 14977 17175 15011
rect 17601 14977 17635 15011
rect 20085 14977 20119 15011
rect 20178 14977 20212 15011
rect 20453 14977 20487 15011
rect 20569 14977 20603 15011
rect 24312 14977 24346 15011
rect 24684 14977 24718 15011
rect 24777 14977 24811 15011
rect 25881 14977 25915 15011
rect 26157 14977 26191 15011
rect 26985 14977 27019 15011
rect 27169 14977 27203 15011
rect 27629 14977 27663 15011
rect 28549 14977 28583 15011
rect 28825 14977 28859 15011
rect 28917 14977 28951 15011
rect 29929 14977 29963 15011
rect 30757 14977 30791 15011
rect 30849 14977 30883 15011
rect 31125 14977 31159 15011
rect 32322 14977 32356 15011
rect 32413 14977 32447 15011
rect 32597 14977 32631 15011
rect 33517 14977 33551 15011
rect 34345 14977 34379 15011
rect 37473 14977 37507 15011
rect 37565 14977 37599 15011
rect 37749 14977 37783 15011
rect 40969 14977 41003 15011
rect 44281 14977 44315 15011
rect 44373 14977 44407 15011
rect 44557 14977 44591 15011
rect 45201 14977 45235 15011
rect 45385 14977 45419 15011
rect 45477 14977 45511 15011
rect 46489 14977 46523 15011
rect 48697 14977 48731 15011
rect 48881 14977 48915 15011
rect 48973 14977 49007 15011
rect 49449 14967 49483 15001
rect 49709 14977 49743 15011
rect 52837 14977 52871 15011
rect 53113 14977 53147 15011
rect 53941 14977 53975 15011
rect 56793 14977 56827 15011
rect 56977 14977 57011 15011
rect 6653 14909 6687 14943
rect 6929 14909 6963 14943
rect 16773 14909 16807 14943
rect 29561 14909 29595 14943
rect 30113 14909 30147 14943
rect 32505 14909 32539 14943
rect 33333 14909 33367 14943
rect 33885 14909 33919 14943
rect 44741 14909 44775 14943
rect 46305 14909 46339 14943
rect 53757 14909 53791 14943
rect 4169 14841 4203 14875
rect 8401 14841 8435 14875
rect 12633 14841 12667 14875
rect 13369 14841 13403 14875
rect 14473 14841 14507 14875
rect 17693 14841 17727 14875
rect 19533 14841 19567 14875
rect 25973 14841 26007 14875
rect 27077 14841 27111 14875
rect 29101 14841 29135 14875
rect 33793 14841 33827 14875
rect 37933 14841 37967 14875
rect 52929 14841 52963 14875
rect 53021 14841 53055 14875
rect 4721 14773 4755 14807
rect 11713 14773 11747 14807
rect 11897 14773 11931 14807
rect 14657 14773 14691 14807
rect 16129 14773 16163 14807
rect 23581 14773 23615 14807
rect 24133 14773 24167 14807
rect 30573 14773 30607 14807
rect 32137 14773 32171 14807
rect 34437 14773 34471 14807
rect 35081 14773 35115 14807
rect 40785 14773 40819 14807
rect 45477 14773 45511 14807
rect 46673 14773 46707 14807
rect 48973 14773 49007 14807
rect 50537 14773 50571 14807
rect 53297 14773 53331 14807
rect 54217 14773 54251 14807
rect 1593 14569 1627 14603
rect 4169 14569 4203 14603
rect 6929 14569 6963 14603
rect 9781 14569 9815 14603
rect 10609 14569 10643 14603
rect 12265 14569 12299 14603
rect 13185 14569 13219 14603
rect 20453 14569 20487 14603
rect 27261 14569 27295 14603
rect 31033 14569 31067 14603
rect 33241 14569 33275 14603
rect 40049 14569 40083 14603
rect 44005 14569 44039 14603
rect 50445 14569 50479 14603
rect 53389 14569 53423 14603
rect 36553 14501 36587 14535
rect 52929 14501 52963 14535
rect 53757 14501 53791 14535
rect 7573 14433 7607 14467
rect 38301 14433 38335 14467
rect 40693 14433 40727 14467
rect 44097 14433 44131 14467
rect 53481 14433 53515 14467
rect 56701 14433 56735 14467
rect 1409 14365 1443 14399
rect 2053 14365 2087 14399
rect 10425 14365 10459 14399
rect 15761 14365 15795 14399
rect 15945 14365 15979 14399
rect 16129 14365 16163 14399
rect 16773 14365 16807 14399
rect 17233 14365 17267 14399
rect 19901 14365 19935 14399
rect 20177 14365 20211 14399
rect 20269 14365 20303 14399
rect 21005 14365 21039 14399
rect 21189 14365 21223 14399
rect 24961 14365 24995 14399
rect 28181 14365 28215 14399
rect 28549 14365 28583 14399
rect 29837 14365 29871 14399
rect 29929 14365 29963 14399
rect 30205 14365 30239 14399
rect 32045 14365 32079 14399
rect 32137 14365 32171 14399
rect 32321 14365 32355 14399
rect 33517 14365 33551 14399
rect 34989 14365 35023 14399
rect 35173 14365 35207 14399
rect 35633 14365 35667 14399
rect 36001 14365 36035 14399
rect 36369 14365 36403 14399
rect 37749 14365 37783 14399
rect 38025 14365 38059 14399
rect 38393 14365 38427 14399
rect 40785 14365 40819 14399
rect 44005 14365 44039 14399
rect 45845 14365 45879 14399
rect 45937 14365 45971 14399
rect 46121 14365 46155 14399
rect 50169 14365 50203 14399
rect 50261 14365 50295 14399
rect 50445 14365 50479 14399
rect 53389 14365 53423 14399
rect 54493 14365 54527 14399
rect 54585 14365 54619 14399
rect 54769 14365 54803 14399
rect 55781 14365 55815 14399
rect 55965 14365 55999 14399
rect 57897 14365 57931 14399
rect 3801 14297 3835 14331
rect 3985 14297 4019 14331
rect 6837 14297 6871 14331
rect 16037 14297 16071 14331
rect 17509 14297 17543 14331
rect 20085 14297 20119 14331
rect 21741 14297 21775 14331
rect 22385 14297 22419 14331
rect 24777 14297 24811 14331
rect 28273 14297 28307 14331
rect 28365 14297 28399 14331
rect 30021 14297 30055 14331
rect 33057 14297 33091 14331
rect 33977 14297 34011 14331
rect 38853 14297 38887 14331
rect 39037 14297 39071 14331
rect 4721 14229 4755 14263
rect 15025 14229 15059 14263
rect 16313 14229 16347 14263
rect 21833 14229 21867 14263
rect 23673 14229 23707 14263
rect 27997 14229 28031 14263
rect 29653 14229 29687 14263
rect 31493 14229 31527 14263
rect 32505 14229 32539 14263
rect 33241 14229 33275 14263
rect 41153 14229 41187 14263
rect 44373 14229 44407 14263
rect 46305 14229 46339 14263
rect 58081 14229 58115 14263
rect 13737 14025 13771 14059
rect 25789 14025 25823 14059
rect 31033 14025 31067 14059
rect 32873 14025 32907 14059
rect 50445 14025 50479 14059
rect 57897 14025 57931 14059
rect 12541 13957 12575 13991
rect 14381 13957 14415 13991
rect 15761 13957 15795 13991
rect 22201 13957 22235 13991
rect 28181 13957 28215 13991
rect 31493 13957 31527 13991
rect 33333 13957 33367 13991
rect 37289 13957 37323 13991
rect 44189 13957 44223 13991
rect 56885 13957 56919 13991
rect 3433 13889 3467 13923
rect 3985 13889 4019 13923
rect 9597 13889 9631 13923
rect 10241 13889 10275 13923
rect 12725 13889 12759 13923
rect 13369 13889 13403 13923
rect 13553 13889 13587 13923
rect 15025 13889 15059 13923
rect 15577 13889 15611 13923
rect 15853 13889 15887 13923
rect 15969 13889 16003 13923
rect 16681 13889 16715 13923
rect 20177 13889 20211 13923
rect 20729 13889 20763 13923
rect 20913 13889 20947 13923
rect 21005 13889 21039 13923
rect 21097 13889 21131 13923
rect 21833 13889 21867 13923
rect 21926 13889 21960 13923
rect 22109 13889 22143 13923
rect 22339 13889 22373 13923
rect 23305 13889 23339 13923
rect 23489 13889 23523 13923
rect 24501 13889 24535 13923
rect 27997 13889 28031 13923
rect 32505 13889 32539 13923
rect 32597 13889 32631 13923
rect 34437 13889 34471 13923
rect 34989 13889 35023 13923
rect 35265 13889 35299 13923
rect 36461 13889 36495 13923
rect 37473 13889 37507 13923
rect 38209 13889 38243 13923
rect 43913 13889 43947 13923
rect 44005 13889 44039 13923
rect 53205 13889 53239 13923
rect 53849 13889 53883 13923
rect 55321 13889 55355 13923
rect 55505 13889 55539 13923
rect 56609 13889 56643 13923
rect 57897 13889 57931 13923
rect 58081 13889 58115 13923
rect 5365 13821 5399 13855
rect 8033 13821 8067 13855
rect 11529 13821 11563 13855
rect 12909 13821 12943 13855
rect 16957 13821 16991 13855
rect 24685 13821 24719 13855
rect 38117 13821 38151 13855
rect 44189 13821 44223 13855
rect 53021 13821 53055 13855
rect 56885 13821 56919 13855
rect 4629 13753 4663 13787
rect 8769 13753 8803 13787
rect 19993 13753 20027 13787
rect 21281 13753 21315 13787
rect 34253 13753 34287 13787
rect 13369 13685 13403 13719
rect 16129 13685 16163 13719
rect 22477 13685 22511 13719
rect 23121 13685 23155 13719
rect 25145 13685 25179 13719
rect 32689 13685 32723 13719
rect 36185 13685 36219 13719
rect 38485 13685 38519 13719
rect 55413 13685 55447 13719
rect 56701 13685 56735 13719
rect 7941 13481 7975 13515
rect 9689 13481 9723 13515
rect 28089 13481 28123 13515
rect 31125 13481 31159 13515
rect 53205 13481 53239 13515
rect 56793 13481 56827 13515
rect 57161 13481 57195 13515
rect 9597 13413 9631 13447
rect 10701 13413 10735 13447
rect 12357 13413 12391 13447
rect 23765 13413 23799 13447
rect 25513 13413 25547 13447
rect 29837 13413 29871 13447
rect 2237 13345 2271 13379
rect 12817 13345 12851 13379
rect 15577 13345 15611 13379
rect 23213 13345 23247 13379
rect 23305 13345 23339 13379
rect 26157 13345 26191 13379
rect 35357 13345 35391 13379
rect 36277 13345 36311 13379
rect 40693 13345 40727 13379
rect 46765 13345 46799 13379
rect 50721 13345 50755 13379
rect 56885 13345 56919 13379
rect 2973 13277 3007 13311
rect 3157 13277 3191 13311
rect 6469 13277 6503 13311
rect 7389 13277 7423 13311
rect 14565 13277 14599 13311
rect 16037 13277 16071 13311
rect 16405 13277 16439 13311
rect 17509 13277 17543 13311
rect 17693 13277 17727 13311
rect 17877 13277 17911 13311
rect 19257 13277 19291 13311
rect 19717 13277 19751 13311
rect 20637 13277 20671 13311
rect 22109 13277 22143 13311
rect 24869 13277 24903 13311
rect 24962 13277 24996 13311
rect 25237 13277 25271 13311
rect 25375 13277 25409 13311
rect 26249 13277 26283 13311
rect 27813 13277 27847 13311
rect 28089 13277 28123 13311
rect 29837 13277 29871 13311
rect 30113 13277 30147 13311
rect 32229 13277 32263 13311
rect 32505 13277 32539 13311
rect 35633 13277 35667 13311
rect 40785 13277 40819 13311
rect 42349 13277 42383 13311
rect 42533 13277 42567 13311
rect 45017 13277 45051 13311
rect 45109 13277 45143 13311
rect 45293 13277 45327 13311
rect 46949 13277 46983 13311
rect 48329 13277 48363 13311
rect 50813 13277 50847 13311
rect 53021 13277 53055 13311
rect 56793 13277 56827 13311
rect 9229 13209 9263 13243
rect 12817 13209 12851 13243
rect 12909 13209 12943 13243
rect 13553 13209 13587 13243
rect 15393 13209 15427 13243
rect 16221 13209 16255 13243
rect 16313 13209 16347 13243
rect 17785 13209 17819 13243
rect 19993 13209 20027 13243
rect 20453 13209 20487 13243
rect 23305 13209 23339 13243
rect 25145 13209 25179 13243
rect 32321 13209 32355 13243
rect 47685 13209 47719 13243
rect 49341 13209 49375 13243
rect 10241 13141 10275 13175
rect 11805 13141 11839 13175
rect 14749 13141 14783 13175
rect 16589 13141 16623 13175
rect 18061 13141 18095 13175
rect 22017 13141 22051 13175
rect 27077 13141 27111 13175
rect 27905 13141 27939 13175
rect 28549 13141 28583 13175
rect 30021 13141 30055 13175
rect 31769 13141 31803 13175
rect 32689 13141 32723 13175
rect 38485 13141 38519 13175
rect 41153 13141 41187 13175
rect 43361 13141 43395 13175
rect 45477 13141 45511 13175
rect 51181 13141 51215 13175
rect 53481 13141 53515 13175
rect 1593 12937 1627 12971
rect 10425 12937 10459 12971
rect 13093 12937 13127 12971
rect 14933 12937 14967 12971
rect 16957 12937 16991 12971
rect 19165 12937 19199 12971
rect 19717 12937 19751 12971
rect 23949 12937 23983 12971
rect 25053 12937 25087 12971
rect 37841 12937 37875 12971
rect 50353 12937 50387 12971
rect 54493 12937 54527 12971
rect 6377 12869 6411 12903
rect 13645 12869 13679 12903
rect 14289 12869 14323 12903
rect 18797 12869 18831 12903
rect 24685 12869 24719 12903
rect 42901 12869 42935 12903
rect 46673 12869 46707 12903
rect 47777 12869 47811 12903
rect 47869 12869 47903 12903
rect 54585 12869 54619 12903
rect 55689 12869 55723 12903
rect 1409 12801 1443 12835
rect 3157 12801 3191 12835
rect 4077 12801 4111 12835
rect 6561 12801 6595 12835
rect 6745 12801 6779 12835
rect 8585 12801 8619 12835
rect 8861 12801 8895 12835
rect 9505 12801 9539 12835
rect 9873 12801 9907 12835
rect 12081 12801 12115 12835
rect 13001 12801 13035 12835
rect 13185 12801 13219 12835
rect 15485 12801 15519 12835
rect 16681 12801 16715 12835
rect 16865 12801 16899 12835
rect 18613 12801 18647 12835
rect 18889 12801 18923 12835
rect 18981 12801 19015 12835
rect 24501 12801 24535 12835
rect 24777 12801 24811 12835
rect 24869 12801 24903 12835
rect 25605 12801 25639 12835
rect 28641 12801 28675 12835
rect 29377 12801 29411 12835
rect 30573 12801 30607 12835
rect 32137 12801 32171 12835
rect 32321 12801 32355 12835
rect 36737 12801 36771 12835
rect 37749 12801 37783 12835
rect 38025 12801 38059 12835
rect 38669 12801 38703 12835
rect 38853 12801 38887 12835
rect 38945 12801 38979 12835
rect 41337 12801 41371 12835
rect 41613 12801 41647 12835
rect 45017 12801 45051 12835
rect 45201 12801 45235 12835
rect 46581 12801 46615 12835
rect 46765 12801 46799 12835
rect 47593 12801 47627 12835
rect 47961 12801 47995 12835
rect 50813 12801 50847 12835
rect 50997 12801 51031 12835
rect 51917 12801 51951 12835
rect 54125 12801 54159 12835
rect 55045 12801 55079 12835
rect 55229 12801 55263 12835
rect 55321 12801 55355 12835
rect 55413 12801 55447 12835
rect 56333 12801 56367 12835
rect 56701 12801 56735 12835
rect 56977 12801 57011 12835
rect 2605 12733 2639 12767
rect 8401 12733 8435 12767
rect 12357 12733 12391 12767
rect 28365 12733 28399 12767
rect 29101 12733 29135 12767
rect 36461 12733 36495 12767
rect 41153 12733 41187 12767
rect 41705 12733 41739 12767
rect 42441 12733 42475 12767
rect 45109 12733 45143 12767
rect 51641 12733 51675 12767
rect 52101 12733 52135 12767
rect 54217 12733 54251 12767
rect 56517 12733 56551 12767
rect 25789 12665 25823 12699
rect 32229 12665 32263 12699
rect 42533 12665 42567 12699
rect 51089 12665 51123 12699
rect 7849 12597 7883 12631
rect 10885 12597 10919 12631
rect 18153 12597 18187 12631
rect 23029 12597 23063 12631
rect 30481 12597 30515 12631
rect 38209 12597 38243 12631
rect 38761 12597 38795 12631
rect 48145 12597 48179 12631
rect 51733 12597 51767 12631
rect 54309 12597 54343 12631
rect 3801 12393 3835 12427
rect 4169 12393 4203 12427
rect 5917 12393 5951 12427
rect 9137 12393 9171 12427
rect 14473 12393 14507 12427
rect 15945 12393 15979 12427
rect 32505 12393 32539 12427
rect 34897 12393 34931 12427
rect 37565 12393 37599 12427
rect 1409 12325 1443 12359
rect 13461 12325 13495 12359
rect 29009 12325 29043 12359
rect 30849 12325 30883 12359
rect 40417 12325 40451 12359
rect 46029 12325 46063 12359
rect 51457 12325 51491 12359
rect 8401 12257 8435 12291
rect 22201 12257 22235 12291
rect 41061 12257 41095 12291
rect 49249 12257 49283 12291
rect 51365 12257 51399 12291
rect 57897 12257 57931 12291
rect 4261 12189 4295 12223
rect 5181 12189 5215 12223
rect 5365 12189 5399 12223
rect 6096 12189 6130 12223
rect 6469 12189 6503 12223
rect 7113 12189 7147 12223
rect 8033 12189 8067 12223
rect 8217 12189 8251 12223
rect 9321 12189 9355 12223
rect 9597 12189 9631 12223
rect 12633 12189 12667 12223
rect 12817 12189 12851 12223
rect 15025 12189 15059 12223
rect 15209 12189 15243 12223
rect 16681 12189 16715 12223
rect 17049 12189 17083 12223
rect 19441 12189 19475 12223
rect 20085 12189 20119 12223
rect 20177 12189 20211 12223
rect 20361 12189 20395 12223
rect 20453 12189 20487 12223
rect 21373 12189 21407 12223
rect 21557 12189 21591 12223
rect 21741 12189 21775 12223
rect 22385 12189 22419 12223
rect 22569 12189 22603 12223
rect 22661 12189 22695 12223
rect 23121 12189 23155 12223
rect 25053 12189 25087 12223
rect 28733 12189 28767 12223
rect 28825 12189 28859 12223
rect 29745 12189 29779 12223
rect 29837 12189 29871 12223
rect 30113 12189 30147 12223
rect 30573 12189 30607 12223
rect 30849 12189 30883 12223
rect 32505 12189 32539 12223
rect 32597 12189 32631 12223
rect 38209 12189 38243 12223
rect 38301 12189 38335 12223
rect 38485 12189 38519 12223
rect 41153 12189 41187 12223
rect 45753 12189 45787 12223
rect 48605 12189 48639 12223
rect 48789 12189 48823 12223
rect 49065 12189 49099 12223
rect 51457 12189 51491 12223
rect 52101 12189 52135 12223
rect 52285 12189 52319 12223
rect 56425 12189 56459 12223
rect 57069 12189 57103 12223
rect 57253 12189 57287 12223
rect 58173 12189 58207 12223
rect 6193 12121 6227 12155
rect 6285 12121 6319 12155
rect 6929 12121 6963 12155
rect 7297 12121 7331 12155
rect 15853 12121 15887 12155
rect 16773 12121 16807 12155
rect 16865 12121 16899 12155
rect 19625 12121 19659 12155
rect 20637 12121 20671 12155
rect 21465 12121 21499 12155
rect 29009 12121 29043 12155
rect 29929 12121 29963 12155
rect 31401 12121 31435 12155
rect 34713 12121 34747 12155
rect 34913 12121 34947 12155
rect 38669 12121 38703 12155
rect 46029 12121 46063 12155
rect 51181 12121 51215 12155
rect 51917 12121 51951 12155
rect 56241 12121 56275 12155
rect 5273 12053 5307 12087
rect 9505 12053 9539 12087
rect 10149 12053 10183 12087
rect 11805 12053 11839 12087
rect 15117 12053 15151 12087
rect 16497 12053 16531 12087
rect 18521 12053 18555 12087
rect 19257 12053 19291 12087
rect 21189 12053 21223 12087
rect 25145 12053 25179 12087
rect 29561 12053 29595 12087
rect 30665 12053 30699 12087
rect 31953 12053 31987 12087
rect 32873 12053 32907 12087
rect 35081 12053 35115 12087
rect 41521 12053 41555 12087
rect 45845 12053 45879 12087
rect 56609 12053 56643 12087
rect 57069 12053 57103 12087
rect 5641 11849 5675 11883
rect 6469 11849 6503 11883
rect 8401 11849 8435 11883
rect 8953 11849 8987 11883
rect 18797 11849 18831 11883
rect 19349 11849 19383 11883
rect 19993 11849 20027 11883
rect 21925 11849 21959 11883
rect 29745 11849 29779 11883
rect 30297 11849 30331 11883
rect 32229 11849 32263 11883
rect 33809 11849 33843 11883
rect 34621 11849 34655 11883
rect 38577 11849 38611 11883
rect 45385 11849 45419 11883
rect 49065 11849 49099 11883
rect 58173 11849 58207 11883
rect 9137 11781 9171 11815
rect 21189 11781 21223 11815
rect 22753 11781 22787 11815
rect 25789 11781 25823 11815
rect 28457 11781 28491 11815
rect 30481 11781 30515 11815
rect 33609 11781 33643 11815
rect 37749 11781 37783 11815
rect 38485 11781 38519 11815
rect 38669 11781 38703 11815
rect 43729 11781 43763 11815
rect 53481 11781 53515 11815
rect 3065 11713 3099 11747
rect 3157 11713 3191 11747
rect 3341 11713 3375 11747
rect 3433 11713 3467 11747
rect 3893 11713 3927 11747
rect 4077 11713 4111 11747
rect 5641 11713 5675 11747
rect 5825 11713 5859 11747
rect 6377 11713 6411 11747
rect 6561 11713 6595 11747
rect 8309 11713 8343 11747
rect 8493 11713 8527 11747
rect 9321 11713 9355 11747
rect 11897 11713 11931 11747
rect 12357 11713 12391 11747
rect 15393 11713 15427 11747
rect 15485 11713 15519 11747
rect 15669 11713 15703 11747
rect 15761 11713 15795 11747
rect 16819 11713 16853 11747
rect 16957 11713 16991 11747
rect 17049 11713 17083 11747
rect 17233 11713 17267 11747
rect 19901 11713 19935 11747
rect 20085 11713 20119 11747
rect 22385 11713 22419 11747
rect 22478 11713 22512 11747
rect 22661 11713 22695 11747
rect 22850 11713 22884 11747
rect 23765 11713 23799 11747
rect 25605 11713 25639 11747
rect 25697 11713 25731 11747
rect 25973 11713 26007 11747
rect 28181 11713 28215 11747
rect 28365 11713 28399 11747
rect 28549 11713 28583 11747
rect 29193 11713 29227 11747
rect 29377 11713 29411 11747
rect 29469 11713 29503 11747
rect 29561 11713 29595 11747
rect 30205 11713 30239 11747
rect 34529 11713 34563 11747
rect 34805 11713 34839 11747
rect 38393 11713 38427 11747
rect 39129 11713 39163 11747
rect 43177 11713 43211 11747
rect 43453 11713 43487 11747
rect 43821 11713 43855 11747
rect 45017 11713 45051 11747
rect 46121 11713 46155 11747
rect 46213 11713 46247 11747
rect 48697 11713 48731 11747
rect 53665 11713 53699 11747
rect 56057 11713 56091 11747
rect 56701 11713 56735 11747
rect 57069 11713 57103 11747
rect 57253 11713 57287 11747
rect 3985 11645 4019 11679
rect 7849 11645 7883 11679
rect 44925 11645 44959 11679
rect 45937 11645 45971 11679
rect 46029 11645 46063 11679
rect 48789 11645 48823 11679
rect 48881 11645 48915 11679
rect 56609 11645 56643 11679
rect 7113 11577 7147 11611
rect 23581 11577 23615 11611
rect 37933 11577 37967 11611
rect 2881 11509 2915 11543
rect 9873 11509 9907 11543
rect 15209 11509 15243 11543
rect 16681 11509 16715 11543
rect 21097 11509 21131 11543
rect 23029 11509 23063 11543
rect 25421 11509 25455 11543
rect 28733 11509 28767 11543
rect 30481 11509 30515 11543
rect 33793 11509 33827 11543
rect 33977 11509 34011 11543
rect 34805 11509 34839 11543
rect 39313 11509 39347 11543
rect 46397 11509 46431 11543
rect 53297 11509 53331 11543
rect 2881 11305 2915 11339
rect 3801 11305 3835 11339
rect 22293 11305 22327 11339
rect 25329 11305 25363 11339
rect 42349 11305 42383 11339
rect 46121 11305 46155 11339
rect 47685 11305 47719 11339
rect 30665 11237 30699 11271
rect 33977 11237 34011 11271
rect 36001 11237 36035 11271
rect 39129 11237 39163 11271
rect 46305 11237 46339 11271
rect 52745 11237 52779 11271
rect 11989 11169 12023 11203
rect 15669 11169 15703 11203
rect 17601 11169 17635 11203
rect 31217 11169 31251 11203
rect 35173 11169 35207 11203
rect 40325 11169 40359 11203
rect 53297 11169 53331 11203
rect 54033 11169 54067 11203
rect 2973 11101 3007 11135
rect 3801 11101 3835 11135
rect 3985 11101 4019 11135
rect 12173 11101 12207 11135
rect 14657 11101 14691 11135
rect 14933 11101 14967 11135
rect 15853 11101 15887 11135
rect 16129 11101 16163 11135
rect 16589 11101 16623 11135
rect 16957 11101 16991 11135
rect 17785 11101 17819 11135
rect 21741 11101 21775 11135
rect 22109 11101 22143 11135
rect 22845 11101 22879 11135
rect 25329 11101 25363 11135
rect 25513 11101 25547 11135
rect 25605 11101 25639 11135
rect 27537 11101 27571 11135
rect 27813 11101 27847 11135
rect 27905 11101 27939 11135
rect 31309 11101 31343 11135
rect 31493 11101 31527 11135
rect 33701 11101 33735 11135
rect 33793 11101 33827 11135
rect 34805 11101 34839 11135
rect 34989 11101 35023 11135
rect 35265 11101 35299 11135
rect 35449 11101 35483 11135
rect 36001 11101 36035 11135
rect 36185 11101 36219 11135
rect 38577 11101 38611 11135
rect 38761 11101 38795 11135
rect 38945 11101 38979 11135
rect 42165 11101 42199 11135
rect 42349 11101 42383 11135
rect 43177 11101 43211 11135
rect 43453 11101 43487 11135
rect 43637 11101 43671 11135
rect 48237 11101 48271 11135
rect 48513 11101 48547 11135
rect 49157 11101 49191 11135
rect 49341 11101 49375 11135
rect 51733 11101 51767 11135
rect 53021 11101 53055 11135
rect 53757 11101 53791 11135
rect 56241 11101 56275 11135
rect 56425 11101 56459 11135
rect 56701 11101 56735 11135
rect 56885 11101 56919 11135
rect 57345 11101 57379 11135
rect 57529 11101 57563 11135
rect 57989 11101 58023 11135
rect 3157 11033 3191 11067
rect 14473 11033 14507 11067
rect 14841 11033 14875 11067
rect 16037 11033 16071 11067
rect 16773 11033 16807 11067
rect 16865 11033 16899 11067
rect 21925 11033 21959 11067
rect 22017 11033 22051 11067
rect 27721 11033 27755 11067
rect 31677 11033 31711 11067
rect 33977 11033 34011 11067
rect 38853 11033 38887 11067
rect 43269 11033 43303 11067
rect 45937 11033 45971 11067
rect 46137 11033 46171 11067
rect 48697 11033 48731 11067
rect 58081 11033 58115 11067
rect 9689 10965 9723 10999
rect 12357 10965 12391 10999
rect 17141 10965 17175 10999
rect 22937 10965 22971 10999
rect 28089 10965 28123 10999
rect 48329 10965 48363 10999
rect 49157 10965 49191 10999
rect 51825 10965 51859 10999
rect 57437 10965 57471 10999
rect 2513 10761 2547 10795
rect 4077 10761 4111 10795
rect 6377 10761 6411 10795
rect 9137 10761 9171 10795
rect 10057 10761 10091 10795
rect 14381 10761 14415 10795
rect 42441 10761 42475 10795
rect 47961 10761 47995 10795
rect 52745 10761 52779 10795
rect 54033 10761 54067 10795
rect 56333 10761 56367 10795
rect 11805 10693 11839 10727
rect 15117 10693 15151 10727
rect 15577 10693 15611 10727
rect 19441 10693 19475 10727
rect 23029 10693 23063 10727
rect 23121 10693 23155 10727
rect 24409 10693 24443 10727
rect 25329 10693 25363 10727
rect 26157 10693 26191 10727
rect 29653 10693 29687 10727
rect 34897 10693 34931 10727
rect 39681 10693 39715 10727
rect 39865 10693 39899 10727
rect 53113 10693 53147 10727
rect 55965 10693 55999 10727
rect 56149 10693 56183 10727
rect 1409 10625 1443 10659
rect 3341 10625 3375 10659
rect 4261 10625 4295 10659
rect 6561 10625 6595 10659
rect 9321 10625 9355 10659
rect 9965 10625 9999 10659
rect 10149 10625 10183 10659
rect 12173 10625 12207 10659
rect 12357 10625 12391 10659
rect 13001 10625 13035 10659
rect 13185 10625 13219 10659
rect 19303 10625 19337 10659
rect 19533 10625 19567 10659
rect 19716 10625 19750 10659
rect 19809 10625 19843 10659
rect 22937 10625 22971 10659
rect 23305 10625 23339 10659
rect 25145 10625 25179 10659
rect 25237 10625 25271 10659
rect 25513 10625 25547 10659
rect 27487 10625 27521 10659
rect 27905 10625 27939 10659
rect 29377 10625 29411 10659
rect 29470 10625 29504 10659
rect 29745 10625 29779 10659
rect 29883 10625 29917 10659
rect 32689 10625 32723 10659
rect 33609 10625 33643 10659
rect 35173 10625 35207 10659
rect 36645 10625 36679 10659
rect 37381 10625 37415 10659
rect 37565 10625 37599 10659
rect 38945 10625 38979 10659
rect 39221 10625 39255 10659
rect 40693 10625 40727 10659
rect 48605 10625 48639 10659
rect 48973 10625 49007 10659
rect 51733 10625 51767 10659
rect 52101 10625 52135 10659
rect 52929 10625 52963 10659
rect 53205 10625 53239 10659
rect 53665 10625 53699 10659
rect 53849 10625 53883 10659
rect 54493 10625 54527 10659
rect 54677 10625 54711 10659
rect 56977 10625 57011 10659
rect 57161 10625 57195 10659
rect 57897 10625 57931 10659
rect 3249 10557 3283 10591
rect 4445 10557 4479 10591
rect 6745 10557 6779 10591
rect 9505 10557 9539 10591
rect 10701 10557 10735 10591
rect 27353 10557 27387 10591
rect 34989 10557 35023 10591
rect 36369 10557 36403 10591
rect 38301 10557 38335 10591
rect 40601 10557 40635 10591
rect 49525 10557 49559 10591
rect 51641 10557 51675 10591
rect 1593 10489 1627 10523
rect 22753 10489 22787 10523
rect 27813 10489 27847 10523
rect 30021 10489 30055 10523
rect 38945 10489 38979 10523
rect 11897 10421 11931 10455
rect 12817 10421 12851 10455
rect 13001 10421 13035 10455
rect 18613 10421 18647 10455
rect 19165 10421 19199 10455
rect 24317 10421 24351 10455
rect 24961 10421 24995 10455
rect 26065 10421 26099 10455
rect 30849 10421 30883 10455
rect 32137 10421 32171 10455
rect 35173 10421 35207 10455
rect 35357 10421 35391 10455
rect 39957 10421 39991 10455
rect 40969 10421 41003 10455
rect 54585 10421 54619 10455
rect 56793 10421 56827 10455
rect 58081 10421 58115 10455
rect 1409 10217 1443 10251
rect 5825 10217 5859 10251
rect 6653 10217 6687 10251
rect 6837 10217 6871 10251
rect 9413 10217 9447 10251
rect 12265 10217 12299 10251
rect 36369 10217 36403 10251
rect 38761 10217 38795 10251
rect 39865 10217 39899 10251
rect 53481 10217 53515 10251
rect 55689 10217 55723 10251
rect 5917 10149 5951 10183
rect 19257 10149 19291 10183
rect 20913 10149 20947 10183
rect 29929 10149 29963 10183
rect 38945 10149 38979 10183
rect 5733 10081 5767 10115
rect 9045 10081 9079 10115
rect 12633 10081 12667 10115
rect 15025 10081 15059 10115
rect 21741 10081 21775 10115
rect 26249 10081 26283 10115
rect 28181 10081 28215 10115
rect 43177 10081 43211 10115
rect 45569 10081 45603 10115
rect 46029 10081 46063 10115
rect 48513 10081 48547 10115
rect 49249 10081 49283 10115
rect 49525 10081 49559 10115
rect 55597 10081 55631 10115
rect 55781 10081 55815 10115
rect 2973 10013 3007 10047
rect 3157 10013 3191 10047
rect 3801 10013 3835 10047
rect 3985 10013 4019 10047
rect 6009 10013 6043 10047
rect 6469 10013 6503 10047
rect 6653 10013 6687 10047
rect 9137 10013 9171 10047
rect 12449 10013 12483 10047
rect 14933 10013 14967 10047
rect 15669 10013 15703 10047
rect 15945 10013 15979 10047
rect 16589 10013 16623 10047
rect 16773 10013 16807 10047
rect 17049 10013 17083 10047
rect 19257 10013 19291 10047
rect 19441 10013 19475 10047
rect 21649 10013 21683 10047
rect 21833 10013 21867 10047
rect 22569 10013 22603 10047
rect 22661 10013 22695 10047
rect 22845 10013 22879 10047
rect 22937 10013 22971 10047
rect 26525 10013 26559 10047
rect 28457 10013 28491 10047
rect 30113 10013 30147 10047
rect 32689 10013 32723 10047
rect 33057 10013 33091 10047
rect 36185 10013 36219 10047
rect 36553 10013 36587 10047
rect 40969 10013 41003 10047
rect 41153 10013 41187 10047
rect 41245 10013 41279 10047
rect 41889 10013 41923 10047
rect 42165 10013 42199 10047
rect 42625 10013 42659 10047
rect 42809 10013 42843 10047
rect 45661 10013 45695 10047
rect 47777 10013 47811 10047
rect 48145 10013 48179 10047
rect 49157 10013 49191 10047
rect 51549 10013 51583 10047
rect 55873 10013 55907 10047
rect 56793 10013 56827 10047
rect 56977 10013 57011 10047
rect 21097 9945 21131 9979
rect 32137 9945 32171 9979
rect 38577 9945 38611 9979
rect 38777 9945 38811 9979
rect 51181 9945 51215 9979
rect 51733 9945 51767 9979
rect 3065 9877 3099 9911
rect 3893 9877 3927 9911
rect 9965 9877 9999 9911
rect 14105 9877 14139 9911
rect 15761 9877 15795 9911
rect 16129 9877 16163 9911
rect 16957 9877 16991 9911
rect 22385 9877 22419 9911
rect 24593 9877 24627 9911
rect 33701 9877 33735 9911
rect 35633 9877 35667 9911
rect 36737 9877 36771 9911
rect 41245 9877 41279 9911
rect 41705 9877 41739 9911
rect 42073 9877 42107 9911
rect 43085 9877 43119 9911
rect 57161 9877 57195 9911
rect 57713 9877 57747 9911
rect 6377 9673 6411 9707
rect 15301 9673 15335 9707
rect 25329 9673 25363 9707
rect 28595 9673 28629 9707
rect 35357 9673 35391 9707
rect 36093 9673 36127 9707
rect 43085 9673 43119 9707
rect 55229 9673 55263 9707
rect 8677 9605 8711 9639
rect 9597 9605 9631 9639
rect 17969 9605 18003 9639
rect 22937 9605 22971 9639
rect 23857 9605 23891 9639
rect 23949 9605 23983 9639
rect 25605 9605 25639 9639
rect 27445 9605 27479 9639
rect 29929 9605 29963 9639
rect 30021 9605 30055 9639
rect 42717 9605 42751 9639
rect 42922 9605 42956 9639
rect 44005 9605 44039 9639
rect 44189 9605 44223 9639
rect 3157 9537 3191 9571
rect 3433 9537 3467 9571
rect 3709 9537 3743 9571
rect 3801 9537 3835 9571
rect 4077 9537 4111 9571
rect 6745 9537 6779 9571
rect 8861 9537 8895 9571
rect 9045 9537 9079 9571
rect 11529 9537 11563 9571
rect 11713 9537 11747 9571
rect 12633 9537 12667 9571
rect 13093 9537 13127 9571
rect 18889 9537 18923 9571
rect 18981 9537 19015 9571
rect 19165 9537 19199 9571
rect 19257 9537 19291 9571
rect 20361 9537 20395 9571
rect 20453 9537 20487 9571
rect 20637 9537 20671 9571
rect 20729 9537 20763 9571
rect 22707 9537 22741 9571
rect 22821 9537 22855 9571
rect 23121 9537 23155 9571
rect 23719 9537 23753 9571
rect 24133 9537 24167 9571
rect 24685 9537 24719 9571
rect 24869 9537 24903 9571
rect 25513 9537 25547 9571
rect 25697 9537 25731 9571
rect 25881 9537 25915 9571
rect 28825 9537 28859 9571
rect 29653 9537 29687 9571
rect 29801 9537 29835 9571
rect 30118 9537 30152 9571
rect 36001 9537 36035 9571
rect 36369 9537 36403 9571
rect 41705 9537 41739 9571
rect 41889 9537 41923 9571
rect 44833 9537 44867 9571
rect 45477 9537 45511 9571
rect 45845 9537 45879 9571
rect 46029 9537 46063 9571
rect 54033 9537 54067 9571
rect 55137 9537 55171 9571
rect 55321 9537 55355 9571
rect 6653 9469 6687 9503
rect 36553 9469 36587 9503
rect 55873 9469 55907 9503
rect 56333 9469 56367 9503
rect 18153 9401 18187 9435
rect 23581 9401 23615 9435
rect 44925 9401 44959 9435
rect 55137 9401 55171 9435
rect 56057 9401 56091 9435
rect 4445 9333 4479 9367
rect 11621 9333 11655 9367
rect 15853 9333 15887 9367
rect 18705 9333 18739 9367
rect 20177 9333 20211 9367
rect 22569 9333 22603 9367
rect 24869 9333 24903 9367
rect 30297 9333 30331 9367
rect 41797 9333 41831 9367
rect 42901 9333 42935 9367
rect 44373 9333 44407 9367
rect 54309 9333 54343 9367
rect 54493 9333 54527 9367
rect 3249 9129 3283 9163
rect 4169 9129 4203 9163
rect 6561 9129 6595 9163
rect 8217 9129 8251 9163
rect 8953 9129 8987 9163
rect 20361 9129 20395 9163
rect 29009 9129 29043 9163
rect 30573 9129 30607 9163
rect 37473 9129 37507 9163
rect 42901 9129 42935 9163
rect 54401 9129 54435 9163
rect 10517 9061 10551 9095
rect 24409 9061 24443 9095
rect 27813 9061 27847 9095
rect 32781 9061 32815 9095
rect 33333 9061 33367 9095
rect 36737 9061 36771 9095
rect 36921 9061 36955 9095
rect 9413 8993 9447 9027
rect 10977 8993 11011 9027
rect 15117 8993 15151 9027
rect 17509 8993 17543 9027
rect 32321 8993 32355 9027
rect 36461 8993 36495 9027
rect 37841 8993 37875 9027
rect 45109 8993 45143 9027
rect 45845 8993 45879 9027
rect 49157 8993 49191 9027
rect 51825 8993 51859 9027
rect 52101 8993 52135 9027
rect 57161 8993 57195 9027
rect 2881 8925 2915 8959
rect 6377 8925 6411 8959
rect 6561 8925 6595 8959
rect 8217 8925 8251 8959
rect 8401 8925 8435 8959
rect 9321 8925 9355 8959
rect 10885 8925 10919 8959
rect 15025 8925 15059 8959
rect 16773 8925 16807 8959
rect 17417 8925 17451 8959
rect 19349 8925 19383 8959
rect 19533 8925 19567 8959
rect 20177 8925 20211 8959
rect 20361 8925 20395 8959
rect 20821 8925 20855 8959
rect 22477 8925 22511 8959
rect 22569 8925 22603 8959
rect 22753 8925 22787 8959
rect 22845 8925 22879 8959
rect 24961 8925 24995 8959
rect 25237 8925 25271 8959
rect 26249 8925 26283 8959
rect 26617 8925 26651 8959
rect 27261 8925 27295 8959
rect 27353 8925 27387 8959
rect 27537 8925 27571 8959
rect 27629 8925 27663 8959
rect 28457 8925 28491 8959
rect 28641 8925 28675 8959
rect 28825 8925 28859 8959
rect 29561 8925 29595 8959
rect 29829 8925 29863 8959
rect 29929 8925 29963 8959
rect 30849 8925 30883 8959
rect 32413 8925 32447 8959
rect 34805 8925 34839 8959
rect 35817 8925 35851 8959
rect 37657 8925 37691 8959
rect 40509 8925 40543 8959
rect 41061 8925 41095 8959
rect 49249 8925 49283 8959
rect 51733 8925 51767 8959
rect 54309 8925 54343 8959
rect 54493 8925 54527 8959
rect 56241 8925 56275 8959
rect 56425 8925 56459 8959
rect 3065 8857 3099 8891
rect 3801 8857 3835 8891
rect 3985 8857 4019 8891
rect 10057 8857 10091 8891
rect 15853 8857 15887 8891
rect 19441 8857 19475 8891
rect 26433 8857 26467 8891
rect 26525 8857 26559 8891
rect 28729 8857 28763 8891
rect 29745 8857 29779 8891
rect 30573 8857 30607 8891
rect 30757 8857 30791 8891
rect 14197 8789 14231 8823
rect 17785 8789 17819 8823
rect 23029 8789 23063 8823
rect 26801 8789 26835 8823
rect 30113 8789 30147 8823
rect 38945 8789 38979 8823
rect 49617 8789 49651 8823
rect 2237 8585 2271 8619
rect 8585 8585 8619 8619
rect 17693 8585 17727 8619
rect 18337 8585 18371 8619
rect 21097 8585 21131 8619
rect 29469 8585 29503 8619
rect 31401 8585 31435 8619
rect 34805 8585 34839 8619
rect 39129 8585 39163 8619
rect 48605 8585 48639 8619
rect 51549 8585 51583 8619
rect 53849 8585 53883 8619
rect 25053 8517 25087 8551
rect 28641 8517 28675 8551
rect 28733 8517 28767 8551
rect 36277 8517 36311 8551
rect 40233 8517 40267 8551
rect 1685 8449 1719 8483
rect 2881 8449 2915 8483
rect 4445 8449 4479 8483
rect 4629 8449 4663 8483
rect 6561 8449 6595 8483
rect 6837 8449 6871 8483
rect 7021 8449 7055 8483
rect 19165 8449 19199 8483
rect 25421 8449 25455 8483
rect 28457 8449 28491 8483
rect 28825 8449 28859 8483
rect 34437 8449 34471 8483
rect 34621 8449 34655 8483
rect 37565 8449 37599 8483
rect 37933 8449 37967 8483
rect 39313 8449 39347 8483
rect 39405 8449 39439 8483
rect 39589 8449 39623 8483
rect 40141 8449 40175 8483
rect 40325 8449 40359 8483
rect 42625 8449 42659 8483
rect 46029 8449 46063 8483
rect 48602 8449 48636 8483
rect 48973 8449 49007 8483
rect 49065 8449 49099 8483
rect 51457 8449 51491 8483
rect 51641 8449 51675 8483
rect 52837 8449 52871 8483
rect 53021 8449 53055 8483
rect 54493 8449 54527 8483
rect 57069 8449 57103 8483
rect 2697 8381 2731 8415
rect 3525 8381 3559 8415
rect 3985 8381 4019 8415
rect 6377 8381 6411 8415
rect 24501 8381 24535 8415
rect 25145 8381 25179 8415
rect 25513 8381 25547 8415
rect 38577 8381 38611 8415
rect 42533 8381 42567 8415
rect 45937 8381 45971 8415
rect 54585 8381 54619 8415
rect 56241 8381 56275 8415
rect 57161 8381 57195 8415
rect 1501 8313 1535 8347
rect 3065 8313 3099 8347
rect 3709 8313 3743 8347
rect 4445 8313 4479 8347
rect 29009 8313 29043 8347
rect 39497 8313 39531 8347
rect 42993 8313 43027 8347
rect 46397 8313 46431 8347
rect 48421 8313 48455 8347
rect 54861 8313 54895 8347
rect 11805 8245 11839 8279
rect 25697 8245 25731 8279
rect 3801 8041 3835 8075
rect 6745 8041 6779 8075
rect 7665 8041 7699 8075
rect 10885 8041 10919 8075
rect 28825 8041 28859 8075
rect 35725 8041 35759 8075
rect 3985 7973 4019 8007
rect 6929 7973 6963 8007
rect 7849 7973 7883 8007
rect 10333 7973 10367 8007
rect 27813 7973 27847 8007
rect 45661 7973 45695 8007
rect 48881 7973 48915 8007
rect 52101 7973 52135 8007
rect 7205 7905 7239 7939
rect 10977 7905 11011 7939
rect 14105 7905 14139 7939
rect 17325 7905 17359 7939
rect 20177 7905 20211 7939
rect 21373 7905 21407 7939
rect 22385 7905 22419 7939
rect 30205 7905 30239 7939
rect 31585 7905 31619 7939
rect 32137 7905 32171 7939
rect 34713 7905 34747 7939
rect 40969 7905 41003 7939
rect 48421 7905 48455 7939
rect 10514 7837 10548 7871
rect 11437 7837 11471 7871
rect 11621 7837 11655 7871
rect 12081 7837 12115 7871
rect 14473 7837 14507 7871
rect 14933 7837 14967 7871
rect 16405 7837 16439 7871
rect 17233 7837 17267 7871
rect 18153 7837 18187 7871
rect 20269 7837 20303 7871
rect 21189 7837 21223 7871
rect 22661 7837 22695 7871
rect 27353 7837 27387 7871
rect 27629 7837 27663 7871
rect 28273 7837 28307 7871
rect 28457 7837 28491 7871
rect 28641 7837 28675 7871
rect 30665 7837 30699 7871
rect 30757 7837 30791 7871
rect 30941 7837 30975 7871
rect 31953 7837 31987 7871
rect 33425 7837 33459 7871
rect 33885 7837 33919 7871
rect 34069 7837 34103 7871
rect 35725 7837 35759 7871
rect 35909 7837 35943 7871
rect 39129 7837 39163 7871
rect 39313 7837 39347 7871
rect 39957 7837 39991 7871
rect 40141 7837 40175 7871
rect 41705 7837 41739 7871
rect 41889 7837 41923 7871
rect 42349 7837 42383 7871
rect 42533 7837 42567 7871
rect 42809 7837 42843 7871
rect 45569 7837 45603 7871
rect 45937 7837 45971 7871
rect 46305 7837 46339 7871
rect 48513 7837 48547 7871
rect 51641 7837 51675 7871
rect 51917 7837 51951 7871
rect 52285 7837 52319 7871
rect 52377 7837 52411 7871
rect 58081 7837 58115 7871
rect 4261 7769 4295 7803
rect 8125 7769 8159 7803
rect 23305 7769 23339 7803
rect 27445 7769 27479 7803
rect 28549 7769 28583 7803
rect 31125 7769 31159 7803
rect 39221 7769 39255 7803
rect 57529 7769 57563 7803
rect 10517 7701 10551 7735
rect 11529 7701 11563 7735
rect 18061 7701 18095 7735
rect 19901 7701 19935 7735
rect 23857 7701 23891 7735
rect 31953 7701 31987 7735
rect 33977 7701 34011 7735
rect 36093 7701 36127 7735
rect 41797 7701 41831 7735
rect 42993 7701 43027 7735
rect 10793 7497 10827 7531
rect 11529 7497 11563 7531
rect 20637 7497 20671 7531
rect 27813 7497 27847 7531
rect 31493 7497 31527 7531
rect 33977 7497 34011 7531
rect 46029 7497 46063 7531
rect 58081 7497 58115 7531
rect 14289 7429 14323 7463
rect 22845 7429 22879 7463
rect 36093 7429 36127 7463
rect 52193 7429 52227 7463
rect 6745 7361 6779 7395
rect 10425 7361 10459 7395
rect 13093 7361 13127 7395
rect 16865 7361 16899 7395
rect 17693 7361 17727 7395
rect 18705 7361 18739 7395
rect 22753 7361 22787 7395
rect 23029 7361 23063 7395
rect 23765 7361 23799 7395
rect 24685 7361 24719 7395
rect 27169 7361 27203 7395
rect 27353 7361 27387 7395
rect 27997 7361 28031 7395
rect 28089 7361 28123 7395
rect 28181 7361 28215 7395
rect 28365 7361 28399 7395
rect 28825 7361 28859 7395
rect 29009 7361 29043 7395
rect 30665 7361 30699 7395
rect 33149 7361 33183 7395
rect 34713 7361 34747 7395
rect 34897 7361 34931 7395
rect 35725 7361 35759 7395
rect 38669 7361 38703 7395
rect 42625 7361 42659 7395
rect 45017 7361 45051 7395
rect 45201 7361 45235 7395
rect 56977 7361 57011 7395
rect 6377 7293 6411 7327
rect 6837 7293 6871 7327
rect 10517 7293 10551 7327
rect 13369 7293 13403 7327
rect 17049 7293 17083 7327
rect 17877 7293 17911 7327
rect 18613 7293 18647 7327
rect 30573 7293 30607 7327
rect 33241 7293 33275 7327
rect 35633 7293 35667 7327
rect 39681 7293 39715 7327
rect 43637 7293 43671 7327
rect 51365 7293 51399 7327
rect 57069 7293 57103 7327
rect 57345 7293 57379 7327
rect 14013 7225 14047 7259
rect 19073 7225 19107 7259
rect 26157 7225 26191 7259
rect 31033 7225 31067 7259
rect 34713 7225 34747 7259
rect 35725 7225 35759 7259
rect 12909 7157 12943 7191
rect 13277 7157 13311 7191
rect 13829 7157 13863 7191
rect 16681 7157 16715 7191
rect 17509 7157 17543 7191
rect 23213 7157 23247 7191
rect 25237 7157 25271 7191
rect 27261 7157 27295 7191
rect 28917 7157 28951 7191
rect 32321 7157 32355 7191
rect 38485 7157 38519 7191
rect 55781 7157 55815 7191
rect 9597 6953 9631 6987
rect 10609 6953 10643 6987
rect 11345 6953 11379 6987
rect 17417 6953 17451 6987
rect 26985 6953 27019 6987
rect 36001 6953 36035 6987
rect 45569 6953 45603 6987
rect 48697 6953 48731 6987
rect 14197 6885 14231 6919
rect 19993 6885 20027 6919
rect 40141 6885 40175 6919
rect 48053 6885 48087 6919
rect 10057 6817 10091 6851
rect 14381 6817 14415 6851
rect 16589 6817 16623 6851
rect 16773 6817 16807 6851
rect 19809 6817 19843 6851
rect 20269 6817 20303 6851
rect 39221 6817 39255 6851
rect 47777 6817 47811 6851
rect 48237 6817 48271 6851
rect 54677 6817 54711 6851
rect 55413 6817 55447 6851
rect 57253 6817 57287 6851
rect 57805 6817 57839 6851
rect 9965 6749 9999 6783
rect 10609 6749 10643 6783
rect 10793 6749 10827 6783
rect 13277 6749 13311 6783
rect 14105 6749 14139 6783
rect 16865 6749 16899 6783
rect 24593 6749 24627 6783
rect 25237 6749 25271 6783
rect 31125 6749 31159 6783
rect 31309 6749 31343 6783
rect 35541 6749 35575 6783
rect 35817 6749 35851 6783
rect 39865 6749 39899 6783
rect 45385 6749 45419 6783
rect 48881 6749 48915 6783
rect 49157 6749 49191 6783
rect 54585 6749 54619 6783
rect 54769 6749 54803 6783
rect 55505 6749 55539 6783
rect 55965 6749 55999 6783
rect 56057 6749 56091 6783
rect 56241 6749 56275 6783
rect 56793 6749 56827 6783
rect 13093 6681 13127 6715
rect 13461 6681 13495 6715
rect 26433 6681 26467 6715
rect 38025 6681 38059 6715
rect 38669 6681 38703 6715
rect 40141 6681 40175 6715
rect 45201 6681 45235 6715
rect 14105 6613 14139 6647
rect 16589 6613 16623 6647
rect 27629 6613 27663 6647
rect 31217 6613 31251 6647
rect 35633 6613 35667 6647
rect 38117 6613 38151 6647
rect 39957 6613 39991 6647
rect 49065 6613 49099 6647
rect 6837 6409 6871 6443
rect 10517 6409 10551 6443
rect 12817 6409 12851 6443
rect 24041 6409 24075 6443
rect 27721 6409 27755 6443
rect 38853 6409 38887 6443
rect 54769 6409 54803 6443
rect 56885 6409 56919 6443
rect 57253 6409 57287 6443
rect 12173 6341 12207 6375
rect 24501 6341 24535 6375
rect 35541 6341 35575 6375
rect 43545 6341 43579 6375
rect 1869 6273 1903 6307
rect 3433 6273 3467 6307
rect 4077 6273 4111 6307
rect 7205 6273 7239 6307
rect 10057 6273 10091 6307
rect 10149 6273 10183 6307
rect 10520 6273 10554 6307
rect 12725 6273 12759 6307
rect 12909 6273 12943 6307
rect 13461 6273 13495 6307
rect 13645 6273 13679 6307
rect 16681 6273 16715 6307
rect 16865 6273 16899 6307
rect 17509 6273 17543 6307
rect 17693 6273 17727 6307
rect 20269 6273 20303 6307
rect 26341 6273 26375 6307
rect 31401 6273 31435 6307
rect 31493 6273 31527 6307
rect 36185 6273 36219 6307
rect 36369 6273 36403 6307
rect 37381 6273 37415 6307
rect 37473 6273 37507 6307
rect 39681 6273 39715 6307
rect 39957 6273 39991 6307
rect 47685 6273 47719 6307
rect 47961 6273 47995 6307
rect 48697 6273 48731 6307
rect 49341 6273 49375 6307
rect 50353 6273 50387 6307
rect 53941 6273 53975 6307
rect 55045 6273 55079 6307
rect 55413 6273 55447 6307
rect 56149 6273 56183 6307
rect 56793 6273 56827 6307
rect 57069 6273 57103 6307
rect 57897 6273 57931 6307
rect 7297 6205 7331 6239
rect 8309 6205 8343 6239
rect 19993 6205 20027 6239
rect 20821 6205 20855 6239
rect 27537 6205 27571 6239
rect 27629 6205 27663 6239
rect 40417 6205 40451 6239
rect 54033 6205 54067 6239
rect 54953 6205 54987 6239
rect 55321 6205 55355 6239
rect 55965 6205 55999 6239
rect 56333 6205 56367 6239
rect 2053 6137 2087 6171
rect 8033 6137 8067 6171
rect 10701 6137 10735 6171
rect 24225 6137 24259 6171
rect 28089 6137 28123 6171
rect 43821 6137 43855 6171
rect 54309 6137 54343 6171
rect 58081 6137 58115 6171
rect 7849 6069 7883 6103
rect 13553 6069 13587 6103
rect 16773 6069 16807 6103
rect 17049 6069 17083 6103
rect 17693 6069 17727 6103
rect 31217 6069 31251 6103
rect 35449 6069 35483 6103
rect 37657 6069 37691 6103
rect 44005 6069 44039 6103
rect 53297 6069 53331 6103
rect 1593 5865 1627 5899
rect 10149 5865 10183 5899
rect 17693 5865 17727 5899
rect 30665 5865 30699 5899
rect 32045 5865 32079 5899
rect 54217 5865 54251 5899
rect 55505 5865 55539 5899
rect 57805 5865 57839 5899
rect 16037 5797 16071 5831
rect 19625 5797 19659 5831
rect 21189 5797 21223 5831
rect 4353 5729 4387 5763
rect 6653 5729 6687 5763
rect 7205 5729 7239 5763
rect 10517 5729 10551 5763
rect 12817 5729 12851 5763
rect 17141 5729 17175 5763
rect 20453 5729 20487 5763
rect 30481 5729 30515 5763
rect 32137 5729 32171 5763
rect 36001 5729 36035 5763
rect 37105 5729 37139 5763
rect 40141 5729 40175 5763
rect 41061 5729 41095 5763
rect 43453 5729 43487 5763
rect 56977 5729 57011 5763
rect 5089 5661 5123 5695
rect 5273 5661 5307 5695
rect 6837 5661 6871 5695
rect 10425 5661 10459 5695
rect 12909 5661 12943 5695
rect 14289 5661 14323 5695
rect 16129 5661 16163 5695
rect 16313 5661 16347 5695
rect 16957 5661 16991 5695
rect 17601 5661 17635 5695
rect 17785 5661 17819 5695
rect 19901 5661 19935 5695
rect 20361 5661 20395 5695
rect 20545 5661 20579 5695
rect 21005 5661 21039 5695
rect 21189 5661 21223 5695
rect 23305 5661 23339 5695
rect 23489 5661 23523 5695
rect 24409 5661 24443 5695
rect 26985 5661 27019 5695
rect 27353 5661 27387 5695
rect 30757 5661 30791 5695
rect 31217 5661 31251 5695
rect 31401 5661 31435 5695
rect 32045 5661 32079 5695
rect 33425 5661 33459 5695
rect 33609 5661 33643 5695
rect 37013 5661 37047 5695
rect 37197 5661 37231 5695
rect 37657 5661 37691 5695
rect 37841 5661 37875 5695
rect 40049 5661 40083 5695
rect 40325 5661 40359 5695
rect 40969 5661 41003 5695
rect 43545 5661 43579 5695
rect 54125 5661 54159 5695
rect 56057 5661 56091 5695
rect 7113 5593 7147 5627
rect 14105 5593 14139 5627
rect 16773 5593 16807 5627
rect 19625 5593 19659 5627
rect 21649 5593 21683 5627
rect 24593 5593 24627 5627
rect 27077 5593 27111 5627
rect 27169 5593 27203 5627
rect 35449 5593 35483 5627
rect 41245 5593 41279 5627
rect 13277 5525 13311 5559
rect 14473 5525 14507 5559
rect 19809 5525 19843 5559
rect 23397 5525 23431 5559
rect 24777 5525 24811 5559
rect 26801 5525 26835 5559
rect 30481 5525 30515 5559
rect 31585 5525 31619 5559
rect 32413 5525 32447 5559
rect 33241 5525 33275 5559
rect 37749 5525 37783 5559
rect 40509 5525 40543 5559
rect 40969 5525 41003 5559
rect 43913 5525 43947 5559
rect 53573 5525 53607 5559
rect 3157 5321 3191 5355
rect 13277 5321 13311 5355
rect 22569 5321 22603 5355
rect 27353 5321 27387 5355
rect 56333 5321 56367 5355
rect 4077 5253 4111 5287
rect 6837 5253 6871 5287
rect 19717 5253 19751 5287
rect 19933 5253 19967 5287
rect 24133 5253 24167 5287
rect 2973 5185 3007 5219
rect 3249 5185 3283 5219
rect 3709 5185 3743 5219
rect 3802 5185 3836 5219
rect 3985 5185 4019 5219
rect 4215 5185 4249 5219
rect 9321 5185 9355 5219
rect 9505 5185 9539 5219
rect 13461 5185 13495 5219
rect 13645 5185 13679 5219
rect 16865 5185 16899 5219
rect 17601 5185 17635 5219
rect 22937 5185 22971 5219
rect 23949 5185 23983 5219
rect 24041 5185 24075 5219
rect 24271 5185 24305 5219
rect 25237 5185 25271 5219
rect 27721 5185 27755 5219
rect 31217 5185 31251 5219
rect 31401 5185 31435 5219
rect 33885 5185 33919 5219
rect 40693 5185 40727 5219
rect 40877 5185 40911 5219
rect 44189 5185 44223 5219
rect 44281 5185 44315 5219
rect 44465 5185 44499 5219
rect 45201 5185 45235 5219
rect 56977 5185 57011 5219
rect 17141 5117 17175 5151
rect 17877 5117 17911 5151
rect 23029 5117 23063 5151
rect 24409 5117 24443 5151
rect 25329 5117 25363 5151
rect 27629 5117 27663 5151
rect 32873 5117 32907 5151
rect 44373 5117 44407 5151
rect 45109 5117 45143 5151
rect 57069 5117 57103 5151
rect 4353 5049 4387 5083
rect 6561 5049 6595 5083
rect 17049 5049 17083 5083
rect 17693 5049 17727 5083
rect 24869 5049 24903 5083
rect 45569 5049 45603 5083
rect 6377 4981 6411 5015
rect 9505 4981 9539 5015
rect 16681 4981 16715 5015
rect 17601 4981 17635 5015
rect 19901 4981 19935 5015
rect 20085 4981 20119 5015
rect 23765 4981 23799 5015
rect 31585 4981 31619 5015
rect 40877 4981 40911 5015
rect 44005 4981 44039 5015
rect 54585 4981 54619 5015
rect 57345 4981 57379 5015
rect 3985 4777 4019 4811
rect 6653 4777 6687 4811
rect 7297 4777 7331 4811
rect 16221 4777 16255 4811
rect 19441 4777 19475 4811
rect 27077 4777 27111 4811
rect 33609 4777 33643 4811
rect 45109 4777 45143 4811
rect 2237 4709 2271 4743
rect 6285 4641 6319 4675
rect 10057 4641 10091 4675
rect 10241 4641 10275 4675
rect 24409 4641 24443 4675
rect 27261 4641 27295 4675
rect 29745 4641 29779 4675
rect 37749 4641 37783 4675
rect 40325 4641 40359 4675
rect 46213 4641 46247 4675
rect 46489 4641 46523 4675
rect 1685 4573 1719 4607
rect 2421 4573 2455 4607
rect 3801 4573 3835 4607
rect 3985 4573 4019 4607
rect 6469 4573 6503 4607
rect 7197 4583 7231 4617
rect 9781 4573 9815 4607
rect 10333 4573 10367 4607
rect 11069 4573 11103 4607
rect 16037 4573 16071 4607
rect 16221 4573 16255 4607
rect 19809 4573 19843 4607
rect 24593 4573 24627 4607
rect 27353 4573 27387 4607
rect 30757 4573 30791 4607
rect 33182 4573 33216 4607
rect 33701 4573 33735 4607
rect 36737 4573 36771 4607
rect 37657 4573 37691 4607
rect 37841 4573 37875 4607
rect 40417 4573 40451 4607
rect 41429 4573 41463 4607
rect 41521 4573 41555 4607
rect 45017 4573 45051 4607
rect 45201 4573 45235 4607
rect 46581 4573 46615 4607
rect 2973 4505 3007 4539
rect 19625 4505 19659 4539
rect 36921 4505 36955 4539
rect 37105 4505 37139 4539
rect 1501 4437 1535 4471
rect 11161 4437 11195 4471
rect 24777 4437 24811 4471
rect 33057 4437 33091 4471
rect 33241 4437 33275 4471
rect 40785 4437 40819 4471
rect 41245 4437 41279 4471
rect 45937 4233 45971 4267
rect 6561 4165 6595 4199
rect 6745 4165 6779 4199
rect 12817 4165 12851 4199
rect 24041 4165 24075 4199
rect 45109 4165 45143 4199
rect 45293 4165 45327 4199
rect 46305 4165 46339 4199
rect 6377 4097 6411 4131
rect 9689 4097 9723 4131
rect 12541 4097 12575 4131
rect 15945 4097 15979 4131
rect 16129 4097 16163 4131
rect 16681 4097 16715 4131
rect 16865 4097 16899 4131
rect 20545 4097 20579 4131
rect 20729 4097 20763 4131
rect 23857 4097 23891 4131
rect 33517 4097 33551 4131
rect 33701 4097 33735 4131
rect 36277 4097 36311 4131
rect 36461 4097 36495 4131
rect 37657 4097 37691 4131
rect 40416 4097 40450 4131
rect 40509 4097 40543 4131
rect 41337 4097 41371 4131
rect 41521 4097 41555 4131
rect 46121 4097 46155 4131
rect 46213 4097 46247 4131
rect 46489 4097 46523 4131
rect 9781 4029 9815 4063
rect 10425 4029 10459 4063
rect 12357 4029 12391 4063
rect 12909 4029 12943 4063
rect 17049 4029 17083 4063
rect 20913 4029 20947 4063
rect 36645 4029 36679 4063
rect 37565 4029 37599 4063
rect 40601 4029 40635 4063
rect 40693 4029 40727 4063
rect 40877 4029 40911 4063
rect 15945 3961 15979 3995
rect 11805 3893 11839 3927
rect 13461 3893 13495 3927
rect 14657 3893 14691 3927
rect 23673 3893 23707 3927
rect 33517 3893 33551 3927
rect 37381 3893 37415 3927
rect 41337 3893 41371 3927
rect 44925 3893 44959 3927
rect 58081 3893 58115 3927
rect 9689 3689 9723 3723
rect 12633 3689 12667 3723
rect 15669 3689 15703 3723
rect 57805 3689 57839 3723
rect 15117 3621 15151 3655
rect 37657 3621 37691 3655
rect 41613 3621 41647 3655
rect 42073 3621 42107 3655
rect 14473 3553 14507 3587
rect 24777 3553 24811 3587
rect 28917 3553 28951 3587
rect 31953 3553 31987 3587
rect 32873 3553 32907 3587
rect 33517 3553 33551 3587
rect 46213 3553 46247 3587
rect 10609 3485 10643 3519
rect 11253 3475 11287 3509
rect 11437 3485 11471 3519
rect 12817 3485 12851 3519
rect 13185 3485 13219 3519
rect 14289 3485 14323 3519
rect 14933 3485 14967 3519
rect 15117 3485 15151 3519
rect 16681 3485 16715 3519
rect 16865 3485 16899 3519
rect 17325 3485 17359 3519
rect 17418 3485 17452 3519
rect 17693 3485 17727 3519
rect 17831 3485 17865 3519
rect 19257 3485 19291 3519
rect 19441 3485 19475 3519
rect 20085 3485 20119 3519
rect 20269 3485 20303 3519
rect 21281 3485 21315 3519
rect 21649 3485 21683 3519
rect 24593 3485 24627 3519
rect 26157 3485 26191 3519
rect 26433 3485 26467 3519
rect 28825 3485 28859 3519
rect 31309 3485 31343 3519
rect 31493 3485 31527 3519
rect 32137 3485 32171 3519
rect 32229 3485 32263 3519
rect 32781 3485 32815 3519
rect 32965 3485 32999 3519
rect 33701 3485 33735 3519
rect 33885 3485 33919 3519
rect 37105 3485 37139 3519
rect 37289 3485 37323 3519
rect 37473 3485 37507 3519
rect 40049 3485 40083 3519
rect 40233 3485 40267 3519
rect 40877 3485 40911 3519
rect 41061 3485 41095 3519
rect 43177 3485 43211 3519
rect 43821 3485 43855 3519
rect 46121 3485 46155 3519
rect 58081 3485 58115 3519
rect 9873 3417 9907 3451
rect 10057 3417 10091 3451
rect 10701 3417 10735 3451
rect 12909 3417 12943 3451
rect 13001 3417 13035 3451
rect 16773 3417 16807 3451
rect 17601 3417 17635 3451
rect 18613 3417 18647 3451
rect 19901 3417 19935 3451
rect 23121 3417 23155 3451
rect 37381 3417 37415 3451
rect 40969 3417 41003 3451
rect 42257 3417 42291 3451
rect 42441 3417 42475 3451
rect 1409 3349 1443 3383
rect 11437 3349 11471 3383
rect 14105 3349 14139 3383
rect 17969 3349 18003 3383
rect 19441 3349 19475 3383
rect 24409 3349 24443 3383
rect 25973 3349 26007 3383
rect 26341 3349 26375 3383
rect 26985 3349 27019 3383
rect 27721 3349 27755 3383
rect 28457 3349 28491 3383
rect 31401 3349 31435 3383
rect 40233 3349 40267 3383
rect 43361 3349 43395 3383
rect 45753 3349 45787 3383
rect 57161 3349 57195 3383
rect 4629 3145 4663 3179
rect 11529 3145 11563 3179
rect 16681 3145 16715 3179
rect 19257 3145 19291 3179
rect 19717 3145 19751 3179
rect 23397 3145 23431 3179
rect 25881 3145 25915 3179
rect 37289 3145 37323 3179
rect 41705 3145 41739 3179
rect 42441 3145 42475 3179
rect 10885 3077 10919 3111
rect 14105 3077 14139 3111
rect 14289 3077 14323 3111
rect 17785 3077 17819 3111
rect 25329 3077 25363 3111
rect 31125 3077 31159 3111
rect 33885 3077 33919 3111
rect 34253 3077 34287 3111
rect 42609 3077 42643 3111
rect 42809 3077 42843 3111
rect 44557 3077 44591 3111
rect 1409 3009 1443 3043
rect 5457 3009 5491 3043
rect 10149 3009 10183 3043
rect 10333 3009 10367 3043
rect 11989 3009 12023 3043
rect 13093 3009 13127 3043
rect 13921 3009 13955 3043
rect 17049 3009 17083 3043
rect 17693 3009 17727 3043
rect 17877 3009 17911 3043
rect 18889 3009 18923 3043
rect 20545 3009 20579 3043
rect 20729 3009 20763 3043
rect 20821 3009 20855 3043
rect 24317 3009 24351 3043
rect 24498 3009 24532 3043
rect 25421 3009 25455 3043
rect 26249 3009 26283 3043
rect 26985 3009 27019 3043
rect 27169 3009 27203 3043
rect 27905 3009 27939 3043
rect 28365 3009 28399 3043
rect 28733 3009 28767 3043
rect 29285 3009 29319 3043
rect 29653 3009 29687 3043
rect 33057 3009 33091 3043
rect 33241 3009 33275 3043
rect 33425 3009 33459 3043
rect 34069 3009 34103 3043
rect 36553 3009 36587 3043
rect 37657 3009 37691 3043
rect 39773 3009 39807 3043
rect 40693 3009 40727 3043
rect 40877 3009 40911 3043
rect 41604 3031 41638 3065
rect 41889 3009 41923 3043
rect 43729 3009 43763 3043
rect 44925 3009 44959 3043
rect 45201 3009 45235 3043
rect 51365 3009 51399 3043
rect 52009 3009 52043 3043
rect 57897 3009 57931 3043
rect 1685 2941 1719 2975
rect 5549 2941 5583 2975
rect 9321 2941 9355 2975
rect 11897 2941 11931 2975
rect 12173 2941 12207 2975
rect 13001 2941 13035 2975
rect 16957 2941 16991 2975
rect 18797 2941 18831 2975
rect 23857 2941 23891 2975
rect 24685 2941 24719 2975
rect 26157 2941 26191 2975
rect 36645 2941 36679 2975
rect 37565 2941 37599 2975
rect 43821 2941 43855 2975
rect 44097 2941 44131 2975
rect 5089 2873 5123 2907
rect 13461 2873 13495 2907
rect 20637 2873 20671 2907
rect 21005 2873 21039 2907
rect 23581 2873 23615 2907
rect 33057 2873 33091 2907
rect 40233 2873 40267 2907
rect 51549 2873 51583 2907
rect 2329 2805 2363 2839
rect 2881 2805 2915 2839
rect 8493 2805 8527 2839
rect 21925 2805 21959 2839
rect 26985 2805 27019 2839
rect 32137 2805 32171 2839
rect 36277 2805 36311 2839
rect 39865 2805 39899 2839
rect 41061 2805 41095 2839
rect 41889 2805 41923 2839
rect 42625 2805 42659 2839
rect 56609 2805 56643 2839
rect 57253 2805 57287 2839
rect 58081 2805 58115 2839
rect 2789 2601 2823 2635
rect 22201 2601 22235 2635
rect 23765 2601 23799 2635
rect 27169 2601 27203 2635
rect 31401 2601 31435 2635
rect 33241 2601 33275 2635
rect 39957 2601 39991 2635
rect 46673 2601 46707 2635
rect 51181 2601 51215 2635
rect 56977 2601 57011 2635
rect 36369 2533 36403 2567
rect 48605 2533 48639 2567
rect 2053 2465 2087 2499
rect 8125 2465 8159 2499
rect 10057 2465 10091 2499
rect 15577 2465 15611 2499
rect 21097 2465 21131 2499
rect 25145 2465 25179 2499
rect 25973 2465 26007 2499
rect 26433 2465 26467 2499
rect 32229 2465 32263 2499
rect 34897 2465 34931 2499
rect 56149 2465 56183 2499
rect 1501 2397 1535 2431
rect 2605 2397 2639 2431
rect 4261 2397 4295 2431
rect 8401 2397 8435 2431
rect 9321 2397 9355 2431
rect 9781 2397 9815 2431
rect 11989 2397 12023 2431
rect 14105 2397 14139 2431
rect 15301 2397 15335 2431
rect 17693 2397 17727 2431
rect 18429 2397 18463 2431
rect 20821 2397 20855 2431
rect 20913 2397 20947 2431
rect 22017 2397 22051 2431
rect 23581 2397 23615 2431
rect 23765 2397 23799 2431
rect 25881 2397 25915 2431
rect 26157 2397 26191 2431
rect 26249 2397 26283 2431
rect 26985 2397 27019 2431
rect 27813 2397 27847 2431
rect 31585 2397 31619 2431
rect 32413 2397 32447 2431
rect 32597 2397 32631 2431
rect 33241 2397 33275 2431
rect 33425 2397 33459 2431
rect 34713 2397 34747 2431
rect 35725 2397 35759 2431
rect 36185 2397 36219 2431
rect 38117 2397 38151 2431
rect 40141 2397 40175 2431
rect 40233 2397 40267 2431
rect 41061 2397 41095 2431
rect 42441 2397 42475 2431
rect 43913 2397 43947 2431
rect 46121 2397 46155 2431
rect 48053 2397 48087 2431
rect 50629 2397 50663 2431
rect 52745 2397 52779 2431
rect 54677 2397 54711 2431
rect 55321 2397 55355 2431
rect 56425 2397 56459 2431
rect 57897 2397 57931 2431
rect 16681 2329 16715 2363
rect 19533 2329 19567 2363
rect 20085 2329 20119 2363
rect 23121 2329 23155 2363
rect 24869 2329 24903 2363
rect 28089 2329 28123 2363
rect 29009 2329 29043 2363
rect 30021 2329 30055 2363
rect 42717 2329 42751 2363
rect 54125 2329 54159 2363
rect 57253 2329 57287 2363
rect 4077 2261 4111 2295
rect 11805 2261 11839 2295
rect 12541 2261 12575 2295
rect 14289 2261 14323 2295
rect 18245 2261 18279 2295
rect 20177 2261 20211 2295
rect 30113 2261 30147 2295
rect 33057 2261 33091 2295
rect 34161 2261 34195 2295
rect 37565 2261 37599 2295
rect 38301 2261 38335 2295
rect 40877 2261 40911 2295
rect 41889 2261 41923 2295
rect 43361 2261 43395 2295
rect 44097 2261 44131 2295
rect 45937 2261 45971 2295
rect 47869 2261 47903 2295
rect 50445 2261 50479 2295
rect 52929 2261 52963 2295
rect 58081 2261 58115 2295
<< metal1 >>
rect 37550 37612 37556 37664
rect 37608 37652 37614 37664
rect 39114 37652 39120 37664
rect 37608 37624 39120 37652
rect 37608 37612 37614 37624
rect 39114 37612 39120 37624
rect 39172 37612 39178 37664
rect 1104 37562 58880 37584
rect 1104 37510 4214 37562
rect 4266 37510 4278 37562
rect 4330 37510 4342 37562
rect 4394 37510 4406 37562
rect 4458 37510 4470 37562
rect 4522 37510 34934 37562
rect 34986 37510 34998 37562
rect 35050 37510 35062 37562
rect 35114 37510 35126 37562
rect 35178 37510 35190 37562
rect 35242 37510 58880 37562
rect 1104 37488 58880 37510
rect 9953 37451 10011 37457
rect 9953 37417 9965 37451
rect 9999 37448 10011 37451
rect 37550 37448 37556 37460
rect 9999 37420 37556 37448
rect 9999 37417 10011 37420
rect 9953 37411 10011 37417
rect 37550 37408 37556 37420
rect 37608 37408 37614 37460
rect 37642 37408 37648 37460
rect 37700 37448 37706 37460
rect 37829 37451 37887 37457
rect 37829 37448 37841 37451
rect 37700 37420 37841 37448
rect 37700 37408 37706 37420
rect 37829 37417 37841 37420
rect 37875 37417 37887 37451
rect 37829 37411 37887 37417
rect 48590 37408 48596 37460
rect 48648 37448 48654 37460
rect 49053 37451 49111 37457
rect 49053 37448 49065 37451
rect 48648 37420 49065 37448
rect 48648 37408 48654 37420
rect 49053 37417 49065 37420
rect 49099 37417 49111 37451
rect 49053 37411 49111 37417
rect 5718 37340 5724 37392
rect 5776 37380 5782 37392
rect 12345 37383 12403 37389
rect 12345 37380 12357 37383
rect 5776 37352 12357 37380
rect 5776 37340 5782 37352
rect 12345 37349 12357 37352
rect 12391 37349 12403 37383
rect 23842 37380 23848 37392
rect 23803 37352 23848 37380
rect 12345 37343 12403 37349
rect 23842 37340 23848 37352
rect 23900 37340 23906 37392
rect 46750 37380 46756 37392
rect 37660 37352 46756 37380
rect 4433 37315 4491 37321
rect 4433 37281 4445 37315
rect 4479 37312 4491 37315
rect 4614 37312 4620 37324
rect 4479 37284 4620 37312
rect 4479 37281 4491 37284
rect 4433 37275 4491 37281
rect 4614 37272 4620 37284
rect 4672 37272 4678 37324
rect 9309 37315 9367 37321
rect 9309 37281 9321 37315
rect 9355 37312 9367 37315
rect 11885 37315 11943 37321
rect 9355 37284 9720 37312
rect 9355 37281 9367 37284
rect 9309 37275 9367 37281
rect 9692 37256 9720 37284
rect 11885 37281 11897 37315
rect 11931 37312 11943 37315
rect 12250 37312 12256 37324
rect 11931 37284 12256 37312
rect 11931 37281 11943 37284
rect 11885 37275 11943 37281
rect 12250 37272 12256 37284
rect 12308 37312 12314 37324
rect 12308 37284 12572 37312
rect 12308 37272 12314 37284
rect 1673 37247 1731 37253
rect 1673 37213 1685 37247
rect 1719 37213 1731 37247
rect 2406 37244 2412 37256
rect 2367 37216 2412 37244
rect 1673 37207 1731 37213
rect 1688 37176 1716 37207
rect 2406 37204 2412 37216
rect 2464 37244 2470 37256
rect 2869 37247 2927 37253
rect 2869 37244 2881 37247
rect 2464 37216 2881 37244
rect 2464 37204 2470 37216
rect 2869 37213 2881 37216
rect 2915 37213 2927 37247
rect 2869 37207 2927 37213
rect 3878 37204 3884 37256
rect 3936 37244 3942 37256
rect 4249 37247 4307 37253
rect 4249 37244 4261 37247
rect 3936 37216 4261 37244
rect 3936 37204 3942 37216
rect 4249 37213 4261 37216
rect 4295 37213 4307 37247
rect 4249 37207 4307 37213
rect 5810 37204 5816 37256
rect 5868 37244 5874 37256
rect 6365 37247 6423 37253
rect 6365 37244 6377 37247
rect 5868 37216 6377 37244
rect 5868 37204 5874 37216
rect 6365 37213 6377 37216
rect 6411 37213 6423 37247
rect 6365 37207 6423 37213
rect 7377 37247 7435 37253
rect 7377 37213 7389 37247
rect 7423 37244 7435 37247
rect 7742 37244 7748 37256
rect 7423 37216 7748 37244
rect 7423 37213 7435 37216
rect 7377 37207 7435 37213
rect 7742 37204 7748 37216
rect 7800 37244 7806 37256
rect 7837 37247 7895 37253
rect 7837 37244 7849 37247
rect 7800 37216 7849 37244
rect 7800 37204 7806 37216
rect 7837 37213 7849 37216
rect 7883 37213 7895 37247
rect 7837 37207 7895 37213
rect 9674 37204 9680 37256
rect 9732 37244 9738 37256
rect 12544 37253 12572 37284
rect 14182 37272 14188 37324
rect 14240 37312 14246 37324
rect 14277 37315 14335 37321
rect 14277 37312 14289 37315
rect 14240 37284 14289 37312
rect 14240 37272 14246 37284
rect 14277 37281 14289 37284
rect 14323 37281 14335 37315
rect 14277 37275 14335 37281
rect 16117 37315 16175 37321
rect 16117 37281 16129 37315
rect 16163 37312 16175 37315
rect 16163 37284 16712 37312
rect 16163 37281 16175 37284
rect 16117 37275 16175 37281
rect 16684 37256 16712 37284
rect 9861 37247 9919 37253
rect 9861 37244 9873 37247
rect 9732 37216 9873 37244
rect 9732 37204 9738 37216
rect 9861 37213 9873 37216
rect 9907 37213 9919 37247
rect 9861 37207 9919 37213
rect 12529 37247 12587 37253
rect 12529 37213 12541 37247
rect 12575 37213 12587 37247
rect 12529 37207 12587 37213
rect 14553 37247 14611 37253
rect 14553 37213 14565 37247
rect 14599 37213 14611 37247
rect 16666 37244 16672 37256
rect 16627 37216 16672 37244
rect 14553 37207 14611 37213
rect 7098 37176 7104 37188
rect 1688 37148 7104 37176
rect 7098 37136 7104 37148
rect 7156 37136 7162 37188
rect 14568 37176 14596 37207
rect 16666 37204 16672 37216
rect 16724 37204 16730 37256
rect 18417 37247 18475 37253
rect 18417 37213 18429 37247
rect 18463 37213 18475 37247
rect 18417 37207 18475 37213
rect 19613 37247 19671 37253
rect 19613 37213 19625 37247
rect 19659 37244 19671 37247
rect 19978 37244 19984 37256
rect 19659 37216 19984 37244
rect 19659 37213 19671 37216
rect 19613 37207 19671 37213
rect 12406 37148 14596 37176
rect 14 37068 20 37120
rect 72 37108 78 37120
rect 1489 37111 1547 37117
rect 1489 37108 1501 37111
rect 72 37080 1501 37108
rect 72 37068 78 37080
rect 1489 37077 1501 37080
rect 1535 37077 1547 37111
rect 1489 37071 1547 37077
rect 1946 37068 1952 37120
rect 2004 37108 2010 37120
rect 2225 37111 2283 37117
rect 2225 37108 2237 37111
rect 2004 37080 2237 37108
rect 2004 37068 2010 37080
rect 2225 37077 2237 37080
rect 2271 37077 2283 37111
rect 2225 37071 2283 37077
rect 5902 37068 5908 37120
rect 5960 37108 5966 37120
rect 6549 37111 6607 37117
rect 6549 37108 6561 37111
rect 5960 37080 6561 37108
rect 5960 37068 5966 37080
rect 6549 37077 6561 37080
rect 6595 37077 6607 37111
rect 8018 37108 8024 37120
rect 7979 37080 8024 37108
rect 6549 37071 6607 37077
rect 8018 37068 8024 37080
rect 8076 37068 8082 37120
rect 11514 37068 11520 37120
rect 11572 37108 11578 37120
rect 12406 37108 12434 37148
rect 11572 37080 12434 37108
rect 11572 37068 11578 37080
rect 16574 37068 16580 37120
rect 16632 37108 16638 37120
rect 16853 37111 16911 37117
rect 16853 37108 16865 37111
rect 16632 37080 16865 37108
rect 16632 37068 16638 37080
rect 16853 37077 16865 37080
rect 16899 37077 16911 37111
rect 16853 37071 16911 37077
rect 18046 37068 18052 37120
rect 18104 37108 18110 37120
rect 18233 37111 18291 37117
rect 18233 37108 18245 37111
rect 18104 37080 18245 37108
rect 18104 37068 18110 37080
rect 18233 37077 18245 37080
rect 18279 37077 18291 37111
rect 18432 37108 18460 37207
rect 19978 37204 19984 37216
rect 20036 37244 20042 37256
rect 20165 37247 20223 37253
rect 20165 37244 20177 37247
rect 20036 37216 20177 37244
rect 20036 37204 20042 37216
rect 20165 37213 20177 37216
rect 20211 37213 20223 37247
rect 23860 37244 23888 37340
rect 28721 37315 28779 37321
rect 28721 37281 28733 37315
rect 28767 37312 28779 37315
rect 28902 37312 28908 37324
rect 28767 37284 28908 37312
rect 28767 37281 28779 37284
rect 28721 37275 28779 37281
rect 28902 37272 28908 37284
rect 28960 37272 28966 37324
rect 29917 37315 29975 37321
rect 29917 37281 29929 37315
rect 29963 37312 29975 37315
rect 30282 37312 30288 37324
rect 29963 37284 30288 37312
rect 29963 37281 29975 37284
rect 29917 37275 29975 37281
rect 30282 37272 30288 37284
rect 30340 37312 30346 37324
rect 30653 37315 30711 37321
rect 30340 37284 30512 37312
rect 30340 37272 30346 37284
rect 24397 37247 24455 37253
rect 24397 37244 24409 37247
rect 20165 37207 20223 37213
rect 22066 37216 23796 37244
rect 23860 37216 24409 37244
rect 20254 37136 20260 37188
rect 20312 37176 20318 37188
rect 20533 37179 20591 37185
rect 20533 37176 20545 37179
rect 20312 37148 20545 37176
rect 20312 37136 20318 37148
rect 20533 37145 20545 37148
rect 20579 37145 20591 37179
rect 20533 37139 20591 37145
rect 22066 37108 22094 37216
rect 22186 37136 22192 37188
rect 22244 37176 22250 37188
rect 22373 37179 22431 37185
rect 22373 37176 22385 37179
rect 22244 37148 22385 37176
rect 22244 37136 22250 37148
rect 22373 37145 22385 37148
rect 22419 37176 22431 37179
rect 22925 37179 22983 37185
rect 22925 37176 22937 37179
rect 22419 37148 22937 37176
rect 22419 37145 22431 37148
rect 22373 37139 22431 37145
rect 22925 37145 22937 37148
rect 22971 37145 22983 37179
rect 23768 37176 23796 37216
rect 24397 37213 24409 37216
rect 24443 37213 24455 37247
rect 24397 37207 24455 37213
rect 25409 37247 25467 37253
rect 25409 37213 25421 37247
rect 25455 37244 25467 37247
rect 25774 37244 25780 37256
rect 25455 37216 25780 37244
rect 25455 37213 25467 37216
rect 25409 37207 25467 37213
rect 25774 37204 25780 37216
rect 25832 37244 25838 37256
rect 25869 37247 25927 37253
rect 25869 37244 25881 37247
rect 25832 37216 25881 37244
rect 25832 37204 25838 37216
rect 25869 37213 25881 37216
rect 25915 37213 25927 37247
rect 25869 37207 25927 37213
rect 27985 37247 28043 37253
rect 27985 37213 27997 37247
rect 28031 37244 28043 37247
rect 28350 37244 28356 37256
rect 28031 37216 28356 37244
rect 28031 37213 28043 37216
rect 27985 37207 28043 37213
rect 28350 37204 28356 37216
rect 28408 37244 28414 37256
rect 30484 37253 30512 37284
rect 30653 37281 30665 37315
rect 30699 37312 30711 37315
rect 37660 37312 37688 37352
rect 46750 37340 46756 37352
rect 46808 37340 46814 37392
rect 43257 37315 43315 37321
rect 43257 37312 43269 37315
rect 30699 37284 37688 37312
rect 41892 37284 43269 37312
rect 30699 37281 30711 37284
rect 30653 37275 30711 37281
rect 41892 37256 41920 37284
rect 43257 37281 43269 37284
rect 43303 37281 43315 37315
rect 43257 37275 43315 37281
rect 47026 37272 47032 37324
rect 47084 37312 47090 37324
rect 48041 37315 48099 37321
rect 48041 37312 48053 37315
rect 47084 37284 48053 37312
rect 47084 37272 47090 37284
rect 48041 37281 48053 37284
rect 48087 37281 48099 37315
rect 48041 37275 48099 37281
rect 52181 37315 52239 37321
rect 52181 37281 52193 37315
rect 52227 37312 52239 37315
rect 52227 37284 52592 37312
rect 52227 37281 52239 37284
rect 52181 37275 52239 37281
rect 52564 37256 52592 37284
rect 28537 37247 28595 37253
rect 28537 37244 28549 37247
rect 28408 37216 28549 37244
rect 28408 37204 28414 37216
rect 28537 37213 28549 37216
rect 28583 37213 28595 37247
rect 28537 37207 28595 37213
rect 30469 37247 30527 37253
rect 30469 37213 30481 37247
rect 30515 37213 30527 37247
rect 32582 37244 32588 37256
rect 32543 37216 32588 37244
rect 30469 37207 30527 37213
rect 32582 37204 32588 37216
rect 32640 37204 32646 37256
rect 33505 37247 33563 37253
rect 33505 37213 33517 37247
rect 33551 37244 33563 37247
rect 33965 37247 34023 37253
rect 33965 37244 33977 37247
rect 33551 37216 33977 37244
rect 33551 37213 33563 37216
rect 33505 37207 33563 37213
rect 33965 37213 33977 37216
rect 34011 37244 34023 37247
rect 34146 37244 34152 37256
rect 34011 37216 34152 37244
rect 34011 37213 34023 37216
rect 33965 37207 34023 37213
rect 34146 37204 34152 37216
rect 34204 37204 34210 37256
rect 35802 37204 35808 37256
rect 35860 37244 35866 37256
rect 35897 37247 35955 37253
rect 35897 37244 35909 37247
rect 35860 37216 35909 37244
rect 35860 37204 35866 37216
rect 35897 37213 35909 37216
rect 35943 37213 35955 37247
rect 35897 37207 35955 37213
rect 36170 37204 36176 37256
rect 36228 37244 36234 37256
rect 37182 37244 37188 37256
rect 36228 37216 37188 37244
rect 36228 37204 36234 37216
rect 37182 37204 37188 37216
rect 37240 37244 37246 37256
rect 37737 37247 37795 37253
rect 37737 37244 37749 37247
rect 37240 37216 37749 37244
rect 37240 37204 37246 37216
rect 37737 37213 37749 37216
rect 37783 37213 37795 37247
rect 39022 37244 39028 37256
rect 38983 37216 39028 37244
rect 37737 37207 37795 37213
rect 39022 37204 39028 37216
rect 39080 37204 39086 37256
rect 39114 37204 39120 37256
rect 39172 37244 39178 37256
rect 40126 37244 40132 37256
rect 39172 37216 39217 37244
rect 40087 37216 40132 37244
rect 39172 37204 39178 37216
rect 40126 37204 40132 37216
rect 40184 37204 40190 37256
rect 40865 37247 40923 37253
rect 40865 37213 40877 37247
rect 40911 37244 40923 37247
rect 41046 37244 41052 37256
rect 40911 37216 41052 37244
rect 40911 37213 40923 37216
rect 40865 37207 40923 37213
rect 41046 37204 41052 37216
rect 41104 37204 41110 37256
rect 41693 37247 41751 37253
rect 41693 37213 41705 37247
rect 41739 37244 41751 37247
rect 41874 37244 41880 37256
rect 41739 37216 41880 37244
rect 41739 37213 41751 37216
rect 41693 37207 41751 37213
rect 41874 37204 41880 37216
rect 41932 37204 41938 37256
rect 42518 37204 42524 37256
rect 42576 37244 42582 37256
rect 42613 37247 42671 37253
rect 42613 37244 42625 37247
rect 42576 37216 42625 37244
rect 42576 37204 42582 37216
rect 42613 37213 42625 37216
rect 42659 37213 42671 37247
rect 42613 37207 42671 37213
rect 42705 37247 42763 37253
rect 42705 37213 42717 37247
rect 42751 37213 42763 37247
rect 42705 37207 42763 37213
rect 46477 37247 46535 37253
rect 46477 37213 46489 37247
rect 46523 37244 46535 37247
rect 47578 37244 47584 37256
rect 46523 37216 47584 37244
rect 46523 37213 46535 37216
rect 46477 37207 46535 37213
rect 28626 37176 28632 37188
rect 23768 37148 28632 37176
rect 22925 37139 22983 37145
rect 28626 37136 28632 37148
rect 28684 37136 28690 37188
rect 34790 37176 34796 37188
rect 34751 37148 34796 37176
rect 34790 37136 34796 37148
rect 34848 37136 34854 37188
rect 34977 37179 35035 37185
rect 34977 37145 34989 37179
rect 35023 37145 35035 37179
rect 35618 37176 35624 37188
rect 35579 37148 35624 37176
rect 34977 37139 35035 37145
rect 22278 37108 22284 37120
rect 18432 37080 22094 37108
rect 22239 37080 22284 37108
rect 18233 37071 18291 37077
rect 22278 37068 22284 37080
rect 22336 37068 22342 37120
rect 24578 37108 24584 37120
rect 24539 37080 24584 37108
rect 24578 37068 24584 37080
rect 24636 37068 24642 37120
rect 26053 37111 26111 37117
rect 26053 37077 26065 37111
rect 26099 37108 26111 37111
rect 26142 37108 26148 37120
rect 26099 37080 26148 37108
rect 26099 37077 26111 37080
rect 26053 37071 26111 37077
rect 26142 37068 26148 37080
rect 26200 37068 26206 37120
rect 32214 37068 32220 37120
rect 32272 37108 32278 37120
rect 32401 37111 32459 37117
rect 32401 37108 32413 37111
rect 32272 37080 32413 37108
rect 32272 37068 32278 37080
rect 32401 37077 32413 37080
rect 32447 37077 32459 37111
rect 32401 37071 32459 37077
rect 34149 37111 34207 37117
rect 34149 37077 34161 37111
rect 34195 37108 34207 37111
rect 34698 37108 34704 37120
rect 34195 37080 34704 37108
rect 34195 37077 34207 37080
rect 34149 37071 34207 37077
rect 34698 37068 34704 37080
rect 34756 37108 34762 37120
rect 34992 37108 35020 37139
rect 35618 37136 35624 37148
rect 35676 37136 35682 37188
rect 36081 37179 36139 37185
rect 36081 37145 36093 37179
rect 36127 37145 36139 37179
rect 36081 37139 36139 37145
rect 34756 37080 35020 37108
rect 35161 37111 35219 37117
rect 34756 37068 34762 37080
rect 35161 37077 35173 37111
rect 35207 37108 35219 37111
rect 35526 37108 35532 37120
rect 35207 37080 35532 37108
rect 35207 37077 35219 37080
rect 35161 37071 35219 37077
rect 35526 37068 35532 37080
rect 35584 37108 35590 37120
rect 35713 37111 35771 37117
rect 35713 37108 35725 37111
rect 35584 37080 35725 37108
rect 35584 37068 35590 37080
rect 35713 37077 35725 37080
rect 35759 37077 35771 37111
rect 36096 37108 36124 37139
rect 38010 37136 38016 37188
rect 38068 37176 38074 37188
rect 42720 37176 42748 37207
rect 47578 37204 47584 37216
rect 47636 37204 47642 37256
rect 48406 37204 48412 37256
rect 48464 37244 48470 37256
rect 48958 37244 48964 37256
rect 48464 37216 48964 37244
rect 48464 37204 48470 37216
rect 48958 37204 48964 37216
rect 49016 37204 49022 37256
rect 50246 37204 50252 37256
rect 50304 37244 50310 37256
rect 50617 37247 50675 37253
rect 50617 37244 50629 37247
rect 50304 37216 50629 37244
rect 50304 37204 50310 37216
rect 50617 37213 50629 37216
rect 50663 37213 50675 37247
rect 50617 37207 50675 37213
rect 52546 37204 52552 37256
rect 52604 37244 52610 37256
rect 52733 37247 52791 37253
rect 52733 37244 52745 37247
rect 52604 37216 52745 37244
rect 52604 37204 52610 37216
rect 52733 37213 52745 37216
rect 52779 37213 52791 37247
rect 54202 37244 54208 37256
rect 54163 37216 54208 37244
rect 52733 37207 52791 37213
rect 54202 37204 54208 37216
rect 54260 37204 54266 37256
rect 55677 37247 55735 37253
rect 55677 37213 55689 37247
rect 55723 37244 55735 37247
rect 56042 37244 56048 37256
rect 55723 37216 56048 37244
rect 55723 37213 55735 37216
rect 55677 37207 55735 37213
rect 56042 37204 56048 37216
rect 56100 37244 56106 37256
rect 56229 37247 56287 37253
rect 56229 37244 56241 37247
rect 56100 37216 56241 37244
rect 56100 37204 56106 37216
rect 56229 37213 56241 37216
rect 56275 37213 56287 37247
rect 56229 37207 56287 37213
rect 57885 37247 57943 37253
rect 57885 37213 57897 37247
rect 57931 37244 57943 37247
rect 57974 37244 57980 37256
rect 57931 37216 57980 37244
rect 57931 37213 57943 37216
rect 57885 37207 57943 37213
rect 57974 37204 57980 37216
rect 58032 37204 58038 37256
rect 43714 37176 43720 37188
rect 38068 37148 39988 37176
rect 38068 37136 38074 37148
rect 38286 37108 38292 37120
rect 36096 37080 38292 37108
rect 35713 37071 35771 37077
rect 38286 37068 38292 37080
rect 38344 37068 38350 37120
rect 38841 37111 38899 37117
rect 38841 37077 38853 37111
rect 38887 37108 38899 37111
rect 39206 37108 39212 37120
rect 38887 37080 39212 37108
rect 38887 37077 38899 37080
rect 38841 37071 38899 37077
rect 39206 37068 39212 37080
rect 39264 37068 39270 37120
rect 39960 37117 39988 37148
rect 41892 37148 43720 37176
rect 39945 37111 40003 37117
rect 39945 37077 39957 37111
rect 39991 37077 40003 37111
rect 39945 37071 40003 37077
rect 40034 37068 40040 37120
rect 40092 37108 40098 37120
rect 41892 37117 41920 37148
rect 43714 37136 43720 37148
rect 43772 37136 43778 37188
rect 46106 37136 46112 37188
rect 46164 37176 46170 37188
rect 46201 37179 46259 37185
rect 46201 37176 46213 37179
rect 46164 37148 46213 37176
rect 46164 37136 46170 37148
rect 46201 37145 46213 37148
rect 46247 37145 46259 37179
rect 46201 37139 46259 37145
rect 46661 37179 46719 37185
rect 46661 37145 46673 37179
rect 46707 37145 46719 37179
rect 46661 37139 46719 37145
rect 40681 37111 40739 37117
rect 40681 37108 40693 37111
rect 40092 37080 40693 37108
rect 40092 37068 40098 37080
rect 40681 37077 40693 37080
rect 40727 37077 40739 37111
rect 40681 37071 40739 37077
rect 41877 37111 41935 37117
rect 41877 37077 41889 37111
rect 41923 37077 41935 37111
rect 41877 37071 41935 37077
rect 42429 37111 42487 37117
rect 42429 37077 42441 37111
rect 42475 37108 42487 37111
rect 42610 37108 42616 37120
rect 42475 37080 42616 37108
rect 42475 37077 42487 37080
rect 42429 37071 42487 37077
rect 42610 37068 42616 37080
rect 42668 37068 42674 37120
rect 46293 37111 46351 37117
rect 46293 37077 46305 37111
rect 46339 37108 46351 37111
rect 46566 37108 46572 37120
rect 46339 37080 46572 37108
rect 46339 37077 46351 37080
rect 46293 37071 46351 37077
rect 46566 37068 46572 37080
rect 46624 37068 46630 37120
rect 46676 37108 46704 37139
rect 46934 37136 46940 37188
rect 46992 37176 46998 37188
rect 48222 37176 48228 37188
rect 46992 37148 48228 37176
rect 46992 37136 46998 37148
rect 48222 37136 48228 37148
rect 48280 37176 48286 37188
rect 48317 37179 48375 37185
rect 48317 37176 48329 37179
rect 48280 37148 48329 37176
rect 48280 37136 48286 37148
rect 48317 37145 48329 37148
rect 48363 37145 48375 37179
rect 56686 37176 56692 37188
rect 56647 37148 56692 37176
rect 48317 37139 48375 37145
rect 56686 37136 56692 37148
rect 56744 37136 56750 37188
rect 50062 37108 50068 37120
rect 46676 37080 50068 37108
rect 50062 37068 50068 37080
rect 50120 37068 50126 37120
rect 50706 37108 50712 37120
rect 50667 37080 50712 37108
rect 50706 37068 50712 37080
rect 50764 37068 50770 37120
rect 52178 37068 52184 37120
rect 52236 37108 52242 37120
rect 52917 37111 52975 37117
rect 52917 37108 52929 37111
rect 52236 37080 52929 37108
rect 52236 37068 52242 37080
rect 52917 37077 52929 37080
rect 52963 37077 52975 37111
rect 52917 37071 52975 37077
rect 54110 37068 54116 37120
rect 54168 37108 54174 37120
rect 54389 37111 54447 37117
rect 54389 37108 54401 37111
rect 54168 37080 54401 37108
rect 54168 37068 54174 37080
rect 54389 37077 54401 37080
rect 54435 37077 54447 37111
rect 54389 37071 54447 37077
rect 56594 37068 56600 37120
rect 56652 37108 56658 37120
rect 58069 37111 58127 37117
rect 58069 37108 58081 37111
rect 56652 37080 58081 37108
rect 56652 37068 56658 37080
rect 58069 37077 58081 37080
rect 58115 37077 58127 37111
rect 58069 37071 58127 37077
rect 58158 37068 58164 37120
rect 58216 37108 58222 37120
rect 59906 37108 59912 37120
rect 58216 37080 59912 37108
rect 58216 37068 58222 37080
rect 59906 37068 59912 37080
rect 59964 37068 59970 37120
rect 1104 37018 58880 37040
rect 1104 36966 19574 37018
rect 19626 36966 19638 37018
rect 19690 36966 19702 37018
rect 19754 36966 19766 37018
rect 19818 36966 19830 37018
rect 19882 36966 50294 37018
rect 50346 36966 50358 37018
rect 50410 36966 50422 37018
rect 50474 36966 50486 37018
rect 50538 36966 50550 37018
rect 50602 36966 58880 37018
rect 1104 36944 58880 36966
rect 1486 36904 1492 36916
rect 1447 36876 1492 36904
rect 1486 36864 1492 36876
rect 1544 36864 1550 36916
rect 3878 36864 3884 36916
rect 3936 36904 3942 36916
rect 3973 36907 4031 36913
rect 3973 36904 3985 36907
rect 3936 36876 3985 36904
rect 3936 36864 3942 36876
rect 3973 36873 3985 36876
rect 4019 36873 4031 36907
rect 3973 36867 4031 36873
rect 4062 36864 4068 36916
rect 4120 36904 4126 36916
rect 24578 36904 24584 36916
rect 4120 36876 24584 36904
rect 4120 36864 4126 36876
rect 24578 36864 24584 36876
rect 24636 36864 24642 36916
rect 26329 36907 26387 36913
rect 26329 36873 26341 36907
rect 26375 36904 26387 36907
rect 32398 36904 32404 36916
rect 26375 36876 32404 36904
rect 26375 36873 26387 36876
rect 26329 36867 26387 36873
rect 32398 36864 32404 36876
rect 32456 36864 32462 36916
rect 37182 36864 37188 36916
rect 37240 36904 37246 36916
rect 37461 36907 37519 36913
rect 37461 36904 37473 36907
rect 37240 36876 37473 36904
rect 37240 36864 37246 36876
rect 37461 36873 37473 36876
rect 37507 36873 37519 36907
rect 37461 36867 37519 36873
rect 39022 36864 39028 36916
rect 39080 36904 39086 36916
rect 39080 36876 39528 36904
rect 39080 36864 39086 36876
rect 8481 36839 8539 36845
rect 8481 36836 8493 36839
rect 6748 36808 8493 36836
rect 6748 36780 6776 36808
rect 8481 36805 8493 36808
rect 8527 36805 8539 36839
rect 14182 36836 14188 36848
rect 14143 36808 14188 36836
rect 8481 36799 8539 36805
rect 14182 36796 14188 36808
rect 14240 36796 14246 36848
rect 20809 36839 20867 36845
rect 20809 36805 20821 36839
rect 20855 36836 20867 36839
rect 26510 36836 26516 36848
rect 20855 36808 26516 36836
rect 20855 36805 20867 36808
rect 20809 36799 20867 36805
rect 26510 36796 26516 36808
rect 26568 36836 26574 36848
rect 28074 36836 28080 36848
rect 26568 36808 27844 36836
rect 28035 36808 28080 36836
rect 26568 36796 26574 36808
rect 1673 36771 1731 36777
rect 1673 36737 1685 36771
rect 1719 36768 1731 36771
rect 2038 36768 2044 36780
rect 1719 36740 2044 36768
rect 1719 36737 1731 36740
rect 1673 36731 1731 36737
rect 2038 36728 2044 36740
rect 2096 36728 2102 36780
rect 5445 36771 5503 36777
rect 5445 36737 5457 36771
rect 5491 36768 5503 36771
rect 6730 36768 6736 36780
rect 5491 36740 6736 36768
rect 5491 36737 5503 36740
rect 5445 36731 5503 36737
rect 6730 36728 6736 36740
rect 6788 36728 6794 36780
rect 7466 36768 7472 36780
rect 7427 36740 7472 36768
rect 7466 36728 7472 36740
rect 7524 36728 7530 36780
rect 8294 36768 8300 36780
rect 8255 36740 8300 36768
rect 8294 36728 8300 36740
rect 8352 36728 8358 36780
rect 8570 36768 8576 36780
rect 8531 36740 8576 36768
rect 8570 36728 8576 36740
rect 8628 36768 8634 36780
rect 9033 36771 9091 36777
rect 9033 36768 9045 36771
rect 8628 36740 9045 36768
rect 8628 36728 8634 36740
rect 9033 36737 9045 36740
rect 9079 36737 9091 36771
rect 9033 36731 9091 36737
rect 20165 36771 20223 36777
rect 20165 36737 20177 36771
rect 20211 36768 20223 36771
rect 21266 36768 21272 36780
rect 20211 36740 21272 36768
rect 20211 36737 20223 36740
rect 20165 36731 20223 36737
rect 21266 36728 21272 36740
rect 21324 36728 21330 36780
rect 22465 36771 22523 36777
rect 22465 36737 22477 36771
rect 22511 36768 22523 36771
rect 23474 36768 23480 36780
rect 22511 36740 23480 36768
rect 22511 36737 22523 36740
rect 22465 36731 22523 36737
rect 23474 36728 23480 36740
rect 23532 36728 23538 36780
rect 23842 36728 23848 36780
rect 23900 36768 23906 36780
rect 24121 36771 24179 36777
rect 24121 36768 24133 36771
rect 23900 36740 24133 36768
rect 23900 36728 23906 36740
rect 24121 36737 24133 36740
rect 24167 36737 24179 36771
rect 24121 36731 24179 36737
rect 24949 36771 25007 36777
rect 24949 36737 24961 36771
rect 24995 36768 25007 36771
rect 26145 36771 26203 36777
rect 26145 36768 26157 36771
rect 24995 36740 26157 36768
rect 24995 36737 25007 36740
rect 24949 36731 25007 36737
rect 26145 36737 26157 36740
rect 26191 36768 26203 36771
rect 26191 36740 27186 36768
rect 26191 36737 26203 36740
rect 26145 36731 26203 36737
rect 5537 36703 5595 36709
rect 5537 36669 5549 36703
rect 5583 36669 5595 36703
rect 5810 36700 5816 36712
rect 5771 36672 5816 36700
rect 5537 36663 5595 36669
rect 5552 36632 5580 36663
rect 5810 36660 5816 36672
rect 5868 36660 5874 36712
rect 7098 36700 7104 36712
rect 7059 36672 7104 36700
rect 7098 36660 7104 36672
rect 7156 36660 7162 36712
rect 7561 36703 7619 36709
rect 7561 36669 7573 36703
rect 7607 36700 7619 36703
rect 8113 36703 8171 36709
rect 8113 36700 8125 36703
rect 7607 36672 8125 36700
rect 7607 36669 7619 36672
rect 7561 36663 7619 36669
rect 8113 36669 8125 36672
rect 8159 36669 8171 36703
rect 8113 36663 8171 36669
rect 19426 36660 19432 36712
rect 19484 36700 19490 36712
rect 19889 36703 19947 36709
rect 19889 36700 19901 36703
rect 19484 36672 19901 36700
rect 19484 36660 19490 36672
rect 19889 36669 19901 36672
rect 19935 36669 19947 36703
rect 19889 36663 19947 36669
rect 21726 36660 21732 36712
rect 21784 36700 21790 36712
rect 22373 36703 22431 36709
rect 22373 36700 22385 36703
rect 21784 36672 22385 36700
rect 21784 36660 21790 36672
rect 22373 36669 22385 36672
rect 22419 36669 22431 36703
rect 24029 36703 24087 36709
rect 24029 36700 24041 36703
rect 22373 36663 22431 36669
rect 22848 36672 24041 36700
rect 22848 36641 22876 36672
rect 24029 36669 24041 36672
rect 24075 36700 24087 36703
rect 24394 36700 24400 36712
rect 24075 36672 24400 36700
rect 24075 36669 24087 36672
rect 24029 36663 24087 36669
rect 24394 36660 24400 36672
rect 24452 36660 24458 36712
rect 25682 36700 25688 36712
rect 25643 36672 25688 36700
rect 25682 36660 25688 36672
rect 25740 36660 25746 36712
rect 26053 36703 26111 36709
rect 26053 36669 26065 36703
rect 26099 36700 26111 36703
rect 26418 36700 26424 36712
rect 26099 36672 26424 36700
rect 26099 36669 26111 36672
rect 26053 36663 26111 36669
rect 26418 36660 26424 36672
rect 26476 36700 26482 36712
rect 27249 36703 27307 36709
rect 27249 36700 27261 36703
rect 26476 36672 27261 36700
rect 26476 36660 26482 36672
rect 27249 36669 27261 36672
rect 27295 36669 27307 36703
rect 27816 36700 27844 36808
rect 28074 36796 28080 36808
rect 28132 36796 28138 36848
rect 38381 36839 38439 36845
rect 38381 36805 38393 36839
rect 38427 36836 38439 36839
rect 38427 36808 38516 36836
rect 38427 36805 38439 36808
rect 38381 36799 38439 36805
rect 27890 36728 27896 36780
rect 27948 36768 27954 36780
rect 28721 36771 28779 36777
rect 28721 36768 28733 36771
rect 27948 36740 28733 36768
rect 27948 36728 27954 36740
rect 28721 36737 28733 36740
rect 28767 36737 28779 36771
rect 28721 36731 28779 36737
rect 31294 36728 31300 36780
rect 31352 36768 31358 36780
rect 32309 36771 32367 36777
rect 32309 36768 32321 36771
rect 31352 36740 32321 36768
rect 31352 36728 31358 36740
rect 32309 36737 32321 36740
rect 32355 36737 32367 36771
rect 34698 36768 34704 36780
rect 34659 36740 34704 36768
rect 32309 36731 32367 36737
rect 34698 36728 34704 36740
rect 34756 36728 34762 36780
rect 34790 36728 34796 36780
rect 34848 36768 34854 36780
rect 34885 36771 34943 36777
rect 34885 36768 34897 36771
rect 34848 36740 34897 36768
rect 34848 36728 34854 36740
rect 34885 36737 34897 36740
rect 34931 36737 34943 36771
rect 35526 36768 35532 36780
rect 35487 36740 35532 36768
rect 34885 36731 34943 36737
rect 35526 36728 35532 36740
rect 35584 36728 35590 36780
rect 38286 36768 38292 36780
rect 38247 36740 38292 36768
rect 38286 36728 38292 36740
rect 38344 36728 38350 36780
rect 28629 36703 28687 36709
rect 28629 36700 28641 36703
rect 27816 36672 28641 36700
rect 27249 36663 27307 36669
rect 28629 36669 28641 36672
rect 28675 36669 28687 36703
rect 28629 36663 28687 36669
rect 31570 36660 31576 36712
rect 31628 36700 31634 36712
rect 32401 36703 32459 36709
rect 32401 36700 32413 36703
rect 31628 36672 32413 36700
rect 31628 36660 31634 36672
rect 32401 36669 32413 36672
rect 32447 36700 32459 36703
rect 33410 36700 33416 36712
rect 32447 36672 33416 36700
rect 32447 36669 32459 36672
rect 32401 36663 32459 36669
rect 33410 36660 33416 36672
rect 33468 36660 33474 36712
rect 22833 36635 22891 36641
rect 5552 36604 6500 36632
rect 6472 36573 6500 36604
rect 22833 36601 22845 36635
rect 22879 36601 22891 36635
rect 22833 36595 22891 36601
rect 23474 36592 23480 36644
rect 23532 36632 23538 36644
rect 30834 36632 30840 36644
rect 23532 36604 30840 36632
rect 23532 36592 23538 36604
rect 30834 36592 30840 36604
rect 30892 36632 30898 36644
rect 33594 36632 33600 36644
rect 30892 36604 33600 36632
rect 30892 36592 30898 36604
rect 33594 36592 33600 36604
rect 33652 36592 33658 36644
rect 38488 36632 38516 36808
rect 38565 36771 38623 36777
rect 38565 36737 38577 36771
rect 38611 36737 38623 36771
rect 38565 36731 38623 36737
rect 39301 36771 39359 36777
rect 39301 36737 39313 36771
rect 39347 36737 39359 36771
rect 39500 36768 39528 36876
rect 40126 36864 40132 36916
rect 40184 36904 40190 36916
rect 47394 36904 47400 36916
rect 40184 36876 47400 36904
rect 40184 36864 40190 36876
rect 47394 36864 47400 36876
rect 47452 36864 47458 36916
rect 47578 36904 47584 36916
rect 47539 36876 47584 36904
rect 47578 36864 47584 36876
rect 47636 36864 47642 36916
rect 48222 36864 48228 36916
rect 48280 36904 48286 36916
rect 48409 36907 48467 36913
rect 48409 36904 48421 36907
rect 48280 36876 48421 36904
rect 48280 36864 48286 36876
rect 48409 36873 48421 36876
rect 48455 36873 48467 36907
rect 48958 36904 48964 36916
rect 48919 36876 48964 36904
rect 48409 36867 48467 36873
rect 48958 36864 48964 36876
rect 49016 36864 49022 36916
rect 50154 36864 50160 36916
rect 50212 36904 50218 36916
rect 50341 36907 50399 36913
rect 50341 36904 50353 36907
rect 50212 36876 50353 36904
rect 50212 36864 50218 36876
rect 50341 36873 50353 36876
rect 50387 36873 50399 36907
rect 50341 36867 50399 36873
rect 57333 36907 57391 36913
rect 57333 36873 57345 36907
rect 57379 36904 57391 36907
rect 57974 36904 57980 36916
rect 57379 36876 57980 36904
rect 57379 36873 57391 36876
rect 57333 36867 57391 36873
rect 57974 36864 57980 36876
rect 58032 36864 58038 36916
rect 41785 36839 41843 36845
rect 41785 36805 41797 36839
rect 41831 36836 41843 36839
rect 43901 36839 43959 36845
rect 43901 36836 43913 36839
rect 41831 36808 43913 36836
rect 41831 36805 41843 36808
rect 41785 36799 41843 36805
rect 40313 36771 40371 36777
rect 40313 36768 40325 36771
rect 39500 36740 40325 36768
rect 39301 36731 39359 36737
rect 40313 36737 40325 36740
rect 40359 36737 40371 36771
rect 40313 36731 40371 36737
rect 40497 36771 40555 36777
rect 40497 36737 40509 36771
rect 40543 36737 40555 36771
rect 40497 36731 40555 36737
rect 41601 36771 41659 36777
rect 41601 36737 41613 36771
rect 41647 36737 41659 36771
rect 41874 36768 41880 36780
rect 41835 36740 41880 36768
rect 41601 36731 41659 36737
rect 38580 36700 38608 36731
rect 39206 36700 39212 36712
rect 38580 36672 39212 36700
rect 39206 36660 39212 36672
rect 39264 36660 39270 36712
rect 39316 36632 39344 36731
rect 40126 36660 40132 36712
rect 40184 36700 40190 36712
rect 40512 36700 40540 36731
rect 40184 36672 40540 36700
rect 41616 36700 41644 36731
rect 41874 36728 41880 36740
rect 41932 36728 41938 36780
rect 42536 36777 42564 36808
rect 43901 36805 43913 36808
rect 43947 36805 43959 36839
rect 46382 36836 46388 36848
rect 46046 36808 46388 36836
rect 43901 36799 43959 36805
rect 46382 36796 46388 36808
rect 46440 36796 46446 36848
rect 56781 36839 56839 36845
rect 56781 36805 56793 36839
rect 56827 36836 56839 36839
rect 57882 36836 57888 36848
rect 56827 36808 57888 36836
rect 56827 36805 56839 36808
rect 56781 36799 56839 36805
rect 57882 36796 57888 36808
rect 57940 36836 57946 36848
rect 58069 36839 58127 36845
rect 58069 36836 58081 36839
rect 57940 36808 58081 36836
rect 57940 36796 57946 36808
rect 58069 36805 58081 36808
rect 58115 36805 58127 36839
rect 58069 36799 58127 36805
rect 42521 36771 42579 36777
rect 42521 36737 42533 36771
rect 42567 36737 42579 36771
rect 42521 36731 42579 36737
rect 42702 36728 42708 36780
rect 42760 36768 42766 36780
rect 43533 36771 43591 36777
rect 43533 36768 43545 36771
rect 42760 36740 43545 36768
rect 42760 36728 42766 36740
rect 43533 36737 43545 36740
rect 43579 36737 43591 36771
rect 43714 36768 43720 36780
rect 43675 36740 43720 36768
rect 43533 36731 43591 36737
rect 43714 36728 43720 36740
rect 43772 36728 43778 36780
rect 46106 36768 46112 36780
rect 46067 36740 46112 36768
rect 46106 36728 46112 36740
rect 46164 36728 46170 36780
rect 46566 36768 46572 36780
rect 46527 36740 46572 36768
rect 46566 36728 46572 36740
rect 46624 36728 46630 36780
rect 47118 36728 47124 36780
rect 47176 36768 47182 36780
rect 47765 36771 47823 36777
rect 47765 36768 47777 36771
rect 47176 36740 47777 36768
rect 47176 36728 47182 36740
rect 47765 36737 47777 36740
rect 47811 36737 47823 36771
rect 47765 36731 47823 36737
rect 42610 36700 42616 36712
rect 41616 36672 42616 36700
rect 40184 36660 40190 36672
rect 42610 36660 42616 36672
rect 42668 36660 42674 36712
rect 47670 36660 47676 36712
rect 47728 36700 47734 36712
rect 47949 36703 48007 36709
rect 47949 36700 47961 36703
rect 47728 36672 47961 36700
rect 47728 36660 47734 36672
rect 47949 36669 47961 36672
rect 47995 36700 48007 36703
rect 56594 36700 56600 36712
rect 47995 36672 56600 36700
rect 47995 36669 48007 36672
rect 47949 36663 48007 36669
rect 56594 36660 56600 36672
rect 56652 36660 56658 36712
rect 40681 36635 40739 36641
rect 40681 36632 40693 36635
rect 38488 36604 40693 36632
rect 40681 36601 40693 36604
rect 40727 36601 40739 36635
rect 57885 36635 57943 36641
rect 57885 36632 57897 36635
rect 40681 36595 40739 36601
rect 56612 36604 57897 36632
rect 56612 36576 56640 36604
rect 57885 36601 57897 36604
rect 57931 36601 57943 36635
rect 57885 36595 57943 36601
rect 6457 36567 6515 36573
rect 6457 36533 6469 36567
rect 6503 36564 6515 36567
rect 6638 36564 6644 36576
rect 6503 36536 6644 36564
rect 6503 36533 6515 36536
rect 6457 36527 6515 36533
rect 6638 36524 6644 36536
rect 6696 36524 6702 36576
rect 29086 36564 29092 36576
rect 29047 36536 29092 36564
rect 29086 36524 29092 36536
rect 29144 36524 29150 36576
rect 30190 36564 30196 36576
rect 30151 36536 30196 36564
rect 30190 36524 30196 36536
rect 30248 36524 30254 36576
rect 32490 36524 32496 36576
rect 32548 36564 32554 36576
rect 32677 36567 32735 36573
rect 32677 36564 32689 36567
rect 32548 36536 32689 36564
rect 32548 36524 32554 36536
rect 32677 36533 32689 36536
rect 32723 36533 32735 36567
rect 32677 36527 32735 36533
rect 35069 36567 35127 36573
rect 35069 36533 35081 36567
rect 35115 36564 35127 36567
rect 35802 36564 35808 36576
rect 35115 36536 35808 36564
rect 35115 36533 35127 36536
rect 35069 36527 35127 36533
rect 35802 36524 35808 36536
rect 35860 36524 35866 36576
rect 35989 36567 36047 36573
rect 35989 36533 36001 36567
rect 36035 36564 36047 36567
rect 36446 36564 36452 36576
rect 36035 36536 36452 36564
rect 36035 36533 36047 36536
rect 35989 36527 36047 36533
rect 36446 36524 36452 36536
rect 36504 36524 36510 36576
rect 38749 36567 38807 36573
rect 38749 36533 38761 36567
rect 38795 36564 38807 36567
rect 39298 36564 39304 36576
rect 38795 36536 39304 36564
rect 38795 36533 38807 36536
rect 38749 36527 38807 36533
rect 39298 36524 39304 36536
rect 39356 36524 39362 36576
rect 39390 36524 39396 36576
rect 39448 36564 39454 36576
rect 39761 36567 39819 36573
rect 39448 36536 39493 36564
rect 39448 36524 39454 36536
rect 39761 36533 39773 36567
rect 39807 36564 39819 36567
rect 40310 36564 40316 36576
rect 39807 36536 40316 36564
rect 39807 36533 39819 36536
rect 39761 36527 39819 36533
rect 40310 36524 40316 36536
rect 40368 36524 40374 36576
rect 41414 36564 41420 36576
rect 41375 36536 41420 36564
rect 41414 36524 41420 36536
rect 41472 36524 41478 36576
rect 42610 36564 42616 36576
rect 42571 36536 42616 36564
rect 42610 36524 42616 36536
rect 42668 36524 42674 36576
rect 42978 36564 42984 36576
rect 42939 36536 42984 36564
rect 42978 36524 42984 36536
rect 43036 36524 43042 36576
rect 56594 36524 56600 36576
rect 56652 36524 56658 36576
rect 1104 36474 58880 36496
rect 1104 36422 4214 36474
rect 4266 36422 4278 36474
rect 4330 36422 4342 36474
rect 4394 36422 4406 36474
rect 4458 36422 4470 36474
rect 4522 36422 34934 36474
rect 34986 36422 34998 36474
rect 35050 36422 35062 36474
rect 35114 36422 35126 36474
rect 35178 36422 35190 36474
rect 35242 36422 58880 36474
rect 1104 36400 58880 36422
rect 8294 36320 8300 36372
rect 8352 36360 8358 36372
rect 8938 36360 8944 36372
rect 8352 36332 8944 36360
rect 8352 36320 8358 36332
rect 8938 36320 8944 36332
rect 8996 36320 9002 36372
rect 19426 36360 19432 36372
rect 19387 36332 19432 36360
rect 19426 36320 19432 36332
rect 19484 36320 19490 36372
rect 21726 36360 21732 36372
rect 21687 36332 21732 36360
rect 21726 36320 21732 36332
rect 21784 36320 21790 36372
rect 23842 36360 23848 36372
rect 23803 36332 23848 36360
rect 23842 36320 23848 36332
rect 23900 36320 23906 36372
rect 24397 36363 24455 36369
rect 24397 36329 24409 36363
rect 24443 36329 24455 36363
rect 24397 36323 24455 36329
rect 24765 36363 24823 36369
rect 24765 36329 24777 36363
rect 24811 36360 24823 36363
rect 25682 36360 25688 36372
rect 24811 36332 25688 36360
rect 24811 36329 24823 36332
rect 24765 36323 24823 36329
rect 6638 36252 6644 36304
rect 6696 36292 6702 36304
rect 7101 36295 7159 36301
rect 7101 36292 7113 36295
rect 6696 36264 7113 36292
rect 6696 36252 6702 36264
rect 7101 36261 7113 36264
rect 7147 36292 7159 36295
rect 8570 36292 8576 36304
rect 7147 36264 8576 36292
rect 7147 36261 7159 36264
rect 7101 36255 7159 36261
rect 8570 36252 8576 36264
rect 8628 36252 8634 36304
rect 21266 36252 21272 36304
rect 21324 36292 21330 36304
rect 21324 36264 22416 36292
rect 21324 36252 21330 36264
rect 9309 36227 9367 36233
rect 9309 36224 9321 36227
rect 8220 36196 9321 36224
rect 1670 36156 1676 36168
rect 1631 36128 1676 36156
rect 1670 36116 1676 36128
rect 1728 36116 1734 36168
rect 8018 36116 8024 36168
rect 8076 36156 8082 36168
rect 8220 36165 8248 36196
rect 9309 36193 9321 36196
rect 9355 36193 9367 36227
rect 9309 36187 9367 36193
rect 19705 36227 19763 36233
rect 19705 36193 19717 36227
rect 19751 36224 19763 36227
rect 20070 36224 20076 36236
rect 19751 36196 20076 36224
rect 19751 36193 19763 36196
rect 19705 36187 19763 36193
rect 20070 36184 20076 36196
rect 20128 36224 20134 36236
rect 22189 36227 22247 36233
rect 22189 36224 22201 36227
rect 20128 36196 22201 36224
rect 20128 36184 20134 36196
rect 8205 36159 8263 36165
rect 8205 36156 8217 36159
rect 8076 36128 8217 36156
rect 8076 36116 8082 36128
rect 8205 36125 8217 36128
rect 8251 36125 8263 36159
rect 8205 36119 8263 36125
rect 8389 36159 8447 36165
rect 8389 36125 8401 36159
rect 8435 36156 8447 36159
rect 8846 36156 8852 36168
rect 8435 36128 8852 36156
rect 8435 36125 8447 36128
rect 8389 36119 8447 36125
rect 7745 36091 7803 36097
rect 7745 36057 7757 36091
rect 7791 36088 7803 36091
rect 8404 36088 8432 36119
rect 8846 36116 8852 36128
rect 8904 36156 8910 36168
rect 9125 36159 9183 36165
rect 9125 36156 9137 36159
rect 8904 36128 9137 36156
rect 8904 36116 8910 36128
rect 9125 36125 9137 36128
rect 9171 36156 9183 36159
rect 9769 36159 9827 36165
rect 9769 36156 9781 36159
rect 9171 36128 9781 36156
rect 9171 36125 9183 36128
rect 9125 36119 9183 36125
rect 9769 36125 9781 36128
rect 9815 36125 9827 36159
rect 19242 36156 19248 36168
rect 19203 36128 19248 36156
rect 9769 36119 9827 36125
rect 19242 36116 19248 36128
rect 19300 36116 19306 36168
rect 19334 36116 19340 36168
rect 19392 36156 19398 36168
rect 19429 36159 19487 36165
rect 19429 36156 19441 36159
rect 19392 36128 19441 36156
rect 19392 36116 19398 36128
rect 19429 36125 19441 36128
rect 19475 36125 19487 36159
rect 21266 36156 21272 36168
rect 21227 36128 21272 36156
rect 19429 36119 19487 36125
rect 21266 36116 21272 36128
rect 21324 36116 21330 36168
rect 21376 36165 21404 36196
rect 22189 36193 22201 36196
rect 22235 36193 22247 36227
rect 22189 36187 22247 36193
rect 21361 36159 21419 36165
rect 21361 36125 21373 36159
rect 21407 36125 21419 36159
rect 21361 36119 21419 36125
rect 21545 36159 21603 36165
rect 21545 36125 21557 36159
rect 21591 36156 21603 36159
rect 22094 36156 22100 36168
rect 21591 36128 22100 36156
rect 21591 36125 21603 36128
rect 21545 36119 21603 36125
rect 22094 36116 22100 36128
rect 22152 36116 22158 36168
rect 22388 36165 22416 36264
rect 24412 36224 24440 36323
rect 25682 36320 25688 36332
rect 25740 36320 25746 36372
rect 26418 36360 26424 36372
rect 26379 36332 26424 36360
rect 26418 36320 26424 36332
rect 26476 36320 26482 36372
rect 28626 36360 28632 36372
rect 28587 36332 28632 36360
rect 28626 36320 28632 36332
rect 28684 36320 28690 36372
rect 31570 36360 31576 36372
rect 31531 36332 31576 36360
rect 31570 36320 31576 36332
rect 31628 36320 31634 36372
rect 33413 36363 33471 36369
rect 33413 36360 33425 36363
rect 31726 36332 33425 36360
rect 27890 36292 27896 36304
rect 23860 36196 24440 36224
rect 26344 36264 27896 36292
rect 23860 36168 23888 36196
rect 22373 36159 22431 36165
rect 22373 36125 22385 36159
rect 22419 36125 22431 36159
rect 23658 36156 23664 36168
rect 23619 36128 23664 36156
rect 22373 36119 22431 36125
rect 23658 36116 23664 36128
rect 23716 36116 23722 36168
rect 23842 36116 23848 36168
rect 23900 36156 23906 36168
rect 24394 36156 24400 36168
rect 23900 36128 23993 36156
rect 24355 36128 24400 36156
rect 23900 36116 23906 36128
rect 24394 36116 24400 36128
rect 24452 36116 24458 36168
rect 24486 36116 24492 36168
rect 24544 36156 24550 36168
rect 26237 36159 26295 36165
rect 24544 36128 24589 36156
rect 24544 36116 24550 36128
rect 26237 36125 26249 36159
rect 26283 36156 26295 36159
rect 26344 36156 26372 36264
rect 27890 36252 27896 36264
rect 27948 36252 27954 36304
rect 31726 36292 31754 36332
rect 33413 36329 33425 36332
rect 33459 36329 33471 36363
rect 33413 36323 33471 36329
rect 38473 36363 38531 36369
rect 38473 36329 38485 36363
rect 38519 36360 38531 36363
rect 39022 36360 39028 36372
rect 38519 36332 39028 36360
rect 38519 36329 38531 36332
rect 38473 36323 38531 36329
rect 39022 36320 39028 36332
rect 39080 36320 39086 36372
rect 41414 36360 41420 36372
rect 39132 36332 41420 36360
rect 30668 36264 31754 36292
rect 32769 36295 32827 36301
rect 30668 36224 30696 36264
rect 32769 36261 32781 36295
rect 32815 36292 32827 36295
rect 34790 36292 34796 36304
rect 32815 36264 34796 36292
rect 32815 36261 32827 36264
rect 32769 36255 32827 36261
rect 34790 36252 34796 36264
rect 34848 36252 34854 36304
rect 35618 36252 35624 36304
rect 35676 36292 35682 36304
rect 35676 36264 38240 36292
rect 35676 36252 35682 36264
rect 28276 36196 30696 36224
rect 26283 36128 26372 36156
rect 26421 36159 26479 36165
rect 26283 36125 26295 36128
rect 26237 36119 26295 36125
rect 26421 36125 26433 36159
rect 26467 36150 26479 36159
rect 26510 36150 26516 36168
rect 26467 36125 26516 36150
rect 26421 36122 26516 36125
rect 26421 36119 26479 36122
rect 26510 36116 26516 36122
rect 26568 36116 26574 36168
rect 7791 36060 8432 36088
rect 22557 36091 22615 36097
rect 7791 36057 7803 36060
rect 7745 36051 7803 36057
rect 22557 36057 22569 36091
rect 22603 36088 22615 36091
rect 28276 36088 28304 36196
rect 28442 36156 28448 36168
rect 28403 36128 28448 36156
rect 28442 36116 28448 36128
rect 28500 36116 28506 36168
rect 28626 36156 28632 36168
rect 28587 36128 28632 36156
rect 28626 36116 28632 36128
rect 28684 36116 28690 36168
rect 29086 36116 29092 36168
rect 29144 36156 29150 36168
rect 30668 36165 30696 36196
rect 30745 36227 30803 36233
rect 30745 36193 30757 36227
rect 30791 36224 30803 36227
rect 32490 36224 32496 36236
rect 30791 36196 31340 36224
rect 32451 36196 32496 36224
rect 30791 36193 30803 36196
rect 30745 36187 30803 36193
rect 31312 36168 31340 36196
rect 32490 36184 32496 36196
rect 32548 36184 32554 36236
rect 33244 36196 35664 36224
rect 29549 36159 29607 36165
rect 29549 36156 29561 36159
rect 29144 36128 29561 36156
rect 29144 36116 29150 36128
rect 29549 36125 29561 36128
rect 29595 36125 29607 36159
rect 29549 36119 29607 36125
rect 29825 36159 29883 36165
rect 29825 36125 29837 36159
rect 29871 36125 29883 36159
rect 29825 36119 29883 36125
rect 30653 36159 30711 36165
rect 30653 36125 30665 36159
rect 30699 36125 30711 36159
rect 30834 36156 30840 36168
rect 30795 36128 30840 36156
rect 30653 36119 30711 36125
rect 22603 36060 28304 36088
rect 28460 36088 28488 36116
rect 29840 36088 29868 36119
rect 30834 36116 30840 36128
rect 30892 36116 30898 36168
rect 31294 36156 31300 36168
rect 31255 36128 31300 36156
rect 31294 36116 31300 36128
rect 31352 36116 31358 36168
rect 32398 36156 32404 36168
rect 32359 36128 32404 36156
rect 32398 36116 32404 36128
rect 32456 36116 32462 36168
rect 28460 36060 29868 36088
rect 30009 36091 30067 36097
rect 22603 36057 22615 36060
rect 22557 36051 22615 36057
rect 30009 36057 30021 36091
rect 30055 36088 30067 36091
rect 33244 36088 33272 36196
rect 33410 36156 33416 36168
rect 33323 36128 33416 36156
rect 33410 36116 33416 36128
rect 33468 36156 33474 36168
rect 34698 36156 34704 36168
rect 33468 36128 34704 36156
rect 33468 36116 33474 36128
rect 34698 36116 34704 36128
rect 34756 36116 34762 36168
rect 30055 36060 33272 36088
rect 30055 36057 30067 36060
rect 30009 36051 30067 36057
rect 1486 36020 1492 36032
rect 1447 35992 1492 36020
rect 1486 35980 1492 35992
rect 1544 35980 1550 36032
rect 8297 36023 8355 36029
rect 8297 35989 8309 36023
rect 8343 36020 8355 36023
rect 8754 36020 8760 36032
rect 8343 35992 8760 36020
rect 8343 35989 8355 35992
rect 8297 35983 8355 35989
rect 8754 35980 8760 35992
rect 8812 35980 8818 36032
rect 23658 35980 23664 36032
rect 23716 36020 23722 36032
rect 24486 36020 24492 36032
rect 23716 35992 24492 36020
rect 23716 35980 23722 35992
rect 24486 35980 24492 35992
rect 24544 35980 24550 36032
rect 29638 36020 29644 36032
rect 29599 35992 29644 36020
rect 29638 35980 29644 35992
rect 29696 35980 29702 36032
rect 31754 35980 31760 36032
rect 31812 36020 31818 36032
rect 33226 36020 33232 36032
rect 31812 35992 31857 36020
rect 33187 35992 33232 36020
rect 31812 35980 31818 35992
rect 33226 35980 33232 35992
rect 33284 35980 33290 36032
rect 33428 36029 33456 36116
rect 33594 36048 33600 36100
rect 33652 36088 33658 36100
rect 35526 36088 35532 36100
rect 33652 36060 33697 36088
rect 35487 36060 35532 36088
rect 33652 36048 33658 36060
rect 35526 36048 35532 36060
rect 35584 36048 35590 36100
rect 35636 36088 35664 36196
rect 36446 36156 36452 36168
rect 36407 36128 36452 36156
rect 36446 36116 36452 36128
rect 36504 36116 36510 36168
rect 37185 36159 37243 36165
rect 37185 36125 37197 36159
rect 37231 36156 37243 36159
rect 37660 36156 37688 36264
rect 38102 36224 38108 36236
rect 38063 36196 38108 36224
rect 38102 36184 38108 36196
rect 38160 36184 38166 36236
rect 38212 36224 38240 36264
rect 39132 36224 39160 36332
rect 41414 36320 41420 36332
rect 41472 36320 41478 36372
rect 47394 36320 47400 36372
rect 47452 36360 47458 36372
rect 48685 36363 48743 36369
rect 48685 36360 48697 36363
rect 47452 36332 48697 36360
rect 47452 36320 47458 36332
rect 48685 36329 48697 36332
rect 48731 36329 48743 36363
rect 48685 36323 48743 36329
rect 39298 36252 39304 36304
rect 39356 36292 39362 36304
rect 46106 36292 46112 36304
rect 39356 36264 46112 36292
rect 39356 36252 39362 36264
rect 46106 36252 46112 36264
rect 46164 36252 46170 36304
rect 41414 36224 41420 36236
rect 38212 36196 39160 36224
rect 41375 36196 41420 36224
rect 41414 36184 41420 36196
rect 41472 36184 41478 36236
rect 49050 36224 49056 36236
rect 49011 36196 49056 36224
rect 49050 36184 49056 36196
rect 49108 36184 49114 36236
rect 38194 36156 38200 36168
rect 37231 36128 37688 36156
rect 38155 36128 38200 36156
rect 37231 36125 37243 36128
rect 37185 36119 37243 36125
rect 38194 36116 38200 36128
rect 38252 36116 38258 36168
rect 38286 36116 38292 36168
rect 38344 36156 38350 36168
rect 39945 36159 40003 36165
rect 39945 36156 39957 36159
rect 38344 36128 39957 36156
rect 38344 36116 38350 36128
rect 39945 36125 39957 36128
rect 39991 36125 40003 36159
rect 40310 36156 40316 36168
rect 40271 36128 40316 36156
rect 39945 36119 40003 36125
rect 40310 36116 40316 36128
rect 40368 36116 40374 36168
rect 42613 36159 42671 36165
rect 42613 36125 42625 36159
rect 42659 36125 42671 36159
rect 42978 36156 42984 36168
rect 42939 36128 42984 36156
rect 42613 36119 42671 36125
rect 41874 36088 41880 36100
rect 35636 36060 41880 36088
rect 41874 36048 41880 36060
rect 41932 36088 41938 36100
rect 42628 36088 42656 36119
rect 42978 36116 42984 36128
rect 43036 36116 43042 36168
rect 47118 36156 47124 36168
rect 47079 36128 47124 36156
rect 47118 36116 47124 36128
rect 47176 36116 47182 36168
rect 47670 36156 47676 36168
rect 47631 36128 47676 36156
rect 47670 36116 47676 36128
rect 47728 36116 47734 36168
rect 48958 36156 48964 36168
rect 48919 36128 48964 36156
rect 48958 36116 48964 36128
rect 49016 36116 49022 36168
rect 58158 36156 58164 36168
rect 58119 36128 58164 36156
rect 58158 36116 58164 36128
rect 58216 36116 58222 36168
rect 41932 36060 42656 36088
rect 44453 36091 44511 36097
rect 41932 36048 41938 36060
rect 44453 36057 44465 36091
rect 44499 36088 44511 36091
rect 44634 36088 44640 36100
rect 44499 36060 44640 36088
rect 44499 36057 44511 36060
rect 44453 36051 44511 36057
rect 44634 36048 44640 36060
rect 44692 36048 44698 36100
rect 46566 36048 46572 36100
rect 46624 36048 46630 36100
rect 57790 36048 57796 36100
rect 57848 36088 57854 36100
rect 57885 36091 57943 36097
rect 57885 36088 57897 36091
rect 57848 36060 57897 36088
rect 57848 36048 57854 36060
rect 57885 36057 57897 36060
rect 57931 36057 57943 36091
rect 57885 36051 57943 36057
rect 33397 36023 33456 36029
rect 33397 35989 33409 36023
rect 33443 35992 33456 36023
rect 39114 36020 39120 36032
rect 39075 35992 39120 36020
rect 33443 35989 33455 35992
rect 33397 35983 33455 35989
rect 39114 35980 39120 35992
rect 39172 36020 39178 36032
rect 40126 36020 40132 36032
rect 39172 35992 40132 36020
rect 39172 35980 39178 35992
rect 40126 35980 40132 35992
rect 40184 35980 40190 36032
rect 1104 35930 58880 35952
rect 1104 35878 19574 35930
rect 19626 35878 19638 35930
rect 19690 35878 19702 35930
rect 19754 35878 19766 35930
rect 19818 35878 19830 35930
rect 19882 35878 50294 35930
rect 50346 35878 50358 35930
rect 50410 35878 50422 35930
rect 50474 35878 50486 35930
rect 50538 35878 50550 35930
rect 50602 35878 58880 35930
rect 1104 35856 58880 35878
rect 6638 35816 6644 35828
rect 6599 35788 6644 35816
rect 6638 35776 6644 35788
rect 6696 35776 6702 35828
rect 6730 35776 6736 35828
rect 6788 35816 6794 35828
rect 8849 35819 8907 35825
rect 8849 35816 8861 35819
rect 6788 35788 8861 35816
rect 6788 35776 6794 35788
rect 8849 35785 8861 35788
rect 8895 35785 8907 35819
rect 8849 35779 8907 35785
rect 16574 35776 16580 35828
rect 16632 35816 16638 35828
rect 17770 35816 17776 35828
rect 16632 35788 17776 35816
rect 16632 35776 16638 35788
rect 17770 35776 17776 35788
rect 17828 35816 17834 35828
rect 28471 35819 28529 35825
rect 17828 35788 26924 35816
rect 17828 35776 17834 35788
rect 6549 35751 6607 35757
rect 6549 35717 6561 35751
rect 6595 35748 6607 35751
rect 7006 35748 7012 35760
rect 6595 35720 7012 35748
rect 6595 35717 6607 35720
rect 6549 35711 6607 35717
rect 7006 35708 7012 35720
rect 7064 35748 7070 35760
rect 7466 35748 7472 35760
rect 7064 35720 7472 35748
rect 7064 35708 7070 35720
rect 7466 35708 7472 35720
rect 7524 35708 7530 35760
rect 8018 35748 8024 35760
rect 7979 35720 8024 35748
rect 8018 35708 8024 35720
rect 8076 35708 8082 35760
rect 9953 35751 10011 35757
rect 9953 35748 9965 35751
rect 8128 35720 9965 35748
rect 8128 35692 8156 35720
rect 9953 35717 9965 35720
rect 9999 35717 10011 35751
rect 9953 35711 10011 35717
rect 18138 35708 18144 35760
rect 18196 35748 18202 35760
rect 19153 35751 19211 35757
rect 19153 35748 19165 35751
rect 18196 35720 19165 35748
rect 18196 35708 18202 35720
rect 19153 35717 19165 35720
rect 19199 35748 19211 35751
rect 19242 35748 19248 35760
rect 19199 35720 19248 35748
rect 19199 35717 19211 35720
rect 19153 35711 19211 35717
rect 19242 35708 19248 35720
rect 19300 35748 19306 35760
rect 19300 35720 19748 35748
rect 19300 35708 19306 35720
rect 6917 35683 6975 35689
rect 6917 35649 6929 35683
rect 6963 35680 6975 35683
rect 7742 35680 7748 35692
rect 6963 35652 7748 35680
rect 6963 35649 6975 35652
rect 6917 35643 6975 35649
rect 7742 35640 7748 35652
rect 7800 35640 7806 35692
rect 7929 35683 7987 35689
rect 7929 35649 7941 35683
rect 7975 35649 7987 35683
rect 8110 35680 8116 35692
rect 8071 35652 8116 35680
rect 7929 35643 7987 35649
rect 7944 35612 7972 35643
rect 8110 35640 8116 35652
rect 8168 35640 8174 35692
rect 8294 35680 8300 35692
rect 8255 35652 8300 35680
rect 8294 35640 8300 35652
rect 8352 35640 8358 35692
rect 8754 35680 8760 35692
rect 8715 35652 8760 35680
rect 8754 35640 8760 35652
rect 8812 35640 8818 35692
rect 8938 35680 8944 35692
rect 8899 35652 8944 35680
rect 8938 35640 8944 35652
rect 8996 35640 9002 35692
rect 11698 35680 11704 35692
rect 11659 35652 11704 35680
rect 11698 35640 11704 35652
rect 11756 35640 11762 35692
rect 11882 35680 11888 35692
rect 11843 35652 11888 35680
rect 11882 35640 11888 35652
rect 11940 35640 11946 35692
rect 19720 35689 19748 35720
rect 22094 35708 22100 35760
rect 22152 35748 22158 35760
rect 23201 35751 23259 35757
rect 23201 35748 23213 35751
rect 22152 35720 23213 35748
rect 22152 35708 22158 35720
rect 23201 35717 23213 35720
rect 23247 35717 23259 35751
rect 23201 35711 23259 35717
rect 23385 35751 23443 35757
rect 23385 35717 23397 35751
rect 23431 35748 23443 35751
rect 23842 35748 23848 35760
rect 23431 35720 23848 35748
rect 23431 35717 23443 35720
rect 23385 35711 23443 35717
rect 23842 35708 23848 35720
rect 23900 35708 23906 35760
rect 18785 35683 18843 35689
rect 18785 35649 18797 35683
rect 18831 35649 18843 35683
rect 18785 35643 18843 35649
rect 19613 35683 19671 35689
rect 19613 35649 19625 35683
rect 19659 35649 19671 35683
rect 19613 35643 19671 35649
rect 19705 35683 19763 35689
rect 19705 35649 19717 35683
rect 19751 35649 19763 35683
rect 19705 35643 19763 35649
rect 8846 35612 8852 35624
rect 7944 35584 8852 35612
rect 8846 35572 8852 35584
rect 8904 35572 8910 35624
rect 18693 35615 18751 35621
rect 18693 35581 18705 35615
rect 18739 35581 18751 35615
rect 18800 35612 18828 35643
rect 19334 35612 19340 35624
rect 18800 35584 19340 35612
rect 18693 35575 18751 35581
rect 5534 35504 5540 35556
rect 5592 35544 5598 35556
rect 6365 35547 6423 35553
rect 6365 35544 6377 35547
rect 5592 35516 6377 35544
rect 5592 35504 5598 35516
rect 6365 35513 6377 35516
rect 6411 35513 6423 35547
rect 6365 35507 6423 35513
rect 11977 35547 12035 35553
rect 11977 35513 11989 35547
rect 12023 35544 12035 35547
rect 12342 35544 12348 35556
rect 12023 35516 12348 35544
rect 12023 35513 12035 35516
rect 11977 35507 12035 35513
rect 12342 35504 12348 35516
rect 12400 35504 12406 35556
rect 18708 35488 18736 35575
rect 19334 35572 19340 35584
rect 19392 35612 19398 35624
rect 19628 35612 19656 35643
rect 21082 35640 21088 35692
rect 21140 35680 21146 35692
rect 23017 35683 23075 35689
rect 23017 35680 23029 35683
rect 21140 35652 23029 35680
rect 21140 35640 21146 35652
rect 23017 35649 23029 35652
rect 23063 35649 23075 35683
rect 26896 35680 26924 35788
rect 28471 35785 28483 35819
rect 28517 35816 28529 35819
rect 28718 35816 28724 35828
rect 28517 35788 28724 35816
rect 28517 35785 28529 35788
rect 28471 35779 28529 35785
rect 28718 35776 28724 35788
rect 28776 35816 28782 35828
rect 29089 35819 29147 35825
rect 29089 35816 29101 35819
rect 28776 35788 29101 35816
rect 28776 35776 28782 35788
rect 29089 35785 29101 35788
rect 29135 35785 29147 35819
rect 29089 35779 29147 35785
rect 32769 35819 32827 35825
rect 32769 35785 32781 35819
rect 32815 35816 32827 35819
rect 38194 35816 38200 35828
rect 32815 35788 38200 35816
rect 32815 35785 32827 35788
rect 32769 35779 32827 35785
rect 38194 35776 38200 35788
rect 38252 35776 38258 35828
rect 40126 35816 40132 35828
rect 40087 35788 40132 35816
rect 40126 35776 40132 35788
rect 40184 35776 40190 35828
rect 46109 35819 46167 35825
rect 46109 35785 46121 35819
rect 46155 35816 46167 35819
rect 47118 35816 47124 35828
rect 46155 35788 47124 35816
rect 46155 35785 46167 35788
rect 46109 35779 46167 35785
rect 47118 35776 47124 35788
rect 47176 35776 47182 35828
rect 49050 35776 49056 35828
rect 49108 35816 49114 35828
rect 49237 35819 49295 35825
rect 49237 35816 49249 35819
rect 49108 35788 49249 35816
rect 49108 35776 49114 35788
rect 49237 35785 49249 35788
rect 49283 35785 49295 35819
rect 58158 35816 58164 35828
rect 58119 35788 58164 35816
rect 49237 35779 49295 35785
rect 58158 35776 58164 35788
rect 58216 35776 58222 35828
rect 27982 35708 27988 35760
rect 28040 35748 28046 35760
rect 28261 35751 28319 35757
rect 28261 35748 28273 35751
rect 28040 35720 28273 35748
rect 28040 35708 28046 35720
rect 28261 35717 28273 35720
rect 28307 35717 28319 35751
rect 50706 35748 50712 35760
rect 28261 35711 28319 35717
rect 28552 35720 50712 35748
rect 28552 35680 28580 35720
rect 50706 35708 50712 35720
rect 50764 35708 50770 35760
rect 26896 35652 28580 35680
rect 29457 35683 29515 35689
rect 23017 35643 23075 35649
rect 29457 35649 29469 35683
rect 29503 35680 29515 35683
rect 29638 35680 29644 35692
rect 29503 35652 29644 35680
rect 29503 35649 29515 35652
rect 29457 35643 29515 35649
rect 29638 35640 29644 35652
rect 29696 35680 29702 35692
rect 30190 35680 30196 35692
rect 29696 35652 30196 35680
rect 29696 35640 29702 35652
rect 30190 35640 30196 35652
rect 30248 35640 30254 35692
rect 31754 35640 31760 35692
rect 31812 35680 31818 35692
rect 32309 35683 32367 35689
rect 32309 35680 32321 35683
rect 31812 35652 32321 35680
rect 31812 35640 31818 35652
rect 32309 35649 32321 35652
rect 32355 35649 32367 35683
rect 32309 35643 32367 35649
rect 32398 35640 32404 35692
rect 32456 35680 32462 35692
rect 32493 35683 32551 35689
rect 32493 35680 32505 35683
rect 32456 35652 32505 35680
rect 32456 35640 32462 35652
rect 32493 35649 32505 35652
rect 32539 35649 32551 35683
rect 32493 35643 32551 35649
rect 32861 35683 32919 35689
rect 32861 35649 32873 35683
rect 32907 35680 32919 35683
rect 33226 35680 33232 35692
rect 32907 35652 33232 35680
rect 32907 35649 32919 35652
rect 32861 35643 32919 35649
rect 33226 35640 33232 35652
rect 33284 35640 33290 35692
rect 45094 35640 45100 35692
rect 45152 35680 45158 35692
rect 45281 35683 45339 35689
rect 45281 35680 45293 35683
rect 45152 35652 45293 35680
rect 45152 35640 45158 35652
rect 45281 35649 45293 35652
rect 45327 35649 45339 35683
rect 45281 35643 45339 35649
rect 49237 35683 49295 35689
rect 49237 35649 49249 35683
rect 49283 35649 49295 35683
rect 49418 35680 49424 35692
rect 49379 35652 49424 35680
rect 49237 35643 49295 35649
rect 24946 35612 24952 35624
rect 19392 35584 19656 35612
rect 19904 35584 24952 35612
rect 19392 35572 19398 35584
rect 19061 35547 19119 35553
rect 19061 35513 19073 35547
rect 19107 35544 19119 35547
rect 19904 35544 19932 35584
rect 24946 35572 24952 35584
rect 25004 35572 25010 35624
rect 29086 35572 29092 35624
rect 29144 35612 29150 35624
rect 29365 35615 29423 35621
rect 29365 35612 29377 35615
rect 29144 35584 29377 35612
rect 29144 35572 29150 35584
rect 29365 35581 29377 35584
rect 29411 35581 29423 35615
rect 29365 35575 29423 35581
rect 43622 35572 43628 35624
rect 43680 35612 43686 35624
rect 45189 35615 45247 35621
rect 45189 35612 45201 35615
rect 43680 35584 45201 35612
rect 43680 35572 43686 35584
rect 45189 35581 45201 35584
rect 45235 35581 45247 35615
rect 49252 35612 49280 35643
rect 49418 35640 49424 35652
rect 49476 35640 49482 35692
rect 49970 35612 49976 35624
rect 49252 35584 49976 35612
rect 45189 35575 45247 35581
rect 49970 35572 49976 35584
rect 50028 35572 50034 35624
rect 19107 35516 19932 35544
rect 19981 35547 20039 35553
rect 19107 35513 19119 35516
rect 19061 35507 19119 35513
rect 19981 35513 19993 35547
rect 20027 35544 20039 35547
rect 23658 35544 23664 35556
rect 20027 35516 23664 35544
rect 20027 35513 20039 35516
rect 19981 35507 20039 35513
rect 23658 35504 23664 35516
rect 23716 35504 23722 35556
rect 28626 35544 28632 35556
rect 28587 35516 28632 35544
rect 28626 35504 28632 35516
rect 28684 35504 28690 35556
rect 7745 35479 7803 35485
rect 7745 35445 7757 35479
rect 7791 35476 7803 35479
rect 7926 35476 7932 35488
rect 7791 35448 7932 35476
rect 7791 35445 7803 35448
rect 7745 35439 7803 35445
rect 7926 35436 7932 35448
rect 7984 35436 7990 35488
rect 8846 35436 8852 35488
rect 8904 35476 8910 35488
rect 9401 35479 9459 35485
rect 9401 35476 9413 35479
rect 8904 35448 9413 35476
rect 8904 35436 8910 35448
rect 9401 35445 9413 35448
rect 9447 35445 9459 35479
rect 9401 35439 9459 35445
rect 12434 35436 12440 35488
rect 12492 35476 12498 35488
rect 12529 35479 12587 35485
rect 12529 35476 12541 35479
rect 12492 35448 12541 35476
rect 12492 35436 12498 35448
rect 12529 35445 12541 35448
rect 12575 35445 12587 35479
rect 18690 35476 18696 35488
rect 18603 35448 18696 35476
rect 12529 35439 12587 35445
rect 18690 35436 18696 35448
rect 18748 35476 18754 35488
rect 19797 35479 19855 35485
rect 19797 35476 19809 35479
rect 18748 35448 19809 35476
rect 18748 35436 18754 35448
rect 19797 35445 19809 35448
rect 19843 35476 19855 35479
rect 20070 35476 20076 35488
rect 19843 35448 20076 35476
rect 19843 35445 19855 35448
rect 19797 35439 19855 35445
rect 20070 35436 20076 35448
rect 20128 35436 20134 35488
rect 28350 35436 28356 35488
rect 28408 35476 28414 35488
rect 28445 35479 28503 35485
rect 28445 35476 28457 35479
rect 28408 35448 28457 35476
rect 28408 35436 28414 35448
rect 28445 35445 28457 35448
rect 28491 35445 28503 35479
rect 30190 35476 30196 35488
rect 30151 35448 30196 35476
rect 28445 35439 28503 35445
rect 30190 35436 30196 35448
rect 30248 35436 30254 35488
rect 41046 35476 41052 35488
rect 41007 35448 41052 35476
rect 41046 35436 41052 35448
rect 41104 35436 41110 35488
rect 1104 35386 58880 35408
rect 1104 35334 4214 35386
rect 4266 35334 4278 35386
rect 4330 35334 4342 35386
rect 4394 35334 4406 35386
rect 4458 35334 4470 35386
rect 4522 35334 34934 35386
rect 34986 35334 34998 35386
rect 35050 35334 35062 35386
rect 35114 35334 35126 35386
rect 35178 35334 35190 35386
rect 35242 35334 58880 35386
rect 1104 35312 58880 35334
rect 6733 35275 6791 35281
rect 6733 35241 6745 35275
rect 6779 35272 6791 35275
rect 7006 35272 7012 35284
rect 6779 35244 7012 35272
rect 6779 35241 6791 35244
rect 6733 35235 6791 35241
rect 7006 35232 7012 35244
rect 7064 35232 7070 35284
rect 7742 35272 7748 35284
rect 7703 35244 7748 35272
rect 7742 35232 7748 35244
rect 7800 35232 7806 35284
rect 9033 35275 9091 35281
rect 9033 35241 9045 35275
rect 9079 35272 9091 35275
rect 9582 35272 9588 35284
rect 9079 35244 9588 35272
rect 9079 35241 9091 35244
rect 9033 35235 9091 35241
rect 7006 35136 7012 35148
rect 6967 35108 7012 35136
rect 7006 35096 7012 35108
rect 7064 35096 7070 35148
rect 8205 35139 8263 35145
rect 8205 35136 8217 35139
rect 7116 35108 8217 35136
rect 7116 35077 7144 35108
rect 8205 35105 8217 35108
rect 8251 35136 8263 35139
rect 8294 35136 8300 35148
rect 8251 35108 8300 35136
rect 8251 35105 8263 35108
rect 8205 35099 8263 35105
rect 8294 35096 8300 35108
rect 8352 35136 8358 35148
rect 9048 35136 9076 35235
rect 9582 35232 9588 35244
rect 9640 35232 9646 35284
rect 11701 35275 11759 35281
rect 11701 35241 11713 35275
rect 11747 35272 11759 35275
rect 11882 35272 11888 35284
rect 11747 35244 11888 35272
rect 11747 35241 11759 35244
rect 11701 35235 11759 35241
rect 11882 35232 11888 35244
rect 11940 35232 11946 35284
rect 16574 35272 16580 35284
rect 16535 35244 16580 35272
rect 16574 35232 16580 35244
rect 16632 35232 16638 35284
rect 18322 35232 18328 35284
rect 18380 35272 18386 35284
rect 18509 35275 18567 35281
rect 18509 35272 18521 35275
rect 18380 35244 18521 35272
rect 18380 35232 18386 35244
rect 18509 35241 18521 35244
rect 18555 35241 18567 35275
rect 18690 35272 18696 35284
rect 18651 35244 18696 35272
rect 18509 35235 18567 35241
rect 18690 35232 18696 35244
rect 18748 35232 18754 35284
rect 22094 35232 22100 35284
rect 22152 35272 22158 35284
rect 22281 35275 22339 35281
rect 22281 35272 22293 35275
rect 22152 35244 22293 35272
rect 22152 35232 22158 35244
rect 22281 35241 22293 35244
rect 22327 35272 22339 35275
rect 25225 35275 25283 35281
rect 22327 35244 23612 35272
rect 22327 35241 22339 35244
rect 22281 35235 22339 35241
rect 22373 35207 22431 35213
rect 22373 35204 22385 35207
rect 21100 35176 22385 35204
rect 8352 35108 9076 35136
rect 10873 35139 10931 35145
rect 8352 35096 8358 35108
rect 10873 35105 10885 35139
rect 10919 35136 10931 35139
rect 11333 35139 11391 35145
rect 11333 35136 11345 35139
rect 10919 35108 11345 35136
rect 10919 35105 10931 35108
rect 10873 35099 10931 35105
rect 11333 35105 11345 35108
rect 11379 35136 11391 35139
rect 12434 35136 12440 35148
rect 11379 35108 12440 35136
rect 11379 35105 11391 35108
rect 11333 35099 11391 35105
rect 12434 35096 12440 35108
rect 12492 35136 12498 35148
rect 12492 35108 13308 35136
rect 12492 35096 12498 35108
rect 7101 35071 7159 35077
rect 7101 35037 7113 35071
rect 7147 35037 7159 35071
rect 7926 35068 7932 35080
rect 7887 35040 7932 35068
rect 7101 35031 7159 35037
rect 7926 35028 7932 35040
rect 7984 35028 7990 35080
rect 8018 35028 8024 35080
rect 8076 35068 8082 35080
rect 8113 35071 8171 35077
rect 8113 35068 8125 35071
rect 8076 35040 8125 35068
rect 8076 35028 8082 35040
rect 8113 35037 8125 35040
rect 8159 35037 8171 35071
rect 11514 35068 11520 35080
rect 11475 35040 11520 35068
rect 8113 35031 8171 35037
rect 11514 35028 11520 35040
rect 11572 35028 11578 35080
rect 12158 35068 12164 35080
rect 12119 35040 12164 35068
rect 12158 35028 12164 35040
rect 12216 35028 12222 35080
rect 12529 35071 12587 35077
rect 12529 35037 12541 35071
rect 12575 35037 12587 35071
rect 12710 35068 12716 35080
rect 12671 35040 12716 35068
rect 12529 35031 12587 35037
rect 12544 35000 12572 35031
rect 12710 35028 12716 35040
rect 12768 35028 12774 35080
rect 13280 35077 13308 35108
rect 13265 35071 13323 35077
rect 13265 35037 13277 35071
rect 13311 35068 13323 35071
rect 16025 35071 16083 35077
rect 16025 35068 16037 35071
rect 13311 35040 16037 35068
rect 13311 35037 13323 35040
rect 13265 35031 13323 35037
rect 16025 35037 16037 35040
rect 16071 35068 16083 35071
rect 17129 35071 17187 35077
rect 17129 35068 17141 35071
rect 16071 35040 17141 35068
rect 16071 35037 16083 35040
rect 16025 35031 16083 35037
rect 17129 35037 17141 35040
rect 17175 35068 17187 35071
rect 17175 35040 18828 35068
rect 17175 35037 17187 35040
rect 17129 35031 17187 35037
rect 12894 35000 12900 35012
rect 12544 34972 12900 35000
rect 12894 34960 12900 34972
rect 12952 35000 12958 35012
rect 15657 35003 15715 35009
rect 15657 35000 15669 35003
rect 12952 34972 15669 35000
rect 12952 34960 12958 34972
rect 15657 34969 15669 34972
rect 15703 34969 15715 35003
rect 15657 34963 15715 34969
rect 15841 35003 15899 35009
rect 15841 34969 15853 35003
rect 15887 35000 15899 35003
rect 16574 35000 16580 35012
rect 15887 34972 16580 35000
rect 15887 34969 15899 34972
rect 15841 34963 15899 34969
rect 16574 34960 16580 34972
rect 16632 34960 16638 35012
rect 17862 34960 17868 35012
rect 17920 35000 17926 35012
rect 18325 35003 18383 35009
rect 18325 35000 18337 35003
rect 17920 34972 18337 35000
rect 17920 34960 17926 34972
rect 18325 34969 18337 34972
rect 18371 34969 18383 35003
rect 18325 34963 18383 34969
rect 12526 34932 12532 34944
rect 12487 34904 12532 34932
rect 12526 34892 12532 34904
rect 12584 34892 12590 34944
rect 18414 34892 18420 34944
rect 18472 34932 18478 34944
rect 18525 34935 18583 34941
rect 18525 34932 18537 34935
rect 18472 34904 18537 34932
rect 18472 34892 18478 34904
rect 18525 34901 18537 34904
rect 18571 34901 18583 34935
rect 18800 34932 18828 35040
rect 20806 35028 20812 35080
rect 20864 35068 20870 35080
rect 21100 35077 21128 35176
rect 22373 35173 22385 35176
rect 22419 35173 22431 35207
rect 22373 35167 22431 35173
rect 21085 35071 21143 35077
rect 21085 35068 21097 35071
rect 20864 35040 21097 35068
rect 20864 35028 20870 35040
rect 21085 35037 21097 35040
rect 21131 35037 21143 35071
rect 21085 35031 21143 35037
rect 21545 35071 21603 35077
rect 21545 35037 21557 35071
rect 21591 35037 21603 35071
rect 23474 35068 23480 35080
rect 23435 35040 23480 35068
rect 21545 35031 21603 35037
rect 20717 35003 20775 35009
rect 20717 34969 20729 35003
rect 20763 35000 20775 35003
rect 21266 35000 21272 35012
rect 20763 34972 21272 35000
rect 20763 34969 20775 34972
rect 20717 34963 20775 34969
rect 21266 34960 21272 34972
rect 21324 34960 21330 35012
rect 21560 35000 21588 35031
rect 23474 35028 23480 35040
rect 23532 35028 23538 35080
rect 23584 35068 23612 35244
rect 25225 35241 25237 35275
rect 25271 35272 25283 35275
rect 27890 35272 27896 35284
rect 25271 35244 27896 35272
rect 25271 35241 25283 35244
rect 25225 35235 25283 35241
rect 27890 35232 27896 35244
rect 27948 35232 27954 35284
rect 28442 35232 28448 35284
rect 28500 35272 28506 35284
rect 28629 35275 28687 35281
rect 28629 35272 28641 35275
rect 28500 35244 28641 35272
rect 28500 35232 28506 35244
rect 28629 35241 28641 35244
rect 28675 35241 28687 35275
rect 28629 35235 28687 35241
rect 32582 35232 32588 35284
rect 32640 35272 32646 35284
rect 32640 35244 35940 35272
rect 32640 35232 32646 35244
rect 24486 35164 24492 35216
rect 24544 35204 24550 35216
rect 34698 35204 34704 35216
rect 24544 35176 25452 35204
rect 34659 35176 34704 35204
rect 24544 35164 24550 35176
rect 23661 35071 23719 35077
rect 23661 35068 23673 35071
rect 23584 35040 23673 35068
rect 23661 35037 23673 35040
rect 23707 35037 23719 35071
rect 25130 35068 25136 35080
rect 25091 35040 25136 35068
rect 23661 35031 23719 35037
rect 25130 35028 25136 35040
rect 25188 35028 25194 35080
rect 25424 35077 25452 35176
rect 34698 35164 34704 35176
rect 34756 35164 34762 35216
rect 35912 35204 35940 35244
rect 35986 35232 35992 35284
rect 36044 35272 36050 35284
rect 37366 35272 37372 35284
rect 36044 35244 37372 35272
rect 36044 35232 36050 35244
rect 37366 35232 37372 35244
rect 37424 35272 37430 35284
rect 37461 35275 37519 35281
rect 37461 35272 37473 35275
rect 37424 35244 37473 35272
rect 37424 35232 37430 35244
rect 37461 35241 37473 35244
rect 37507 35241 37519 35275
rect 43622 35272 43628 35284
rect 43583 35244 43628 35272
rect 37461 35235 37519 35241
rect 43622 35232 43628 35244
rect 43680 35232 43686 35284
rect 53561 35207 53619 35213
rect 35912 35176 45554 35204
rect 35161 35139 35219 35145
rect 25516 35108 28580 35136
rect 25409 35071 25467 35077
rect 25409 35037 25421 35071
rect 25455 35037 25467 35071
rect 25409 35031 25467 35037
rect 22646 35000 22652 35012
rect 21560 34972 22652 35000
rect 22646 34960 22652 34972
rect 22704 35000 22710 35012
rect 22741 35003 22799 35009
rect 22741 35000 22753 35003
rect 22704 34972 22753 35000
rect 22704 34960 22710 34972
rect 22741 34969 22753 34972
rect 22787 34969 22799 35003
rect 22741 34963 22799 34969
rect 23845 35003 23903 35009
rect 23845 34969 23857 35003
rect 23891 35000 23903 35003
rect 25516 35000 25544 35108
rect 25593 35071 25651 35077
rect 25593 35037 25605 35071
rect 25639 35037 25651 35071
rect 28350 35068 28356 35080
rect 28311 35040 28356 35068
rect 25593 35031 25651 35037
rect 23891 34972 25544 35000
rect 23891 34969 23903 34972
rect 23845 34963 23903 34969
rect 22186 34932 22192 34944
rect 18800 34904 22192 34932
rect 18525 34895 18583 34901
rect 22186 34892 22192 34904
rect 22244 34892 22250 34944
rect 24946 34892 24952 34944
rect 25004 34932 25010 34944
rect 25608 34932 25636 35031
rect 28350 35028 28356 35040
rect 28408 35028 28414 35080
rect 25004 34904 25636 34932
rect 25004 34892 25010 34904
rect 27982 34892 27988 34944
rect 28040 34932 28046 34944
rect 28445 34935 28503 34941
rect 28445 34932 28457 34935
rect 28040 34904 28457 34932
rect 28040 34892 28046 34904
rect 28445 34901 28457 34904
rect 28491 34901 28503 34935
rect 28552 34932 28580 35108
rect 35161 35105 35173 35139
rect 35207 35136 35219 35139
rect 35894 35136 35900 35148
rect 35207 35108 35900 35136
rect 35207 35105 35219 35108
rect 35161 35099 35219 35105
rect 35894 35096 35900 35108
rect 35952 35096 35958 35148
rect 37182 35096 37188 35148
rect 37240 35136 37246 35148
rect 37553 35139 37611 35145
rect 37553 35136 37565 35139
rect 37240 35108 37565 35136
rect 37240 35096 37246 35108
rect 37553 35105 37565 35108
rect 37599 35105 37611 35139
rect 43254 35136 43260 35148
rect 43215 35108 43260 35136
rect 37553 35099 37611 35105
rect 43254 35096 43260 35108
rect 43312 35096 43318 35148
rect 45526 35136 45554 35176
rect 53561 35173 53573 35207
rect 53607 35204 53619 35207
rect 54202 35204 54208 35216
rect 53607 35176 54208 35204
rect 53607 35173 53619 35176
rect 53561 35167 53619 35173
rect 54202 35164 54208 35176
rect 54260 35164 54266 35216
rect 47581 35139 47639 35145
rect 47581 35136 47593 35139
rect 45526 35108 47593 35136
rect 47581 35105 47593 35108
rect 47627 35105 47639 35139
rect 49510 35136 49516 35148
rect 47581 35099 47639 35105
rect 48608 35108 49516 35136
rect 48504 35080 48556 35086
rect 28629 35071 28687 35077
rect 28629 35037 28641 35071
rect 28675 35068 28687 35071
rect 28718 35068 28724 35080
rect 28675 35040 28724 35068
rect 28675 35037 28687 35040
rect 28629 35031 28687 35037
rect 28718 35028 28724 35040
rect 28776 35028 28782 35080
rect 35069 35071 35127 35077
rect 35069 35037 35081 35071
rect 35115 35068 35127 35071
rect 35342 35068 35348 35080
rect 35115 35040 35348 35068
rect 35115 35037 35127 35040
rect 35069 35031 35127 35037
rect 35342 35028 35348 35040
rect 35400 35028 35406 35080
rect 37458 35068 37464 35080
rect 37419 35040 37464 35068
rect 37458 35028 37464 35040
rect 37516 35028 37522 35080
rect 43346 35068 43352 35080
rect 43307 35040 43352 35068
rect 43346 35028 43352 35040
rect 43404 35028 43410 35080
rect 48608 35077 48636 35108
rect 49510 35096 49516 35108
rect 49568 35096 49574 35148
rect 52178 35096 52184 35148
rect 52236 35136 52242 35148
rect 53101 35139 53159 35145
rect 53101 35136 53113 35139
rect 52236 35108 53113 35136
rect 52236 35096 52242 35108
rect 53101 35105 53113 35108
rect 53147 35105 53159 35139
rect 57882 35136 57888 35148
rect 57843 35108 57888 35136
rect 53101 35099 53159 35105
rect 57882 35096 57888 35108
rect 57940 35096 57946 35148
rect 48593 35071 48651 35077
rect 48593 35037 48605 35071
rect 48639 35037 48651 35071
rect 48593 35031 48651 35037
rect 48504 35022 48556 35028
rect 28902 34960 28908 35012
rect 28960 35000 28966 35012
rect 40310 35000 40316 35012
rect 28960 34972 40316 35000
rect 28960 34960 28966 34972
rect 40310 34960 40316 34972
rect 40368 34960 40374 35012
rect 35986 34932 35992 34944
rect 28552 34904 35992 34932
rect 28445 34895 28503 34901
rect 35986 34892 35992 34904
rect 36044 34892 36050 34944
rect 37829 34935 37887 34941
rect 37829 34901 37841 34935
rect 37875 34932 37887 34935
rect 38930 34932 38936 34944
rect 37875 34904 38936 34932
rect 37875 34901 37887 34904
rect 37829 34895 37887 34901
rect 38930 34892 38936 34904
rect 38988 34892 38994 34944
rect 48406 34892 48412 34944
rect 48464 34932 48470 34944
rect 48608 34932 48636 35031
rect 49050 35028 49056 35080
rect 49108 35068 49114 35080
rect 49145 35071 49203 35077
rect 49145 35068 49157 35071
rect 49108 35040 49157 35068
rect 49108 35028 49114 35040
rect 49145 35037 49157 35040
rect 49191 35037 49203 35071
rect 49145 35031 49203 35037
rect 49329 35071 49387 35077
rect 49329 35037 49341 35071
rect 49375 35037 49387 35071
rect 49329 35031 49387 35037
rect 53193 35071 53251 35077
rect 53193 35037 53205 35071
rect 53239 35068 53251 35071
rect 53558 35068 53564 35080
rect 53239 35040 53564 35068
rect 53239 35037 53251 35040
rect 53193 35031 53251 35037
rect 48682 34960 48688 35012
rect 48740 35000 48746 35012
rect 49344 35000 49372 35031
rect 53558 35028 53564 35040
rect 53616 35028 53622 35080
rect 58158 35068 58164 35080
rect 58119 35040 58164 35068
rect 58158 35028 58164 35040
rect 58216 35028 58222 35080
rect 50157 35003 50215 35009
rect 50157 35000 50169 35003
rect 48740 34972 50169 35000
rect 48740 34960 48746 34972
rect 50157 34969 50169 34972
rect 50203 34969 50215 35003
rect 50157 34963 50215 34969
rect 48464 34904 48636 34932
rect 49329 34935 49387 34941
rect 48464 34892 48470 34904
rect 49329 34901 49341 34935
rect 49375 34932 49387 34935
rect 49970 34932 49976 34944
rect 49375 34904 49976 34932
rect 49375 34901 49387 34904
rect 49329 34895 49387 34901
rect 49970 34892 49976 34904
rect 50028 34892 50034 34944
rect 1104 34842 58880 34864
rect 1104 34790 19574 34842
rect 19626 34790 19638 34842
rect 19690 34790 19702 34842
rect 19754 34790 19766 34842
rect 19818 34790 19830 34842
rect 19882 34790 50294 34842
rect 50346 34790 50358 34842
rect 50410 34790 50422 34842
rect 50474 34790 50486 34842
rect 50538 34790 50550 34842
rect 50602 34790 58880 34842
rect 1104 34768 58880 34790
rect 8294 34688 8300 34740
rect 8352 34728 8358 34740
rect 8481 34731 8539 34737
rect 8481 34728 8493 34731
rect 8352 34700 8493 34728
rect 8352 34688 8358 34700
rect 8481 34697 8493 34700
rect 8527 34697 8539 34731
rect 8481 34691 8539 34697
rect 16853 34731 16911 34737
rect 16853 34697 16865 34731
rect 16899 34728 16911 34731
rect 18138 34728 18144 34740
rect 16899 34700 18144 34728
rect 16899 34697 16911 34700
rect 16853 34691 16911 34697
rect 18138 34688 18144 34700
rect 18196 34688 18202 34740
rect 18239 34731 18297 34737
rect 18239 34697 18251 34731
rect 18285 34728 18297 34731
rect 19334 34728 19340 34740
rect 18285 34700 19340 34728
rect 18285 34697 18297 34700
rect 18239 34691 18297 34697
rect 19334 34688 19340 34700
rect 19392 34688 19398 34740
rect 20257 34731 20315 34737
rect 20257 34697 20269 34731
rect 20303 34728 20315 34731
rect 20806 34728 20812 34740
rect 20303 34700 20812 34728
rect 20303 34697 20315 34700
rect 20257 34691 20315 34697
rect 20806 34688 20812 34700
rect 20864 34688 20870 34740
rect 21082 34728 21088 34740
rect 21043 34700 21088 34728
rect 21082 34688 21088 34700
rect 21140 34688 21146 34740
rect 22186 34688 22192 34740
rect 22244 34728 22250 34740
rect 48590 34728 48596 34740
rect 22244 34700 48596 34728
rect 22244 34688 22250 34700
rect 48590 34688 48596 34700
rect 48648 34688 48654 34740
rect 48777 34731 48835 34737
rect 48777 34697 48789 34731
rect 48823 34728 48835 34731
rect 48958 34728 48964 34740
rect 48823 34700 48964 34728
rect 48823 34697 48835 34700
rect 48777 34691 48835 34697
rect 48958 34688 48964 34700
rect 49016 34688 49022 34740
rect 52178 34728 52184 34740
rect 52139 34700 52184 34728
rect 52178 34688 52184 34700
rect 52236 34688 52242 34740
rect 53558 34728 53564 34740
rect 53519 34700 53564 34728
rect 53558 34688 53564 34700
rect 53616 34688 53622 34740
rect 58158 34728 58164 34740
rect 58119 34700 58164 34728
rect 58158 34688 58164 34700
rect 58216 34688 58222 34740
rect 10781 34663 10839 34669
rect 10781 34629 10793 34663
rect 10827 34660 10839 34663
rect 11701 34663 11759 34669
rect 11701 34660 11713 34663
rect 10827 34632 11713 34660
rect 10827 34629 10839 34632
rect 10781 34623 10839 34629
rect 11701 34629 11713 34632
rect 11747 34660 11759 34663
rect 12434 34660 12440 34672
rect 11747 34632 12440 34660
rect 11747 34629 11759 34632
rect 11701 34623 11759 34629
rect 12434 34620 12440 34632
rect 12492 34620 12498 34672
rect 15286 34620 15292 34672
rect 15344 34660 15350 34672
rect 16482 34660 16488 34672
rect 15344 34632 16488 34660
rect 15344 34620 15350 34632
rect 16482 34620 16488 34632
rect 16540 34660 16546 34672
rect 20717 34663 20775 34669
rect 16540 34632 16896 34660
rect 16540 34620 16546 34632
rect 7834 34592 7840 34604
rect 7795 34564 7840 34592
rect 7834 34552 7840 34564
rect 7892 34552 7898 34604
rect 8021 34595 8079 34601
rect 8021 34561 8033 34595
rect 8067 34592 8079 34595
rect 9490 34592 9496 34604
rect 8067 34564 9496 34592
rect 8067 34561 8079 34564
rect 8021 34555 8079 34561
rect 9490 34552 9496 34564
rect 9548 34592 9554 34604
rect 10597 34595 10655 34601
rect 10597 34592 10609 34595
rect 9548 34564 10609 34592
rect 9548 34552 9554 34564
rect 10597 34561 10609 34564
rect 10643 34592 10655 34595
rect 11514 34592 11520 34604
rect 10643 34564 11520 34592
rect 10643 34561 10655 34564
rect 10597 34555 10655 34561
rect 11514 34552 11520 34564
rect 11572 34552 11578 34604
rect 12342 34592 12348 34604
rect 12303 34564 12348 34592
rect 12342 34552 12348 34564
rect 12400 34552 12406 34604
rect 12526 34552 12532 34604
rect 12584 34592 12590 34604
rect 12713 34595 12771 34601
rect 12713 34592 12725 34595
rect 12584 34564 12725 34592
rect 12584 34552 12590 34564
rect 12713 34561 12725 34564
rect 12759 34561 12771 34595
rect 12713 34555 12771 34561
rect 15473 34595 15531 34601
rect 15473 34561 15485 34595
rect 15519 34592 15531 34595
rect 15838 34592 15844 34604
rect 15519 34564 15844 34592
rect 15519 34561 15531 34564
rect 15473 34555 15531 34561
rect 15838 34552 15844 34564
rect 15896 34592 15902 34604
rect 16868 34601 16896 34632
rect 20717 34629 20729 34663
rect 20763 34629 20775 34663
rect 20717 34623 20775 34629
rect 20933 34663 20991 34669
rect 20933 34629 20945 34663
rect 20979 34660 20991 34663
rect 22646 34660 22652 34672
rect 20979 34632 22652 34660
rect 20979 34629 20991 34632
rect 20933 34623 20991 34629
rect 16669 34595 16727 34601
rect 16669 34592 16681 34595
rect 15896 34564 16681 34592
rect 15896 34552 15902 34564
rect 16669 34561 16681 34564
rect 16715 34561 16727 34595
rect 16669 34555 16727 34561
rect 16853 34595 16911 34601
rect 16853 34561 16865 34595
rect 16899 34561 16911 34595
rect 16853 34555 16911 34561
rect 17402 34552 17408 34604
rect 17460 34592 17466 34604
rect 17862 34592 17868 34604
rect 17460 34564 17868 34592
rect 17460 34552 17466 34564
rect 17862 34552 17868 34564
rect 17920 34592 17926 34604
rect 18141 34595 18199 34601
rect 18141 34592 18153 34595
rect 17920 34564 18153 34592
rect 17920 34552 17926 34564
rect 18141 34561 18153 34564
rect 18187 34561 18199 34595
rect 18322 34592 18328 34604
rect 18283 34564 18328 34592
rect 18141 34555 18199 34561
rect 18322 34552 18328 34564
rect 18380 34552 18386 34604
rect 18414 34552 18420 34604
rect 18472 34592 18478 34604
rect 20073 34595 20131 34601
rect 18472 34564 18517 34592
rect 18472 34552 18478 34564
rect 20073 34561 20085 34595
rect 20119 34561 20131 34595
rect 20073 34555 20131 34561
rect 7006 34484 7012 34536
rect 7064 34524 7070 34536
rect 7193 34527 7251 34533
rect 7193 34524 7205 34527
rect 7064 34496 7205 34524
rect 7064 34484 7070 34496
rect 7193 34493 7205 34496
rect 7239 34524 7251 34527
rect 7926 34524 7932 34536
rect 7239 34496 7932 34524
rect 7239 34493 7251 34496
rect 7193 34487 7251 34493
rect 7926 34484 7932 34496
rect 7984 34524 7990 34536
rect 9033 34527 9091 34533
rect 9033 34524 9045 34527
rect 7984 34496 9045 34524
rect 7984 34484 7990 34496
rect 9033 34493 9045 34496
rect 9079 34493 9091 34527
rect 9033 34487 9091 34493
rect 10965 34527 11023 34533
rect 10965 34493 10977 34527
rect 11011 34524 11023 34527
rect 11606 34524 11612 34536
rect 11011 34496 11612 34524
rect 11011 34493 11023 34496
rect 10965 34487 11023 34493
rect 11606 34484 11612 34496
rect 11664 34484 11670 34536
rect 15194 34524 15200 34536
rect 15155 34496 15200 34524
rect 15194 34484 15200 34496
rect 15252 34484 15258 34536
rect 16114 34524 16120 34536
rect 16075 34496 16120 34524
rect 16114 34484 16120 34496
rect 16172 34484 16178 34536
rect 11146 34416 11152 34468
rect 11204 34456 11210 34468
rect 11517 34459 11575 34465
rect 11517 34456 11529 34459
rect 11204 34428 11529 34456
rect 11204 34416 11210 34428
rect 11517 34425 11529 34428
rect 11563 34425 11575 34459
rect 11517 34419 11575 34425
rect 18322 34416 18328 34468
rect 18380 34456 18386 34468
rect 20088 34456 20116 34555
rect 20162 34552 20168 34604
rect 20220 34592 20226 34604
rect 20257 34595 20315 34601
rect 20257 34592 20269 34595
rect 20220 34564 20269 34592
rect 20220 34552 20226 34564
rect 20257 34561 20269 34564
rect 20303 34592 20315 34595
rect 20732 34592 20760 34623
rect 22646 34620 22652 34632
rect 22704 34620 22710 34672
rect 24486 34620 24492 34672
rect 24544 34660 24550 34672
rect 25041 34663 25099 34669
rect 25041 34660 25053 34663
rect 24544 34632 25053 34660
rect 24544 34620 24550 34632
rect 25041 34629 25053 34632
rect 25087 34629 25099 34663
rect 27890 34660 27896 34672
rect 27851 34632 27896 34660
rect 25041 34623 25099 34629
rect 27890 34620 27896 34632
rect 27948 34620 27954 34672
rect 34790 34620 34796 34672
rect 34848 34660 34854 34672
rect 35161 34663 35219 34669
rect 35161 34660 35173 34663
rect 34848 34632 35173 34660
rect 34848 34620 34854 34632
rect 35161 34629 35173 34632
rect 35207 34629 35219 34663
rect 35161 34623 35219 34629
rect 35345 34663 35403 34669
rect 35345 34629 35357 34663
rect 35391 34660 35403 34663
rect 39117 34663 39175 34669
rect 35391 34632 39068 34660
rect 35391 34629 35403 34632
rect 35345 34623 35403 34629
rect 24946 34592 24952 34604
rect 20303 34564 20760 34592
rect 24907 34564 24952 34592
rect 20303 34561 20315 34564
rect 20257 34555 20315 34561
rect 24946 34552 24952 34564
rect 25004 34552 25010 34604
rect 25130 34552 25136 34604
rect 25188 34592 25194 34604
rect 25225 34595 25283 34601
rect 25225 34592 25237 34595
rect 25188 34564 25237 34592
rect 25188 34552 25194 34564
rect 25225 34561 25237 34564
rect 25271 34561 25283 34595
rect 25225 34555 25283 34561
rect 25409 34595 25467 34601
rect 25409 34561 25421 34595
rect 25455 34592 25467 34595
rect 27709 34595 27767 34601
rect 27709 34592 27721 34595
rect 25455 34564 27721 34592
rect 25455 34561 25467 34564
rect 25409 34555 25467 34561
rect 27709 34561 27721 34564
rect 27755 34592 27767 34595
rect 27798 34592 27804 34604
rect 27755 34564 27804 34592
rect 27755 34561 27767 34564
rect 27709 34555 27767 34561
rect 27798 34552 27804 34564
rect 27856 34552 27862 34604
rect 27985 34595 28043 34601
rect 27985 34561 27997 34595
rect 28031 34592 28043 34595
rect 28442 34592 28448 34604
rect 28031 34564 28448 34592
rect 28031 34561 28043 34564
rect 27985 34555 28043 34561
rect 27249 34527 27307 34533
rect 27249 34493 27261 34527
rect 27295 34524 27307 34527
rect 28000 34524 28028 34555
rect 28442 34552 28448 34564
rect 28500 34552 28506 34604
rect 32398 34592 32404 34604
rect 32359 34564 32404 34592
rect 32398 34552 32404 34564
rect 32456 34552 32462 34604
rect 32766 34592 32772 34604
rect 32727 34564 32772 34592
rect 32766 34552 32772 34564
rect 32824 34552 32830 34604
rect 34977 34595 35035 34601
rect 34977 34561 34989 34595
rect 35023 34561 35035 34595
rect 35176 34592 35204 34623
rect 35805 34595 35863 34601
rect 35805 34592 35817 34595
rect 35176 34564 35817 34592
rect 34977 34555 35035 34561
rect 35805 34561 35817 34564
rect 35851 34561 35863 34595
rect 35986 34592 35992 34604
rect 35947 34564 35992 34592
rect 35805 34555 35863 34561
rect 27295 34496 28028 34524
rect 34992 34524 35020 34555
rect 35986 34552 35992 34564
rect 36044 34552 36050 34604
rect 37826 34592 37832 34604
rect 37787 34564 37832 34592
rect 37826 34552 37832 34564
rect 37884 34552 37890 34604
rect 38194 34552 38200 34604
rect 38252 34592 38258 34604
rect 38657 34595 38715 34601
rect 38657 34592 38669 34595
rect 38252 34564 38669 34592
rect 38252 34552 38258 34564
rect 38657 34561 38669 34564
rect 38703 34561 38715 34595
rect 38930 34592 38936 34604
rect 38891 34564 38936 34592
rect 38657 34555 38715 34561
rect 38930 34552 38936 34564
rect 38988 34552 38994 34604
rect 39040 34592 39068 34632
rect 39117 34629 39129 34663
rect 39163 34660 39175 34663
rect 39163 34632 40264 34660
rect 39163 34629 39175 34632
rect 39117 34623 39175 34629
rect 40034 34592 40040 34604
rect 39040 34564 39896 34592
rect 39995 34564 40040 34592
rect 35342 34524 35348 34536
rect 34992 34496 35348 34524
rect 27295 34493 27307 34496
rect 27249 34487 27307 34493
rect 35342 34484 35348 34496
rect 35400 34484 35406 34536
rect 37458 34484 37464 34536
rect 37516 34524 37522 34536
rect 37921 34527 37979 34533
rect 37921 34524 37933 34527
rect 37516 34496 37933 34524
rect 37516 34484 37522 34496
rect 37921 34493 37933 34496
rect 37967 34524 37979 34527
rect 38286 34524 38292 34536
rect 37967 34496 38292 34524
rect 37967 34493 37979 34496
rect 37921 34487 37979 34493
rect 38286 34484 38292 34496
rect 38344 34524 38350 34536
rect 39669 34527 39727 34533
rect 39669 34524 39681 34527
rect 38344 34496 39681 34524
rect 38344 34484 38350 34496
rect 39669 34493 39681 34496
rect 39715 34493 39727 34527
rect 39868 34524 39896 34564
rect 40034 34552 40040 34564
rect 40092 34552 40098 34604
rect 40126 34524 40132 34536
rect 39868 34496 39988 34524
rect 40087 34496 40132 34524
rect 39669 34487 39727 34493
rect 27982 34456 27988 34468
rect 18380 34428 20944 34456
rect 27943 34428 27988 34456
rect 18380 34416 18386 34428
rect 7650 34388 7656 34400
rect 7611 34360 7656 34388
rect 7650 34348 7656 34360
rect 7708 34348 7714 34400
rect 14090 34348 14096 34400
rect 14148 34388 14154 34400
rect 20916 34397 20944 34428
rect 27982 34416 27988 34428
rect 28040 34416 28046 34468
rect 33594 34456 33600 34468
rect 33555 34428 33600 34456
rect 33594 34416 33600 34428
rect 33652 34416 33658 34468
rect 35894 34456 35900 34468
rect 35855 34428 35900 34456
rect 35894 34416 35900 34428
rect 35952 34416 35958 34468
rect 38378 34416 38384 34468
rect 38436 34456 38442 34468
rect 38749 34459 38807 34465
rect 38749 34456 38761 34459
rect 38436 34428 38761 34456
rect 38436 34416 38442 34428
rect 38749 34425 38761 34428
rect 38795 34425 38807 34459
rect 39960 34456 39988 34496
rect 40126 34484 40132 34496
rect 40184 34484 40190 34536
rect 40236 34524 40264 34632
rect 40310 34620 40316 34672
rect 40368 34660 40374 34672
rect 48682 34660 48688 34672
rect 40368 34632 48688 34660
rect 40368 34620 40374 34632
rect 48682 34620 48688 34632
rect 48740 34620 48746 34672
rect 48792 34632 50384 34660
rect 42886 34552 42892 34604
rect 42944 34592 42950 34604
rect 42981 34595 43039 34601
rect 42981 34592 42993 34595
rect 42944 34564 42993 34592
rect 42944 34552 42950 34564
rect 42981 34561 42993 34564
rect 43027 34561 43039 34595
rect 42981 34555 43039 34561
rect 43162 34552 43168 34604
rect 43220 34592 43226 34604
rect 43220 34564 43265 34592
rect 43220 34552 43226 34564
rect 48406 34552 48412 34604
rect 48464 34592 48470 34604
rect 48501 34595 48559 34601
rect 48501 34592 48513 34595
rect 48464 34564 48513 34592
rect 48464 34552 48470 34564
rect 48501 34561 48513 34564
rect 48547 34561 48559 34595
rect 48501 34555 48559 34561
rect 45094 34524 45100 34536
rect 40236 34496 45100 34524
rect 45094 34484 45100 34496
rect 45152 34484 45158 34536
rect 48792 34533 48820 34632
rect 49697 34595 49755 34601
rect 49697 34592 49709 34595
rect 48976 34564 49709 34592
rect 48777 34527 48835 34533
rect 48777 34493 48789 34527
rect 48823 34524 48835 34527
rect 48866 34524 48872 34536
rect 48823 34496 48872 34524
rect 48823 34493 48835 34496
rect 48777 34487 48835 34493
rect 48866 34484 48872 34496
rect 48924 34484 48930 34536
rect 40310 34456 40316 34468
rect 39960 34428 40316 34456
rect 38749 34419 38807 34425
rect 40310 34416 40316 34428
rect 40368 34416 40374 34468
rect 43165 34459 43223 34465
rect 43165 34425 43177 34459
rect 43211 34456 43223 34459
rect 43254 34456 43260 34468
rect 43211 34428 43260 34456
rect 43211 34425 43223 34428
rect 43165 34419 43223 34425
rect 43254 34416 43260 34428
rect 43312 34416 43318 34468
rect 48498 34416 48504 34468
rect 48556 34456 48562 34468
rect 48593 34459 48651 34465
rect 48593 34456 48605 34459
rect 48556 34428 48605 34456
rect 48556 34416 48562 34428
rect 48593 34425 48605 34428
rect 48639 34456 48651 34459
rect 48976 34456 49004 34564
rect 49697 34561 49709 34564
rect 49743 34561 49755 34595
rect 49970 34592 49976 34604
rect 49931 34564 49976 34592
rect 49697 34555 49755 34561
rect 49970 34552 49976 34564
rect 50028 34552 50034 34604
rect 50356 34601 50384 34632
rect 52454 34620 52460 34672
rect 52512 34660 52518 34672
rect 53009 34663 53067 34669
rect 53009 34660 53021 34663
rect 52512 34632 53021 34660
rect 52512 34620 52518 34632
rect 53009 34629 53021 34632
rect 53055 34660 53067 34663
rect 54113 34663 54171 34669
rect 54113 34660 54125 34663
rect 53055 34632 54125 34660
rect 53055 34629 53067 34632
rect 53009 34623 53067 34629
rect 54113 34629 54125 34632
rect 54159 34629 54171 34663
rect 54113 34623 54171 34629
rect 50341 34595 50399 34601
rect 50341 34561 50353 34595
rect 50387 34561 50399 34595
rect 50341 34555 50399 34561
rect 51997 34595 52055 34601
rect 51997 34561 52009 34595
rect 52043 34561 52055 34595
rect 51997 34555 52055 34561
rect 52181 34595 52239 34601
rect 52181 34561 52193 34595
rect 52227 34592 52239 34595
rect 52227 34564 52316 34592
rect 52227 34561 52239 34564
rect 52181 34555 52239 34561
rect 49421 34527 49479 34533
rect 49421 34493 49433 34527
rect 49467 34524 49479 34527
rect 49510 34524 49516 34536
rect 49467 34496 49516 34524
rect 49467 34493 49479 34496
rect 49421 34487 49479 34493
rect 49510 34484 49516 34496
rect 49568 34484 49574 34536
rect 48639 34428 49004 34456
rect 50709 34459 50767 34465
rect 48639 34425 48651 34428
rect 48593 34419 48651 34425
rect 50709 34425 50721 34459
rect 50755 34456 50767 34459
rect 52012 34456 52040 34555
rect 52178 34456 52184 34468
rect 50755 34428 52184 34456
rect 50755 34425 50767 34428
rect 50709 34419 50767 34425
rect 52178 34416 52184 34428
rect 52236 34416 52242 34468
rect 14185 34391 14243 34397
rect 14185 34388 14197 34391
rect 14148 34360 14197 34388
rect 14148 34348 14154 34360
rect 14185 34357 14197 34360
rect 14231 34357 14243 34391
rect 14185 34351 14243 34357
rect 20901 34391 20959 34397
rect 20901 34357 20913 34391
rect 20947 34357 20959 34391
rect 28442 34388 28448 34400
rect 28403 34360 28448 34388
rect 20901 34351 20959 34357
rect 28442 34348 28448 34360
rect 28500 34348 28506 34400
rect 38102 34388 38108 34400
rect 38063 34360 38108 34388
rect 38102 34348 38108 34360
rect 38160 34348 38166 34400
rect 49418 34348 49424 34400
rect 49476 34388 49482 34400
rect 52288 34388 52316 34564
rect 52638 34552 52644 34604
rect 52696 34592 52702 34604
rect 52733 34595 52791 34601
rect 52733 34592 52745 34595
rect 52696 34564 52745 34592
rect 52696 34552 52702 34564
rect 52733 34561 52745 34564
rect 52779 34561 52791 34595
rect 52733 34555 52791 34561
rect 52822 34552 52828 34604
rect 52880 34592 52886 34604
rect 53466 34592 53472 34604
rect 52880 34564 52925 34592
rect 53427 34564 53472 34592
rect 52880 34552 52886 34564
rect 53466 34552 53472 34564
rect 53524 34552 53530 34604
rect 53653 34595 53711 34601
rect 53653 34561 53665 34595
rect 53699 34561 53711 34595
rect 53653 34555 53711 34561
rect 53668 34524 53696 34555
rect 53024 34496 53696 34524
rect 53024 34465 53052 34496
rect 53009 34459 53067 34465
rect 53009 34425 53021 34459
rect 53055 34425 53067 34459
rect 53009 34419 53067 34425
rect 52914 34388 52920 34400
rect 49476 34360 52920 34388
rect 49476 34348 49482 34360
rect 52914 34348 52920 34360
rect 52972 34348 52978 34400
rect 1104 34298 58880 34320
rect 1104 34246 4214 34298
rect 4266 34246 4278 34298
rect 4330 34246 4342 34298
rect 4394 34246 4406 34298
rect 4458 34246 4470 34298
rect 4522 34246 34934 34298
rect 34986 34246 34998 34298
rect 35050 34246 35062 34298
rect 35114 34246 35126 34298
rect 35178 34246 35190 34298
rect 35242 34246 58880 34298
rect 1104 34224 58880 34246
rect 10873 34187 10931 34193
rect 10873 34153 10885 34187
rect 10919 34184 10931 34187
rect 11698 34184 11704 34196
rect 10919 34156 11704 34184
rect 10919 34153 10931 34156
rect 10873 34147 10931 34153
rect 11698 34144 11704 34156
rect 11756 34144 11762 34196
rect 15194 34184 15200 34196
rect 15155 34156 15200 34184
rect 15194 34144 15200 34156
rect 15252 34144 15258 34196
rect 16025 34187 16083 34193
rect 16025 34153 16037 34187
rect 16071 34184 16083 34187
rect 17402 34184 17408 34196
rect 16071 34156 17408 34184
rect 16071 34153 16083 34156
rect 16025 34147 16083 34153
rect 17402 34144 17408 34156
rect 17460 34144 17466 34196
rect 18414 34144 18420 34196
rect 18472 34184 18478 34196
rect 19245 34187 19303 34193
rect 19245 34184 19257 34187
rect 18472 34156 19257 34184
rect 18472 34144 18478 34156
rect 19245 34153 19257 34156
rect 19291 34153 19303 34187
rect 25130 34184 25136 34196
rect 25091 34156 25136 34184
rect 19245 34147 19303 34153
rect 25130 34144 25136 34156
rect 25188 34144 25194 34196
rect 27614 34144 27620 34196
rect 27672 34184 27678 34196
rect 27890 34184 27896 34196
rect 27672 34156 27896 34184
rect 27672 34144 27678 34156
rect 27890 34144 27896 34156
rect 27948 34144 27954 34196
rect 28534 34184 28540 34196
rect 28495 34156 28540 34184
rect 28534 34144 28540 34156
rect 28592 34144 28598 34196
rect 32766 34184 32772 34196
rect 32232 34156 32772 34184
rect 11790 34116 11796 34128
rect 11532 34088 11796 34116
rect 11532 34057 11560 34088
rect 11790 34076 11796 34088
rect 11848 34116 11854 34128
rect 12158 34116 12164 34128
rect 11848 34088 12164 34116
rect 11848 34076 11854 34088
rect 12158 34076 12164 34088
rect 12216 34076 12222 34128
rect 16114 34076 16120 34128
rect 16172 34116 16178 34128
rect 24946 34116 24952 34128
rect 16172 34088 24952 34116
rect 16172 34076 16178 34088
rect 24946 34076 24952 34088
rect 25004 34076 25010 34128
rect 28350 34076 28356 34128
rect 28408 34116 28414 34128
rect 28905 34119 28963 34125
rect 28905 34116 28917 34119
rect 28408 34088 28917 34116
rect 28408 34076 28414 34088
rect 28905 34085 28917 34088
rect 28951 34085 28963 34119
rect 28905 34079 28963 34085
rect 11517 34051 11575 34057
rect 11517 34017 11529 34051
rect 11563 34017 11575 34051
rect 11517 34011 11575 34017
rect 11701 34051 11759 34057
rect 11701 34017 11713 34051
rect 11747 34048 11759 34051
rect 11882 34048 11888 34060
rect 11747 34020 11888 34048
rect 11747 34017 11759 34020
rect 11701 34011 11759 34017
rect 11882 34008 11888 34020
rect 11940 34008 11946 34060
rect 12066 34008 12072 34060
rect 12124 34048 12130 34060
rect 22278 34048 22284 34060
rect 12124 34020 22284 34048
rect 12124 34008 12130 34020
rect 22278 34008 22284 34020
rect 22336 34008 22342 34060
rect 22646 34048 22652 34060
rect 22607 34020 22652 34048
rect 22646 34008 22652 34020
rect 22704 34008 22710 34060
rect 23382 34048 23388 34060
rect 23343 34020 23388 34048
rect 23382 34008 23388 34020
rect 23440 34008 23446 34060
rect 32232 34057 32260 34156
rect 32766 34144 32772 34156
rect 32824 34144 32830 34196
rect 33137 34187 33195 34193
rect 33137 34153 33149 34187
rect 33183 34184 33195 34187
rect 34790 34184 34796 34196
rect 33183 34156 34796 34184
rect 33183 34153 33195 34156
rect 33137 34147 33195 34153
rect 34790 34144 34796 34156
rect 34848 34144 34854 34196
rect 38378 34184 38384 34196
rect 38339 34156 38384 34184
rect 38378 34144 38384 34156
rect 38436 34144 38442 34196
rect 40037 34187 40095 34193
rect 40037 34153 40049 34187
rect 40083 34184 40095 34187
rect 40126 34184 40132 34196
rect 40083 34156 40132 34184
rect 40083 34153 40095 34156
rect 40037 34147 40095 34153
rect 40126 34144 40132 34156
rect 40184 34144 40190 34196
rect 43162 34144 43168 34196
rect 43220 34184 43226 34196
rect 43809 34187 43867 34193
rect 43809 34184 43821 34187
rect 43220 34156 43821 34184
rect 43220 34144 43226 34156
rect 43809 34153 43821 34156
rect 43855 34153 43867 34187
rect 48682 34184 48688 34196
rect 48643 34156 48688 34184
rect 43809 34147 43867 34153
rect 48682 34144 48688 34156
rect 48740 34144 48746 34196
rect 49418 34144 49424 34196
rect 49476 34184 49482 34196
rect 49513 34187 49571 34193
rect 49513 34184 49525 34187
rect 49476 34156 49525 34184
rect 49476 34144 49482 34156
rect 49513 34153 49525 34156
rect 49559 34153 49571 34187
rect 49513 34147 49571 34153
rect 38286 34116 38292 34128
rect 38247 34088 38292 34116
rect 38286 34076 38292 34088
rect 38344 34076 38350 34128
rect 40218 34076 40224 34128
rect 40276 34116 40282 34128
rect 42245 34119 42303 34125
rect 40276 34088 42196 34116
rect 40276 34076 40282 34088
rect 32217 34051 32275 34057
rect 32217 34017 32229 34051
rect 32263 34017 32275 34051
rect 35894 34048 35900 34060
rect 35855 34020 35900 34048
rect 32217 34011 32275 34017
rect 35894 34008 35900 34020
rect 35952 34008 35958 34060
rect 37277 34051 37335 34057
rect 37277 34017 37289 34051
rect 37323 34048 37335 34051
rect 37826 34048 37832 34060
rect 37323 34020 37832 34048
rect 37323 34017 37335 34020
rect 37277 34011 37335 34017
rect 37826 34008 37832 34020
rect 37884 34048 37890 34060
rect 37921 34051 37979 34057
rect 37921 34048 37933 34051
rect 37884 34020 37933 34048
rect 37884 34008 37890 34020
rect 37921 34017 37933 34020
rect 37967 34017 37979 34051
rect 37921 34011 37979 34017
rect 39960 34020 40816 34048
rect 35440 33992 35492 33998
rect 39960 33992 39988 34020
rect 7834 33940 7840 33992
rect 7892 33980 7898 33992
rect 8113 33983 8171 33989
rect 8113 33980 8125 33983
rect 7892 33952 8125 33980
rect 7892 33940 7898 33952
rect 8113 33949 8125 33952
rect 8159 33949 8171 33983
rect 8113 33943 8171 33949
rect 8128 33912 8156 33943
rect 8202 33940 8208 33992
rect 8260 33980 8266 33992
rect 8389 33983 8447 33989
rect 8389 33980 8401 33983
rect 8260 33952 8401 33980
rect 8260 33940 8266 33952
rect 8389 33949 8401 33952
rect 8435 33980 8447 33983
rect 9122 33980 9128 33992
rect 8435 33952 9128 33980
rect 8435 33949 8447 33952
rect 8389 33943 8447 33949
rect 9122 33940 9128 33952
rect 9180 33940 9186 33992
rect 9309 33983 9367 33989
rect 9309 33949 9321 33983
rect 9355 33980 9367 33983
rect 9766 33980 9772 33992
rect 9355 33952 9772 33980
rect 9355 33949 9367 33952
rect 9309 33943 9367 33949
rect 9766 33940 9772 33952
rect 9824 33980 9830 33992
rect 10873 33983 10931 33989
rect 10873 33980 10885 33983
rect 9824 33952 10885 33980
rect 9824 33940 9830 33952
rect 10873 33949 10885 33952
rect 10919 33949 10931 33983
rect 10873 33943 10931 33949
rect 11057 33983 11115 33989
rect 11057 33949 11069 33983
rect 11103 33980 11115 33983
rect 11146 33980 11152 33992
rect 11103 33952 11152 33980
rect 11103 33949 11115 33952
rect 11057 33943 11115 33949
rect 11146 33940 11152 33952
rect 11204 33940 11210 33992
rect 11606 33940 11612 33992
rect 11664 33980 11670 33992
rect 12437 33983 12495 33989
rect 12437 33980 12449 33983
rect 11664 33952 12449 33980
rect 11664 33940 11670 33952
rect 12437 33949 12449 33952
rect 12483 33949 12495 33983
rect 12437 33943 12495 33949
rect 12621 33983 12679 33989
rect 12621 33949 12633 33983
rect 12667 33949 12679 33983
rect 12894 33980 12900 33992
rect 12855 33952 12900 33980
rect 12621 33943 12679 33949
rect 8294 33912 8300 33924
rect 8128 33884 8300 33912
rect 8294 33872 8300 33884
rect 8352 33872 8358 33924
rect 9490 33912 9496 33924
rect 9451 33884 9496 33912
rect 9490 33872 9496 33884
rect 9548 33872 9554 33924
rect 12069 33915 12127 33921
rect 12069 33881 12081 33915
rect 12115 33881 12127 33915
rect 12636 33912 12664 33943
rect 12894 33940 12900 33952
rect 12952 33940 12958 33992
rect 14182 33940 14188 33992
rect 14240 33980 14246 33992
rect 15013 33983 15071 33989
rect 15013 33980 15025 33983
rect 14240 33952 15025 33980
rect 14240 33940 14246 33952
rect 15013 33949 15025 33952
rect 15059 33949 15071 33983
rect 15013 33943 15071 33949
rect 15197 33983 15255 33989
rect 15197 33949 15209 33983
rect 15243 33980 15255 33983
rect 15286 33980 15292 33992
rect 15243 33952 15292 33980
rect 15243 33949 15255 33952
rect 15197 33943 15255 33949
rect 12710 33912 12716 33924
rect 12623 33884 12716 33912
rect 12069 33875 12127 33881
rect 7282 33804 7288 33856
rect 7340 33844 7346 33856
rect 12084 33844 12112 33875
rect 12710 33872 12716 33884
rect 12768 33912 12774 33924
rect 13722 33912 13728 33924
rect 12768 33884 13728 33912
rect 12768 33872 12774 33884
rect 13722 33872 13728 33884
rect 13780 33872 13786 33924
rect 15028 33912 15056 33943
rect 15286 33940 15292 33952
rect 15344 33940 15350 33992
rect 15657 33983 15715 33989
rect 15657 33949 15669 33983
rect 15703 33949 15715 33983
rect 15838 33980 15844 33992
rect 15799 33952 15844 33980
rect 15657 33943 15715 33949
rect 15672 33912 15700 33943
rect 15838 33940 15844 33952
rect 15896 33940 15902 33992
rect 18414 33980 18420 33992
rect 18375 33952 18420 33980
rect 18414 33940 18420 33952
rect 18472 33980 18478 33992
rect 18693 33983 18751 33989
rect 18472 33952 18644 33980
rect 18472 33940 18478 33952
rect 18506 33912 18512 33924
rect 15028 33884 15700 33912
rect 18467 33884 18512 33912
rect 18506 33872 18512 33884
rect 18564 33872 18570 33924
rect 7340 33816 12112 33844
rect 7340 33804 7346 33816
rect 18322 33804 18328 33856
rect 18380 33844 18386 33856
rect 18417 33847 18475 33853
rect 18417 33844 18429 33847
rect 18380 33816 18429 33844
rect 18380 33804 18386 33816
rect 18417 33813 18429 33816
rect 18463 33813 18475 33847
rect 18616 33844 18644 33952
rect 18693 33949 18705 33983
rect 18739 33980 18751 33983
rect 19242 33980 19248 33992
rect 18739 33952 19248 33980
rect 18739 33949 18751 33952
rect 18693 33943 18751 33949
rect 19242 33940 19248 33952
rect 19300 33980 19306 33992
rect 19429 33983 19487 33989
rect 19429 33980 19441 33983
rect 19300 33952 19441 33980
rect 19300 33940 19306 33952
rect 19429 33949 19441 33952
rect 19475 33949 19487 33983
rect 19429 33943 19487 33949
rect 19705 33983 19763 33989
rect 19705 33949 19717 33983
rect 19751 33949 19763 33983
rect 19705 33943 19763 33949
rect 18782 33872 18788 33924
rect 18840 33912 18846 33924
rect 19720 33912 19748 33943
rect 23198 33940 23204 33992
rect 23256 33980 23262 33992
rect 23256 33952 23301 33980
rect 23256 33940 23262 33952
rect 28258 33940 28264 33992
rect 28316 33980 28322 33992
rect 28537 33983 28595 33989
rect 28537 33980 28549 33983
rect 28316 33952 28549 33980
rect 28316 33940 28322 33952
rect 28537 33949 28549 33952
rect 28583 33949 28595 33983
rect 28537 33943 28595 33949
rect 28629 33983 28687 33989
rect 28629 33949 28641 33983
rect 28675 33949 28687 33983
rect 28629 33943 28687 33949
rect 24670 33912 24676 33924
rect 18840 33884 19748 33912
rect 24631 33884 24676 33912
rect 18840 33872 18846 33884
rect 24670 33872 24676 33884
rect 24728 33872 24734 33924
rect 27706 33912 27712 33924
rect 27667 33884 27712 33912
rect 27706 33872 27712 33884
rect 27764 33872 27770 33924
rect 27798 33872 27804 33924
rect 27856 33912 27862 33924
rect 27909 33915 27967 33921
rect 27909 33912 27921 33915
rect 27856 33884 27921 33912
rect 27856 33872 27862 33884
rect 27909 33881 27921 33884
rect 27955 33881 27967 33915
rect 28644 33912 28672 33943
rect 31110 33940 31116 33992
rect 31168 33980 31174 33992
rect 31205 33983 31263 33989
rect 31205 33980 31217 33983
rect 31168 33952 31217 33980
rect 31168 33940 31174 33952
rect 31205 33949 31217 33952
rect 31251 33949 31263 33983
rect 31386 33980 31392 33992
rect 31347 33952 31392 33980
rect 31205 33943 31263 33949
rect 31386 33940 31392 33952
rect 31444 33940 31450 33992
rect 32398 33940 32404 33992
rect 32456 33980 32462 33992
rect 32677 33983 32735 33989
rect 32677 33980 32689 33983
rect 32456 33952 32689 33980
rect 32456 33940 32462 33952
rect 32677 33949 32689 33952
rect 32723 33949 32735 33983
rect 32677 33943 32735 33949
rect 37182 33980 37188 33992
rect 37143 33952 37188 33980
rect 37182 33940 37188 33952
rect 37240 33940 37246 33992
rect 37366 33980 37372 33992
rect 37327 33952 37372 33980
rect 37366 33940 37372 33952
rect 37424 33940 37430 33992
rect 39942 33980 39948 33992
rect 39903 33952 39948 33980
rect 39942 33940 39948 33952
rect 40000 33940 40006 33992
rect 40129 33983 40187 33989
rect 40129 33949 40141 33983
rect 40175 33980 40187 33983
rect 40310 33980 40316 33992
rect 40175 33952 40316 33980
rect 40175 33949 40187 33952
rect 40129 33943 40187 33949
rect 40310 33940 40316 33952
rect 40368 33940 40374 33992
rect 40788 33989 40816 34020
rect 40972 33989 41000 34088
rect 41782 34048 41788 34060
rect 41743 34020 41788 34048
rect 41782 34008 41788 34020
rect 41840 34008 41846 34060
rect 40773 33983 40831 33989
rect 40773 33949 40785 33983
rect 40819 33949 40831 33983
rect 40773 33943 40831 33949
rect 40957 33983 41015 33989
rect 40957 33949 40969 33983
rect 41003 33949 41015 33983
rect 40957 33943 41015 33949
rect 41877 33983 41935 33989
rect 41877 33949 41889 33983
rect 41923 33949 41935 33983
rect 42168 33980 42196 34088
rect 42245 34085 42257 34119
rect 42291 34085 42303 34119
rect 42245 34079 42303 34085
rect 42260 34048 42288 34079
rect 42886 34076 42892 34128
rect 42944 34116 42950 34128
rect 44177 34119 44235 34125
rect 42944 34088 43944 34116
rect 42944 34076 42950 34088
rect 43916 34057 43944 34088
rect 44177 34085 44189 34119
rect 44223 34085 44235 34119
rect 44177 34079 44235 34085
rect 43901 34051 43959 34057
rect 42260 34020 43208 34048
rect 42886 33980 42892 33992
rect 42168 33952 42892 33980
rect 41877 33943 41935 33949
rect 35440 33934 35492 33940
rect 35342 33912 35348 33924
rect 27909 33875 27967 33881
rect 28092 33884 28672 33912
rect 35255 33884 35348 33912
rect 28092 33856 28120 33884
rect 35342 33872 35348 33884
rect 35400 33872 35406 33924
rect 19613 33847 19671 33853
rect 19613 33844 19625 33847
rect 18616 33816 19625 33844
rect 18417 33807 18475 33813
rect 19613 33813 19625 33816
rect 19659 33844 19671 33847
rect 20162 33844 20168 33856
rect 19659 33816 20168 33844
rect 19659 33813 19671 33816
rect 19613 33807 19671 33813
rect 20162 33804 20168 33816
rect 20220 33804 20226 33856
rect 28074 33844 28080 33856
rect 28035 33816 28080 33844
rect 28074 33804 28080 33816
rect 28132 33804 28138 33856
rect 35360 33844 35388 33872
rect 37200 33844 37228 33940
rect 35360 33816 37228 33844
rect 40328 33844 40356 33940
rect 40865 33915 40923 33921
rect 40865 33881 40877 33915
rect 40911 33912 40923 33915
rect 41892 33912 41920 33943
rect 42886 33940 42892 33952
rect 42944 33940 42950 33992
rect 43180 33989 43208 34020
rect 43901 34017 43913 34051
rect 43947 34017 43959 34051
rect 43901 34011 43959 34017
rect 42981 33983 43039 33989
rect 42981 33949 42993 33983
rect 43027 33949 43039 33983
rect 42981 33943 43039 33949
rect 43165 33983 43223 33989
rect 43165 33949 43177 33983
rect 43211 33980 43223 33983
rect 43346 33980 43352 33992
rect 43211 33952 43352 33980
rect 43211 33949 43223 33952
rect 43165 33943 43223 33949
rect 42610 33912 42616 33924
rect 40911 33884 42616 33912
rect 40911 33881 40923 33884
rect 40865 33875 40923 33881
rect 42610 33872 42616 33884
rect 42668 33872 42674 33924
rect 42996 33844 43024 33943
rect 43346 33940 43352 33952
rect 43404 33980 43410 33992
rect 43809 33983 43867 33989
rect 43809 33980 43821 33983
rect 43404 33952 43821 33980
rect 43404 33940 43410 33952
rect 43809 33949 43821 33952
rect 43855 33949 43867 33983
rect 44192 33980 44220 34079
rect 46934 34076 46940 34128
rect 46992 34116 46998 34128
rect 50709 34119 50767 34125
rect 50709 34116 50721 34119
rect 46992 34088 50721 34116
rect 46992 34076 46998 34088
rect 50709 34085 50721 34088
rect 50755 34085 50767 34119
rect 50709 34079 50767 34085
rect 50724 34048 50752 34079
rect 52454 34048 52460 34060
rect 50724 34020 52460 34048
rect 45002 33980 45008 33992
rect 44192 33952 45008 33980
rect 43809 33943 43867 33949
rect 45002 33940 45008 33952
rect 45060 33940 45066 33992
rect 45094 33940 45100 33992
rect 45152 33980 45158 33992
rect 45281 33983 45339 33989
rect 45152 33952 45197 33980
rect 45152 33940 45158 33952
rect 45281 33949 45293 33983
rect 45327 33949 45339 33983
rect 45281 33943 45339 33949
rect 45296 33912 45324 33943
rect 48682 33940 48688 33992
rect 48740 33980 48746 33992
rect 49421 33983 49479 33989
rect 49421 33980 49433 33983
rect 48740 33952 49433 33980
rect 48740 33940 48746 33952
rect 49421 33949 49433 33952
rect 49467 33949 49479 33983
rect 51258 33980 51264 33992
rect 51219 33952 51264 33980
rect 49421 33943 49479 33949
rect 51258 33940 51264 33952
rect 51316 33940 51322 33992
rect 51552 33989 51580 34020
rect 52454 34008 52460 34020
rect 52512 34008 52518 34060
rect 53466 34048 53472 34060
rect 53427 34020 53472 34048
rect 53466 34008 53472 34020
rect 53524 34008 53530 34060
rect 51537 33983 51595 33989
rect 51537 33949 51549 33983
rect 51583 33949 51595 33983
rect 52178 33980 52184 33992
rect 52139 33952 52184 33980
rect 51537 33943 51595 33949
rect 52178 33940 52184 33952
rect 52236 33940 52242 33992
rect 52549 33983 52607 33989
rect 52549 33949 52561 33983
rect 52595 33949 52607 33983
rect 52914 33980 52920 33992
rect 52875 33952 52920 33980
rect 52549 33943 52607 33949
rect 43364 33884 45324 33912
rect 43364 33856 43392 33884
rect 49050 33872 49056 33924
rect 49108 33912 49114 33924
rect 49237 33915 49295 33921
rect 49237 33912 49249 33915
rect 49108 33884 49249 33912
rect 49108 33872 49114 33884
rect 49237 33881 49249 33884
rect 49283 33881 49295 33915
rect 49237 33875 49295 33881
rect 51721 33915 51779 33921
rect 51721 33881 51733 33915
rect 51767 33912 51779 33915
rect 52564 33912 52592 33943
rect 52914 33940 52920 33952
rect 52972 33940 52978 33992
rect 51767 33884 52592 33912
rect 53561 33915 53619 33921
rect 51767 33881 51779 33884
rect 51721 33875 51779 33881
rect 53561 33881 53573 33915
rect 53607 33912 53619 33915
rect 55582 33912 55588 33924
rect 53607 33884 55588 33912
rect 53607 33881 53619 33884
rect 53561 33875 53619 33881
rect 55582 33872 55588 33884
rect 55640 33872 55646 33924
rect 43162 33844 43168 33856
rect 40328 33816 43168 33844
rect 43162 33804 43168 33816
rect 43220 33804 43226 33856
rect 43346 33844 43352 33856
rect 43307 33816 43352 33844
rect 43346 33804 43352 33816
rect 43404 33804 43410 33856
rect 45465 33847 45523 33853
rect 45465 33813 45477 33847
rect 45511 33844 45523 33847
rect 45830 33844 45836 33856
rect 45511 33816 45836 33844
rect 45511 33813 45523 33816
rect 45465 33807 45523 33813
rect 45830 33804 45836 33816
rect 45888 33804 45894 33856
rect 51353 33847 51411 33853
rect 51353 33813 51365 33847
rect 51399 33844 51411 33847
rect 52178 33844 52184 33856
rect 51399 33816 52184 33844
rect 51399 33813 51411 33816
rect 51353 33807 51411 33813
rect 52178 33804 52184 33816
rect 52236 33804 52242 33856
rect 1104 33754 58880 33776
rect 1104 33702 19574 33754
rect 19626 33702 19638 33754
rect 19690 33702 19702 33754
rect 19754 33702 19766 33754
rect 19818 33702 19830 33754
rect 19882 33702 50294 33754
rect 50346 33702 50358 33754
rect 50410 33702 50422 33754
rect 50474 33702 50486 33754
rect 50538 33702 50550 33754
rect 50602 33702 58880 33754
rect 1104 33680 58880 33702
rect 11790 33640 11796 33652
rect 11751 33612 11796 33640
rect 11790 33600 11796 33612
rect 11848 33600 11854 33652
rect 17770 33640 17776 33652
rect 17144 33612 17776 33640
rect 17144 33584 17172 33612
rect 17770 33600 17776 33612
rect 17828 33640 17834 33652
rect 17957 33643 18015 33649
rect 17957 33640 17969 33643
rect 17828 33612 17969 33640
rect 17828 33600 17834 33612
rect 17957 33609 17969 33612
rect 18003 33609 18015 33643
rect 27614 33640 27620 33652
rect 27575 33612 27620 33640
rect 17957 33603 18015 33609
rect 27614 33600 27620 33612
rect 27672 33600 27678 33652
rect 27798 33600 27804 33652
rect 27856 33600 27862 33652
rect 31021 33643 31079 33649
rect 31021 33609 31033 33643
rect 31067 33640 31079 33643
rect 31386 33640 31392 33652
rect 31067 33612 31392 33640
rect 31067 33609 31079 33612
rect 31021 33603 31079 33609
rect 31386 33600 31392 33612
rect 31444 33600 31450 33652
rect 35710 33600 35716 33652
rect 35768 33640 35774 33652
rect 57977 33643 58035 33649
rect 57977 33640 57989 33643
rect 35768 33612 57989 33640
rect 35768 33600 35774 33612
rect 57977 33609 57989 33612
rect 58023 33609 58035 33643
rect 57977 33603 58035 33609
rect 8481 33575 8539 33581
rect 8481 33572 8493 33575
rect 6748 33544 8493 33572
rect 1578 33464 1584 33516
rect 1636 33504 1642 33516
rect 6748 33513 6776 33544
rect 8481 33541 8493 33544
rect 8527 33541 8539 33575
rect 9122 33572 9128 33584
rect 9035 33544 9128 33572
rect 8481 33535 8539 33541
rect 9122 33532 9128 33544
rect 9180 33572 9186 33584
rect 9677 33575 9735 33581
rect 9677 33572 9689 33575
rect 9180 33544 9689 33572
rect 9180 33532 9186 33544
rect 9677 33541 9689 33544
rect 9723 33572 9735 33575
rect 12066 33572 12072 33584
rect 9723 33544 12072 33572
rect 9723 33541 9735 33544
rect 9677 33535 9735 33541
rect 12066 33532 12072 33544
rect 12124 33532 12130 33584
rect 17126 33572 17132 33584
rect 17039 33544 17132 33572
rect 17126 33532 17132 33544
rect 17184 33532 17190 33584
rect 23293 33575 23351 33581
rect 23293 33541 23305 33575
rect 23339 33572 23351 33575
rect 23382 33572 23388 33584
rect 23339 33544 23388 33572
rect 23339 33541 23351 33544
rect 23293 33535 23351 33541
rect 23382 33532 23388 33544
rect 23440 33572 23446 33584
rect 25314 33572 25320 33584
rect 23440 33544 25320 33572
rect 23440 33532 23446 33544
rect 25314 33532 25320 33544
rect 25372 33532 25378 33584
rect 27816 33572 27844 33600
rect 28442 33572 28448 33584
rect 27540 33544 27844 33572
rect 27908 33544 28448 33572
rect 1857 33507 1915 33513
rect 1857 33504 1869 33507
rect 1636 33476 1869 33504
rect 1636 33464 1642 33476
rect 1857 33473 1869 33476
rect 1903 33473 1915 33507
rect 1857 33467 1915 33473
rect 6733 33507 6791 33513
rect 6733 33473 6745 33507
rect 6779 33473 6791 33507
rect 6733 33467 6791 33473
rect 6917 33507 6975 33513
rect 6917 33473 6929 33507
rect 6963 33504 6975 33507
rect 7561 33507 7619 33513
rect 6963 33476 7420 33504
rect 6963 33473 6975 33476
rect 6917 33467 6975 33473
rect 6641 33371 6699 33377
rect 6641 33337 6653 33371
rect 6687 33368 6699 33371
rect 7098 33368 7104 33380
rect 6687 33340 7104 33368
rect 6687 33337 6699 33340
rect 6641 33331 6699 33337
rect 7098 33328 7104 33340
rect 7156 33328 7162 33380
rect 7392 33368 7420 33476
rect 7561 33473 7573 33507
rect 7607 33504 7619 33507
rect 8202 33504 8208 33516
rect 7607 33476 8208 33504
rect 7607 33473 7619 33476
rect 7561 33467 7619 33473
rect 8202 33464 8208 33476
rect 8260 33464 8266 33516
rect 8294 33464 8300 33516
rect 8352 33504 8358 33516
rect 8389 33507 8447 33513
rect 8389 33504 8401 33507
rect 8352 33476 8401 33504
rect 8352 33464 8358 33476
rect 8389 33473 8401 33476
rect 8435 33473 8447 33507
rect 8389 33467 8447 33473
rect 8573 33507 8631 33513
rect 8573 33473 8585 33507
rect 8619 33504 8631 33507
rect 9766 33504 9772 33516
rect 8619 33476 9772 33504
rect 8619 33473 8631 33476
rect 8573 33467 8631 33473
rect 9766 33464 9772 33476
rect 9824 33464 9830 33516
rect 11606 33464 11612 33516
rect 11664 33504 11670 33516
rect 11977 33507 12035 33513
rect 11977 33504 11989 33507
rect 11664 33476 11989 33504
rect 11664 33464 11670 33476
rect 11977 33473 11989 33476
rect 12023 33473 12035 33507
rect 11977 33467 12035 33473
rect 22462 33464 22468 33516
rect 22520 33504 22526 33516
rect 23017 33507 23075 33513
rect 23017 33504 23029 33507
rect 22520 33476 23029 33504
rect 22520 33464 22526 33476
rect 23017 33473 23029 33476
rect 23063 33473 23075 33507
rect 23198 33504 23204 33516
rect 23159 33476 23204 33504
rect 23017 33467 23075 33473
rect 23198 33464 23204 33476
rect 23256 33464 23262 33516
rect 24670 33464 24676 33516
rect 24728 33504 24734 33516
rect 27540 33513 27568 33544
rect 24857 33507 24915 33513
rect 24857 33504 24869 33507
rect 24728 33476 24869 33504
rect 24728 33464 24734 33476
rect 24857 33473 24869 33476
rect 24903 33473 24915 33507
rect 24857 33467 24915 33473
rect 27525 33507 27583 33513
rect 27525 33473 27537 33507
rect 27571 33473 27583 33507
rect 27525 33467 27583 33473
rect 27706 33464 27712 33516
rect 27764 33504 27770 33516
rect 27801 33507 27859 33513
rect 27801 33504 27813 33507
rect 27764 33476 27813 33504
rect 27764 33464 27770 33476
rect 27801 33473 27813 33476
rect 27847 33504 27859 33507
rect 27908 33504 27936 33544
rect 28442 33532 28448 33544
rect 28500 33572 28506 33584
rect 28902 33572 28908 33584
rect 28500 33544 28908 33572
rect 28500 33532 28506 33544
rect 28902 33532 28908 33544
rect 28960 33532 28966 33584
rect 29089 33575 29147 33581
rect 29089 33541 29101 33575
rect 29135 33572 29147 33575
rect 42521 33575 42579 33581
rect 29135 33544 41414 33572
rect 29135 33541 29147 33544
rect 29089 33535 29147 33541
rect 28626 33504 28632 33516
rect 27847 33476 27936 33504
rect 28587 33476 28632 33504
rect 27847 33473 27859 33476
rect 27801 33467 27859 33473
rect 28626 33464 28632 33476
rect 28684 33464 28690 33516
rect 30929 33507 30987 33513
rect 30929 33473 30941 33507
rect 30975 33473 30987 33507
rect 31202 33504 31208 33516
rect 31163 33476 31208 33504
rect 30929 33467 30987 33473
rect 7469 33439 7527 33445
rect 7469 33405 7481 33439
rect 7515 33436 7527 33439
rect 8938 33436 8944 33448
rect 7515 33408 8944 33436
rect 7515 33405 7527 33408
rect 7469 33399 7527 33405
rect 8938 33396 8944 33408
rect 8996 33396 9002 33448
rect 12158 33436 12164 33448
rect 12071 33408 12164 33436
rect 12158 33396 12164 33408
rect 12216 33436 12222 33448
rect 17405 33439 17463 33445
rect 17405 33436 17417 33439
rect 12216 33408 17417 33436
rect 12216 33396 12222 33408
rect 17405 33405 17417 33408
rect 17451 33405 17463 33439
rect 24946 33436 24952 33448
rect 24907 33408 24952 33436
rect 17405 33399 17463 33405
rect 24946 33396 24952 33408
rect 25004 33396 25010 33448
rect 27065 33439 27123 33445
rect 27065 33405 27077 33439
rect 27111 33436 27123 33439
rect 27724 33436 27752 33464
rect 27111 33408 27752 33436
rect 27111 33405 27123 33408
rect 27065 33399 27123 33405
rect 28350 33396 28356 33448
rect 28408 33436 28414 33448
rect 28537 33439 28595 33445
rect 28537 33436 28549 33439
rect 28408 33408 28549 33436
rect 28408 33396 28414 33408
rect 28537 33405 28549 33408
rect 28583 33405 28595 33439
rect 30944 33436 30972 33467
rect 31202 33464 31208 33476
rect 31260 33464 31266 33516
rect 31389 33507 31447 33513
rect 31389 33473 31401 33507
rect 31435 33504 31447 33507
rect 35434 33504 35440 33516
rect 31435 33476 35440 33504
rect 31435 33473 31447 33476
rect 31389 33467 31447 33473
rect 35434 33464 35440 33476
rect 35492 33504 35498 33516
rect 35713 33507 35771 33513
rect 35713 33504 35725 33507
rect 35492 33476 35725 33504
rect 35492 33464 35498 33476
rect 35713 33473 35725 33476
rect 35759 33473 35771 33507
rect 35713 33467 35771 33473
rect 31110 33436 31116 33448
rect 30944 33408 31116 33436
rect 28537 33399 28595 33405
rect 31110 33396 31116 33408
rect 31168 33396 31174 33448
rect 36173 33439 36231 33445
rect 36173 33405 36185 33439
rect 36219 33436 36231 33439
rect 39942 33436 39948 33448
rect 36219 33408 39948 33436
rect 36219 33405 36231 33408
rect 36173 33399 36231 33405
rect 39942 33396 39948 33408
rect 40000 33396 40006 33448
rect 41386 33436 41414 33544
rect 42521 33541 42533 33575
rect 42567 33572 42579 33575
rect 48409 33575 48467 33581
rect 42567 33544 44956 33572
rect 42567 33541 42579 33544
rect 42521 33535 42579 33541
rect 44928 33516 44956 33544
rect 48409 33541 48421 33575
rect 48455 33572 48467 33575
rect 48498 33572 48504 33584
rect 48455 33544 48504 33572
rect 48455 33541 48467 33544
rect 48409 33535 48467 33541
rect 48498 33532 48504 33544
rect 48556 33532 48562 33584
rect 52181 33575 52239 33581
rect 52181 33541 52193 33575
rect 52227 33572 52239 33575
rect 52454 33572 52460 33584
rect 52227 33544 52460 33572
rect 52227 33541 52239 33544
rect 52181 33535 52239 33541
rect 52454 33532 52460 33544
rect 52512 33572 52518 33584
rect 52733 33575 52791 33581
rect 52733 33572 52745 33575
rect 52512 33544 52745 33572
rect 52512 33532 52518 33544
rect 52733 33541 52745 33544
rect 52779 33541 52791 33575
rect 52933 33575 52991 33581
rect 52933 33572 52945 33575
rect 52733 33535 52791 33541
rect 52840 33544 52945 33572
rect 41782 33464 41788 33516
rect 41840 33504 41846 33516
rect 42429 33507 42487 33513
rect 42429 33504 42441 33507
rect 41840 33476 42441 33504
rect 41840 33464 41846 33476
rect 42429 33473 42441 33476
rect 42475 33473 42487 33507
rect 42610 33504 42616 33516
rect 42571 33476 42616 33504
rect 42429 33467 42487 33473
rect 42610 33464 42616 33476
rect 42668 33464 42674 33516
rect 43346 33464 43352 33516
rect 43404 33504 43410 33516
rect 44637 33507 44695 33513
rect 44637 33504 44649 33507
rect 43404 33476 44649 33504
rect 43404 33464 43410 33476
rect 44637 33473 44649 33476
rect 44683 33473 44695 33507
rect 44637 33467 44695 33473
rect 44726 33464 44732 33516
rect 44784 33464 44790 33516
rect 44910 33504 44916 33516
rect 44823 33476 44916 33504
rect 44910 33464 44916 33476
rect 44968 33464 44974 33516
rect 45094 33504 45100 33516
rect 45055 33476 45100 33504
rect 45094 33464 45100 33476
rect 45152 33464 45158 33516
rect 45186 33464 45192 33516
rect 45244 33504 45250 33516
rect 45465 33507 45523 33513
rect 45465 33504 45477 33507
rect 45244 33476 45477 33504
rect 45244 33464 45250 33476
rect 45465 33473 45477 33476
rect 45511 33473 45523 33507
rect 48958 33504 48964 33516
rect 48919 33476 48964 33504
rect 45465 33467 45523 33473
rect 48958 33464 48964 33476
rect 49016 33464 49022 33516
rect 49326 33504 49332 33516
rect 49068 33476 49332 33504
rect 44744 33436 44772 33464
rect 41386 33408 44772 33436
rect 45002 33396 45008 33448
rect 45060 33436 45066 33448
rect 45373 33439 45431 33445
rect 45373 33436 45385 33439
rect 45060 33408 45385 33436
rect 45060 33396 45066 33408
rect 45373 33405 45385 33408
rect 45419 33405 45431 33439
rect 45373 33399 45431 33405
rect 47949 33439 48007 33445
rect 47949 33405 47961 33439
rect 47995 33436 48007 33439
rect 49068 33436 49096 33476
rect 49326 33464 49332 33476
rect 49384 33464 49390 33516
rect 51258 33464 51264 33516
rect 51316 33504 51322 33516
rect 52638 33504 52644 33516
rect 51316 33476 52644 33504
rect 51316 33464 51322 33476
rect 52638 33464 52644 33476
rect 52696 33504 52702 33516
rect 52840 33504 52868 33544
rect 52933 33541 52945 33544
rect 52979 33541 52991 33575
rect 52933 33535 52991 33541
rect 58158 33504 58164 33516
rect 52696 33476 52868 33504
rect 58119 33476 58164 33504
rect 52696 33464 52702 33476
rect 58158 33464 58164 33476
rect 58216 33464 58222 33516
rect 47995 33408 49096 33436
rect 47995 33405 48007 33408
rect 47949 33399 48007 33405
rect 7650 33368 7656 33380
rect 7392 33340 7656 33368
rect 7650 33328 7656 33340
rect 7708 33328 7714 33380
rect 7929 33371 7987 33377
rect 7929 33337 7941 33371
rect 7975 33368 7987 33371
rect 8110 33368 8116 33380
rect 7975 33340 8116 33368
rect 7975 33337 7987 33340
rect 7929 33331 7987 33337
rect 8110 33328 8116 33340
rect 8168 33328 8174 33380
rect 25225 33371 25283 33377
rect 25225 33337 25237 33371
rect 25271 33368 25283 33371
rect 26326 33368 26332 33380
rect 25271 33340 26332 33368
rect 25271 33337 25283 33340
rect 25225 33331 25283 33337
rect 26326 33328 26332 33340
rect 26384 33328 26390 33380
rect 32398 33368 32404 33380
rect 26896 33340 32404 33368
rect 1762 33260 1768 33312
rect 1820 33300 1826 33312
rect 1949 33303 2007 33309
rect 1949 33300 1961 33303
rect 1820 33272 1961 33300
rect 1820 33260 1826 33272
rect 1949 33269 1961 33272
rect 1995 33269 2007 33303
rect 1949 33263 2007 33269
rect 22833 33303 22891 33309
rect 22833 33269 22845 33303
rect 22879 33300 22891 33303
rect 26896 33300 26924 33340
rect 32398 33328 32404 33340
rect 32456 33328 32462 33380
rect 44729 33371 44787 33377
rect 44729 33337 44741 33371
rect 44775 33368 44787 33371
rect 45554 33368 45560 33380
rect 44775 33340 45560 33368
rect 44775 33337 44787 33340
rect 44729 33331 44787 33337
rect 45554 33328 45560 33340
rect 45612 33328 45618 33380
rect 53101 33371 53159 33377
rect 53101 33337 53113 33371
rect 53147 33368 53159 33371
rect 53466 33368 53472 33380
rect 53147 33340 53472 33368
rect 53147 33337 53159 33340
rect 53101 33331 53159 33337
rect 53466 33328 53472 33340
rect 53524 33328 53530 33380
rect 22879 33272 26924 33300
rect 27801 33303 27859 33309
rect 22879 33269 22891 33272
rect 22833 33263 22891 33269
rect 27801 33269 27813 33303
rect 27847 33300 27859 33303
rect 27982 33300 27988 33312
rect 27847 33272 27988 33300
rect 27847 33269 27859 33272
rect 27801 33263 27859 33269
rect 27982 33260 27988 33272
rect 28040 33300 28046 33312
rect 28534 33300 28540 33312
rect 28040 33272 28540 33300
rect 28040 33260 28046 33272
rect 28534 33260 28540 33272
rect 28592 33260 28598 33312
rect 30190 33260 30196 33312
rect 30248 33300 30254 33312
rect 35710 33300 35716 33312
rect 30248 33272 35716 33300
rect 30248 33260 30254 33272
rect 35710 33260 35716 33272
rect 35768 33260 35774 33312
rect 35894 33300 35900 33312
rect 35855 33272 35900 33300
rect 35894 33260 35900 33272
rect 35952 33260 35958 33312
rect 52178 33260 52184 33312
rect 52236 33300 52242 33312
rect 52822 33300 52828 33312
rect 52236 33272 52828 33300
rect 52236 33260 52242 33272
rect 52822 33260 52828 33272
rect 52880 33300 52886 33312
rect 52917 33303 52975 33309
rect 52917 33300 52929 33303
rect 52880 33272 52929 33300
rect 52880 33260 52886 33272
rect 52917 33269 52929 33272
rect 52963 33269 52975 33303
rect 52917 33263 52975 33269
rect 1104 33210 58880 33232
rect 1104 33158 4214 33210
rect 4266 33158 4278 33210
rect 4330 33158 4342 33210
rect 4394 33158 4406 33210
rect 4458 33158 4470 33210
rect 4522 33158 34934 33210
rect 34986 33158 34998 33210
rect 35050 33158 35062 33210
rect 35114 33158 35126 33210
rect 35178 33158 35190 33210
rect 35242 33158 58880 33210
rect 1104 33136 58880 33158
rect 1578 33096 1584 33108
rect 1539 33068 1584 33096
rect 1578 33056 1584 33068
rect 1636 33056 1642 33108
rect 8938 33096 8944 33108
rect 8899 33068 8944 33096
rect 8938 33056 8944 33068
rect 8996 33056 9002 33108
rect 18414 33056 18420 33108
rect 18472 33096 18478 33108
rect 18509 33099 18567 33105
rect 18509 33096 18521 33099
rect 18472 33068 18521 33096
rect 18472 33056 18478 33068
rect 18509 33065 18521 33068
rect 18555 33065 18567 33099
rect 18509 33059 18567 33065
rect 27982 33056 27988 33108
rect 28040 33096 28046 33108
rect 28077 33099 28135 33105
rect 28077 33096 28089 33099
rect 28040 33068 28089 33096
rect 28040 33056 28046 33068
rect 28077 33065 28089 33068
rect 28123 33065 28135 33099
rect 28077 33059 28135 33065
rect 28169 33099 28227 33105
rect 28169 33065 28181 33099
rect 28215 33096 28227 33099
rect 28626 33096 28632 33108
rect 28215 33068 28632 33096
rect 28215 33065 28227 33068
rect 28169 33059 28227 33065
rect 28626 33056 28632 33068
rect 28684 33056 28690 33108
rect 48866 33096 48872 33108
rect 48827 33068 48872 33096
rect 48866 33056 48872 33068
rect 48924 33056 48930 33108
rect 58158 33096 58164 33108
rect 58119 33068 58164 33096
rect 58158 33056 58164 33068
rect 58216 33056 58222 33108
rect 16669 33031 16727 33037
rect 16669 32997 16681 33031
rect 16715 33028 16727 33031
rect 17126 33028 17132 33040
rect 16715 33000 17132 33028
rect 16715 32997 16727 33000
rect 16669 32991 16727 32997
rect 17126 32988 17132 33000
rect 17184 32988 17190 33040
rect 19242 33028 19248 33040
rect 19203 33000 19248 33028
rect 19242 32988 19248 33000
rect 19300 32988 19306 33040
rect 27525 33031 27583 33037
rect 27525 32997 27537 33031
rect 27571 32997 27583 33031
rect 27525 32991 27583 32997
rect 7650 32960 7656 32972
rect 7611 32932 7656 32960
rect 7650 32920 7656 32932
rect 7708 32920 7714 32972
rect 18782 32920 18788 32972
rect 18840 32960 18846 32972
rect 19521 32963 19579 32969
rect 19521 32960 19533 32963
rect 18840 32932 19533 32960
rect 18840 32920 18846 32932
rect 19521 32929 19533 32932
rect 19567 32929 19579 32963
rect 19521 32923 19579 32929
rect 22833 32963 22891 32969
rect 22833 32929 22845 32963
rect 22879 32960 22891 32963
rect 23198 32960 23204 32972
rect 22879 32932 23204 32960
rect 22879 32929 22891 32932
rect 22833 32923 22891 32929
rect 23198 32920 23204 32932
rect 23256 32920 23262 32972
rect 26326 32960 26332 32972
rect 26287 32932 26332 32960
rect 26326 32920 26332 32932
rect 26384 32960 26390 32972
rect 27540 32960 27568 32991
rect 38654 32988 38660 33040
rect 38712 33028 38718 33040
rect 38749 33031 38807 33037
rect 38749 33028 38761 33031
rect 38712 33000 38761 33028
rect 38712 32988 38718 33000
rect 38749 32997 38761 33000
rect 38795 32997 38807 33031
rect 38749 32991 38807 32997
rect 28258 32960 28264 32972
rect 26384 32932 27292 32960
rect 27540 32932 28264 32960
rect 26384 32920 26390 32932
rect 7098 32892 7104 32904
rect 7059 32864 7104 32892
rect 7098 32852 7104 32864
rect 7156 32852 7162 32904
rect 7282 32892 7288 32904
rect 7243 32864 7288 32892
rect 7282 32852 7288 32864
rect 7340 32852 7346 32904
rect 8110 32892 8116 32904
rect 8071 32864 8116 32892
rect 8110 32852 8116 32864
rect 8168 32852 8174 32904
rect 11146 32852 11152 32904
rect 11204 32892 11210 32904
rect 11606 32892 11612 32904
rect 11204 32864 11612 32892
rect 11204 32852 11210 32864
rect 11606 32852 11612 32864
rect 11664 32852 11670 32904
rect 11974 32892 11980 32904
rect 11887 32864 11980 32892
rect 11974 32852 11980 32864
rect 12032 32892 12038 32904
rect 12158 32892 12164 32904
rect 12032 32864 12164 32892
rect 12032 32852 12038 32864
rect 12158 32852 12164 32864
rect 12216 32852 12222 32904
rect 16485 32895 16543 32901
rect 16485 32861 16497 32895
rect 16531 32892 16543 32895
rect 16574 32892 16580 32904
rect 16531 32864 16580 32892
rect 16531 32861 16543 32864
rect 16485 32855 16543 32861
rect 16574 32852 16580 32864
rect 16632 32852 16638 32904
rect 16761 32895 16819 32901
rect 16761 32861 16773 32895
rect 16807 32892 16819 32895
rect 16807 32864 17356 32892
rect 16807 32861 16819 32864
rect 16761 32855 16819 32861
rect 10870 32784 10876 32836
rect 10928 32824 10934 32836
rect 17218 32824 17224 32836
rect 10928 32796 17224 32824
rect 10928 32784 10934 32796
rect 17218 32784 17224 32796
rect 17276 32784 17282 32836
rect 7285 32759 7343 32765
rect 7285 32725 7297 32759
rect 7331 32756 7343 32759
rect 7374 32756 7380 32768
rect 7331 32728 7380 32756
rect 7331 32725 7343 32728
rect 7285 32719 7343 32725
rect 7374 32716 7380 32728
rect 7432 32716 7438 32768
rect 8110 32716 8116 32768
rect 8168 32756 8174 32768
rect 8297 32759 8355 32765
rect 8297 32756 8309 32759
rect 8168 32728 8309 32756
rect 8168 32716 8174 32728
rect 8297 32725 8309 32728
rect 8343 32725 8355 32759
rect 8297 32719 8355 32725
rect 12621 32759 12679 32765
rect 12621 32725 12633 32759
rect 12667 32756 12679 32759
rect 13262 32756 13268 32768
rect 12667 32728 13268 32756
rect 12667 32725 12679 32728
rect 12621 32719 12679 32725
rect 13262 32716 13268 32728
rect 13320 32716 13326 32768
rect 13722 32716 13728 32768
rect 13780 32756 13786 32768
rect 17328 32765 17356 32864
rect 18322 32852 18328 32904
rect 18380 32892 18386 32904
rect 18417 32895 18475 32901
rect 18417 32892 18429 32895
rect 18380 32864 18429 32892
rect 18380 32852 18386 32864
rect 18417 32861 18429 32864
rect 18463 32861 18475 32895
rect 18417 32855 18475 32861
rect 18506 32852 18512 32904
rect 18564 32892 18570 32904
rect 18564 32864 18609 32892
rect 18564 32852 18570 32864
rect 19334 32852 19340 32904
rect 19392 32892 19398 32904
rect 19613 32895 19671 32901
rect 19613 32892 19625 32895
rect 19392 32864 19625 32892
rect 19392 32852 19398 32864
rect 19613 32861 19625 32864
rect 19659 32892 19671 32895
rect 22002 32892 22008 32904
rect 19659 32864 20392 32892
rect 21963 32864 22008 32892
rect 19659 32861 19671 32864
rect 19613 32855 19671 32861
rect 18230 32824 18236 32836
rect 18191 32796 18236 32824
rect 18230 32784 18236 32796
rect 18288 32784 18294 32836
rect 16301 32759 16359 32765
rect 16301 32756 16313 32759
rect 13780 32728 16313 32756
rect 13780 32716 13786 32728
rect 16301 32725 16313 32728
rect 16347 32725 16359 32759
rect 16301 32719 16359 32725
rect 17313 32759 17371 32765
rect 17313 32725 17325 32759
rect 17359 32756 17371 32759
rect 17586 32756 17592 32768
rect 17359 32728 17592 32756
rect 17359 32725 17371 32728
rect 17313 32719 17371 32725
rect 17586 32716 17592 32728
rect 17644 32716 17650 32768
rect 20364 32765 20392 32864
rect 22002 32852 22008 32864
rect 22060 32852 22066 32904
rect 22278 32892 22284 32904
rect 22239 32864 22284 32892
rect 22278 32852 22284 32864
rect 22336 32852 22342 32904
rect 27264 32901 27292 32932
rect 28258 32920 28264 32932
rect 28316 32920 28322 32972
rect 30466 32960 30472 32972
rect 30427 32932 30472 32960
rect 30466 32920 30472 32932
rect 30524 32920 30530 32972
rect 31297 32963 31355 32969
rect 31297 32929 31309 32963
rect 31343 32960 31355 32963
rect 31386 32960 31392 32972
rect 31343 32932 31392 32960
rect 31343 32929 31355 32932
rect 31297 32923 31355 32929
rect 31386 32920 31392 32932
rect 31444 32920 31450 32972
rect 35805 32963 35863 32969
rect 35805 32929 35817 32963
rect 35851 32960 35863 32963
rect 35894 32960 35900 32972
rect 35851 32932 35900 32960
rect 35851 32929 35863 32932
rect 35805 32923 35863 32929
rect 35894 32920 35900 32932
rect 35952 32920 35958 32972
rect 49326 32960 49332 32972
rect 48792 32932 49332 32960
rect 48792 32904 48820 32932
rect 49326 32920 49332 32932
rect 49384 32960 49390 32972
rect 49421 32963 49479 32969
rect 49421 32960 49433 32963
rect 49384 32932 49433 32960
rect 49384 32920 49390 32932
rect 49421 32929 49433 32932
rect 49467 32929 49479 32963
rect 49421 32923 49479 32929
rect 26421 32895 26479 32901
rect 26421 32861 26433 32895
rect 26467 32861 26479 32895
rect 26421 32855 26479 32861
rect 27249 32895 27307 32901
rect 27249 32861 27261 32895
rect 27295 32861 27307 32895
rect 27982 32892 27988 32904
rect 27943 32864 27988 32892
rect 27249 32855 27307 32861
rect 26436 32824 26464 32855
rect 27982 32852 27988 32864
rect 28040 32852 28046 32904
rect 30650 32852 30656 32904
rect 30708 32852 30714 32904
rect 34514 32852 34520 32904
rect 34572 32892 34578 32904
rect 34793 32895 34851 32901
rect 34793 32892 34805 32895
rect 34572 32864 34805 32892
rect 34572 32852 34578 32864
rect 34793 32861 34805 32864
rect 34839 32861 34851 32895
rect 34793 32855 34851 32861
rect 35161 32895 35219 32901
rect 35161 32861 35173 32895
rect 35207 32892 35219 32895
rect 35710 32892 35716 32904
rect 35207 32864 35716 32892
rect 35207 32861 35219 32864
rect 35161 32855 35219 32861
rect 35710 32852 35716 32864
rect 35768 32852 35774 32904
rect 37274 32852 37280 32904
rect 37332 32892 37338 32904
rect 37921 32895 37979 32901
rect 37921 32892 37933 32895
rect 37332 32864 37933 32892
rect 37332 32852 37338 32864
rect 37921 32861 37933 32864
rect 37967 32892 37979 32895
rect 37967 32864 41414 32892
rect 37967 32861 37979 32864
rect 37921 32855 37979 32861
rect 27522 32824 27528 32836
rect 26436 32796 27384 32824
rect 27483 32796 27528 32824
rect 20349 32759 20407 32765
rect 20349 32725 20361 32759
rect 20395 32756 20407 32759
rect 24762 32756 24768 32768
rect 20395 32728 24768 32756
rect 20395 32725 20407 32728
rect 20349 32719 20407 32725
rect 24762 32716 24768 32728
rect 24820 32716 24826 32768
rect 26789 32759 26847 32765
rect 26789 32725 26801 32759
rect 26835 32756 26847 32759
rect 26970 32756 26976 32768
rect 26835 32728 26976 32756
rect 26835 32725 26847 32728
rect 26789 32719 26847 32725
rect 26970 32716 26976 32728
rect 27028 32716 27034 32768
rect 27356 32765 27384 32796
rect 27522 32784 27528 32796
rect 27580 32784 27586 32836
rect 38286 32784 38292 32836
rect 38344 32824 38350 32836
rect 38473 32827 38531 32833
rect 38473 32824 38485 32827
rect 38344 32796 38485 32824
rect 38344 32784 38350 32796
rect 38473 32793 38485 32796
rect 38519 32793 38531 32827
rect 41386 32824 41414 32864
rect 44910 32852 44916 32904
rect 44968 32892 44974 32904
rect 45005 32895 45063 32901
rect 45005 32892 45017 32895
rect 44968 32864 45017 32892
rect 44968 32852 44974 32864
rect 45005 32861 45017 32864
rect 45051 32861 45063 32895
rect 45186 32892 45192 32904
rect 45147 32864 45192 32892
rect 45005 32855 45063 32861
rect 45186 32852 45192 32864
rect 45244 32852 45250 32904
rect 45830 32892 45836 32904
rect 45791 32864 45836 32892
rect 45830 32852 45836 32864
rect 45888 32852 45894 32904
rect 46198 32892 46204 32904
rect 46159 32864 46204 32892
rect 46198 32852 46204 32864
rect 46256 32852 46262 32904
rect 48774 32892 48780 32904
rect 48735 32864 48780 32892
rect 48774 32852 48780 32864
rect 48832 32852 48838 32904
rect 48958 32892 48964 32904
rect 48919 32864 48964 32892
rect 48958 32852 48964 32864
rect 49016 32852 49022 32904
rect 47026 32824 47032 32836
rect 41386 32796 47032 32824
rect 38473 32787 38531 32793
rect 47026 32784 47032 32796
rect 47084 32784 47090 32836
rect 47673 32827 47731 32833
rect 47673 32793 47685 32827
rect 47719 32824 47731 32827
rect 52914 32824 52920 32836
rect 47719 32796 52920 32824
rect 47719 32793 47731 32796
rect 47673 32787 47731 32793
rect 52914 32784 52920 32796
rect 52972 32784 52978 32836
rect 27341 32759 27399 32765
rect 27341 32725 27353 32759
rect 27387 32756 27399 32759
rect 27890 32756 27896 32768
rect 27387 32728 27896 32756
rect 27387 32725 27399 32728
rect 27341 32719 27399 32725
rect 27890 32716 27896 32728
rect 27948 32716 27954 32768
rect 33594 32716 33600 32768
rect 33652 32756 33658 32768
rect 35526 32756 35532 32768
rect 33652 32728 35532 32756
rect 33652 32716 33658 32728
rect 35526 32716 35532 32728
rect 35584 32716 35590 32768
rect 38933 32759 38991 32765
rect 38933 32725 38945 32759
rect 38979 32756 38991 32759
rect 39022 32756 39028 32768
rect 38979 32728 39028 32756
rect 38979 32725 38991 32728
rect 38933 32719 38991 32725
rect 39022 32716 39028 32728
rect 39080 32716 39086 32768
rect 45097 32759 45155 32765
rect 45097 32725 45109 32759
rect 45143 32756 45155 32759
rect 45646 32756 45652 32768
rect 45143 32728 45652 32756
rect 45143 32725 45155 32728
rect 45097 32719 45155 32725
rect 45646 32716 45652 32728
rect 45704 32716 45710 32768
rect 1104 32666 58880 32688
rect 1104 32614 19574 32666
rect 19626 32614 19638 32666
rect 19690 32614 19702 32666
rect 19754 32614 19766 32666
rect 19818 32614 19830 32666
rect 19882 32614 50294 32666
rect 50346 32614 50358 32666
rect 50410 32614 50422 32666
rect 50474 32614 50486 32666
rect 50538 32614 50550 32666
rect 50602 32614 58880 32666
rect 1104 32592 58880 32614
rect 2222 32512 2228 32564
rect 2280 32552 2286 32564
rect 33594 32552 33600 32564
rect 2280 32524 33600 32552
rect 2280 32512 2286 32524
rect 33594 32512 33600 32524
rect 33652 32512 33658 32564
rect 37458 32552 37464 32564
rect 33796 32524 37464 32552
rect 8938 32444 8944 32496
rect 8996 32484 9002 32496
rect 9306 32484 9312 32496
rect 8996 32456 9312 32484
rect 8996 32444 9002 32456
rect 9306 32444 9312 32456
rect 9364 32484 9370 32496
rect 9493 32487 9551 32493
rect 9493 32484 9505 32487
rect 9364 32456 9505 32484
rect 9364 32444 9370 32456
rect 9493 32453 9505 32456
rect 9539 32453 9551 32487
rect 9493 32447 9551 32453
rect 15289 32487 15347 32493
rect 15289 32453 15301 32487
rect 15335 32484 15347 32487
rect 15838 32484 15844 32496
rect 15335 32456 15844 32484
rect 15335 32453 15347 32456
rect 15289 32447 15347 32453
rect 15838 32444 15844 32456
rect 15896 32444 15902 32496
rect 16868 32456 18552 32484
rect 7374 32416 7380 32428
rect 7335 32388 7380 32416
rect 7374 32376 7380 32388
rect 7432 32376 7438 32428
rect 8110 32416 8116 32428
rect 8071 32388 8116 32416
rect 8110 32376 8116 32388
rect 8168 32376 8174 32428
rect 10410 32416 10416 32428
rect 10371 32388 10416 32416
rect 10410 32376 10416 32388
rect 10468 32376 10474 32428
rect 13262 32416 13268 32428
rect 13223 32388 13268 32416
rect 13262 32376 13268 32388
rect 13320 32376 13326 32428
rect 13722 32376 13728 32428
rect 13780 32416 13786 32428
rect 13909 32419 13967 32425
rect 13909 32416 13921 32419
rect 13780 32388 13921 32416
rect 13780 32376 13786 32388
rect 13909 32385 13921 32388
rect 13955 32385 13967 32419
rect 15194 32416 15200 32428
rect 15155 32388 15200 32416
rect 13909 32379 13967 32385
rect 15194 32376 15200 32388
rect 15252 32376 15258 32428
rect 15381 32419 15439 32425
rect 15381 32385 15393 32419
rect 15427 32385 15439 32419
rect 15381 32379 15439 32385
rect 9033 32351 9091 32357
rect 9033 32317 9045 32351
rect 9079 32348 9091 32351
rect 10226 32348 10232 32360
rect 9079 32320 10232 32348
rect 9079 32317 9091 32320
rect 9033 32311 9091 32317
rect 10226 32308 10232 32320
rect 10284 32308 10290 32360
rect 10686 32348 10692 32360
rect 10647 32320 10692 32348
rect 10686 32308 10692 32320
rect 10744 32308 10750 32360
rect 15102 32308 15108 32360
rect 15160 32348 15166 32360
rect 15396 32348 15424 32379
rect 15654 32376 15660 32428
rect 15712 32416 15718 32428
rect 16669 32419 16727 32425
rect 16669 32416 16681 32419
rect 15712 32388 16681 32416
rect 15712 32376 15718 32388
rect 16669 32385 16681 32388
rect 16715 32385 16727 32419
rect 16669 32379 16727 32385
rect 16868 32348 16896 32456
rect 18524 32428 18552 32456
rect 18598 32444 18604 32496
rect 18656 32484 18662 32496
rect 18693 32487 18751 32493
rect 18693 32484 18705 32487
rect 18656 32456 18705 32484
rect 18656 32444 18662 32456
rect 18693 32453 18705 32456
rect 18739 32453 18751 32487
rect 24394 32484 24400 32496
rect 24355 32456 24400 32484
rect 18693 32447 18751 32453
rect 24394 32444 24400 32456
rect 24452 32444 24458 32496
rect 24581 32487 24639 32493
rect 24581 32453 24593 32487
rect 24627 32484 24639 32487
rect 24670 32484 24676 32496
rect 24627 32456 24676 32484
rect 24627 32453 24639 32456
rect 24581 32447 24639 32453
rect 24670 32444 24676 32456
rect 24728 32444 24734 32496
rect 24762 32444 24768 32496
rect 24820 32484 24826 32496
rect 30561 32487 30619 32493
rect 24820 32456 28994 32484
rect 24820 32444 24826 32456
rect 18230 32416 18236 32428
rect 18191 32388 18236 32416
rect 18230 32376 18236 32388
rect 18288 32376 18294 32428
rect 18322 32376 18328 32428
rect 18380 32416 18386 32428
rect 18380 32388 18425 32416
rect 18380 32376 18386 32388
rect 18506 32376 18512 32428
rect 18564 32416 18570 32428
rect 24210 32416 24216 32428
rect 18564 32388 18657 32416
rect 21100 32388 24216 32416
rect 18564 32376 18570 32388
rect 15160 32320 16896 32348
rect 17129 32351 17187 32357
rect 15160 32308 15166 32320
rect 17129 32317 17141 32351
rect 17175 32348 17187 32351
rect 21100 32348 21128 32388
rect 24210 32376 24216 32388
rect 24268 32416 24274 32428
rect 24268 32388 24361 32416
rect 24268 32376 24274 32388
rect 22002 32348 22008 32360
rect 17175 32320 21128 32348
rect 21963 32320 22008 32348
rect 17175 32317 17187 32320
rect 17129 32311 17187 32317
rect 22002 32308 22008 32320
rect 22060 32308 22066 32360
rect 22462 32348 22468 32360
rect 22423 32320 22468 32348
rect 22462 32308 22468 32320
rect 22520 32308 22526 32360
rect 8386 32240 8392 32292
rect 8444 32280 8450 32292
rect 15286 32280 15292 32292
rect 8444 32252 15292 32280
rect 8444 32240 8450 32252
rect 15286 32240 15292 32252
rect 15344 32240 15350 32292
rect 16206 32240 16212 32292
rect 16264 32280 16270 32292
rect 22094 32280 22100 32292
rect 16264 32252 22100 32280
rect 16264 32240 16270 32252
rect 22094 32240 22100 32252
rect 22152 32240 22158 32292
rect 22278 32280 22284 32292
rect 22239 32252 22284 32280
rect 22278 32240 22284 32252
rect 22336 32240 22342 32292
rect 28966 32280 28994 32456
rect 30561 32453 30573 32487
rect 30607 32484 30619 32487
rect 31202 32484 31208 32496
rect 30607 32456 31208 32484
rect 30607 32453 30619 32456
rect 30561 32447 30619 32453
rect 31202 32444 31208 32456
rect 31260 32444 31266 32496
rect 33796 32484 33824 32524
rect 37458 32512 37464 32524
rect 37516 32512 37522 32564
rect 38286 32552 38292 32564
rect 38247 32524 38292 32552
rect 38286 32512 38292 32524
rect 38344 32512 38350 32564
rect 40034 32552 40040 32564
rect 39995 32524 40040 32552
rect 40034 32512 40040 32524
rect 40092 32512 40098 32564
rect 45557 32555 45615 32561
rect 45557 32521 45569 32555
rect 45603 32552 45615 32555
rect 46198 32552 46204 32564
rect 45603 32524 46204 32552
rect 45603 32521 45615 32524
rect 45557 32515 45615 32521
rect 46198 32512 46204 32524
rect 46256 32512 46262 32564
rect 48958 32512 48964 32564
rect 49016 32552 49022 32564
rect 49513 32555 49571 32561
rect 49513 32552 49525 32555
rect 49016 32524 49525 32552
rect 49016 32512 49022 32524
rect 49513 32521 49525 32524
rect 49559 32521 49571 32555
rect 49513 32515 49571 32521
rect 31726 32456 33824 32484
rect 33873 32487 33931 32493
rect 30466 32416 30472 32428
rect 30427 32388 30472 32416
rect 30466 32376 30472 32388
rect 30524 32376 30530 32428
rect 30650 32416 30656 32428
rect 30611 32388 30656 32416
rect 30650 32376 30656 32388
rect 30708 32376 30714 32428
rect 31726 32348 31754 32456
rect 33873 32453 33885 32487
rect 33919 32484 33931 32487
rect 34609 32487 34667 32493
rect 33919 32456 34560 32484
rect 33919 32453 33931 32456
rect 33873 32447 33931 32453
rect 34532 32428 34560 32456
rect 34609 32453 34621 32487
rect 34655 32484 34667 32487
rect 35710 32484 35716 32496
rect 34655 32456 35716 32484
rect 34655 32453 34667 32456
rect 34609 32447 34667 32453
rect 35710 32444 35716 32456
rect 35768 32444 35774 32496
rect 56686 32484 56692 32496
rect 35820 32456 56692 32484
rect 33778 32416 33784 32428
rect 33739 32388 33784 32416
rect 33778 32376 33784 32388
rect 33836 32376 33842 32428
rect 33962 32416 33968 32428
rect 33923 32388 33968 32416
rect 33962 32376 33968 32388
rect 34020 32376 34026 32428
rect 34514 32416 34520 32428
rect 34475 32388 34520 32416
rect 34514 32376 34520 32388
rect 34572 32376 34578 32428
rect 34793 32419 34851 32425
rect 34793 32385 34805 32419
rect 34839 32385 34851 32419
rect 34793 32379 34851 32385
rect 30944 32320 31754 32348
rect 30944 32280 30972 32320
rect 34146 32308 34152 32360
rect 34204 32348 34210 32360
rect 34808 32348 34836 32379
rect 35820 32348 35848 32456
rect 56686 32444 56692 32456
rect 56744 32444 56750 32496
rect 37274 32416 37280 32428
rect 37235 32388 37280 32416
rect 37274 32376 37280 32388
rect 37332 32376 37338 32428
rect 38194 32416 38200 32428
rect 38155 32388 38200 32416
rect 38194 32376 38200 32388
rect 38252 32376 38258 32428
rect 38381 32419 38439 32425
rect 38381 32385 38393 32419
rect 38427 32385 38439 32419
rect 39022 32416 39028 32428
rect 38983 32388 39028 32416
rect 38381 32379 38439 32385
rect 37458 32348 37464 32360
rect 34204 32320 34836 32348
rect 34900 32320 35848 32348
rect 37419 32320 37464 32348
rect 34204 32308 34210 32320
rect 34900 32280 34928 32320
rect 37458 32308 37464 32320
rect 37516 32308 37522 32360
rect 24504 32252 28028 32280
rect 28966 32252 30972 32280
rect 31726 32252 34928 32280
rect 34977 32283 35035 32289
rect 10502 32212 10508 32224
rect 10463 32184 10508 32212
rect 10502 32172 10508 32184
rect 10560 32172 10566 32224
rect 10597 32215 10655 32221
rect 10597 32181 10609 32215
rect 10643 32212 10655 32215
rect 14274 32212 14280 32224
rect 10643 32184 14280 32212
rect 10643 32181 10655 32184
rect 10597 32175 10655 32181
rect 14274 32172 14280 32184
rect 14332 32172 14338 32224
rect 14369 32215 14427 32221
rect 14369 32181 14381 32215
rect 14415 32212 14427 32215
rect 14458 32212 14464 32224
rect 14415 32184 14464 32212
rect 14415 32181 14427 32184
rect 14369 32175 14427 32181
rect 14458 32172 14464 32184
rect 14516 32172 14522 32224
rect 16482 32172 16488 32224
rect 16540 32212 16546 32224
rect 16761 32215 16819 32221
rect 16761 32212 16773 32215
rect 16540 32184 16773 32212
rect 16540 32172 16546 32184
rect 16761 32181 16773 32184
rect 16807 32181 16819 32215
rect 16761 32175 16819 32181
rect 17126 32172 17132 32224
rect 17184 32212 17190 32224
rect 17589 32215 17647 32221
rect 17589 32212 17601 32215
rect 17184 32184 17601 32212
rect 17184 32172 17190 32184
rect 17589 32181 17601 32184
rect 17635 32181 17647 32215
rect 17589 32175 17647 32181
rect 21174 32172 21180 32224
rect 21232 32212 21238 32224
rect 24504 32212 24532 32252
rect 21232 32184 24532 32212
rect 27065 32215 27123 32221
rect 21232 32172 21238 32184
rect 27065 32181 27077 32215
rect 27111 32212 27123 32215
rect 27709 32215 27767 32221
rect 27709 32212 27721 32215
rect 27111 32184 27721 32212
rect 27111 32181 27123 32184
rect 27065 32175 27123 32181
rect 27709 32181 27721 32184
rect 27755 32212 27767 32215
rect 27890 32212 27896 32224
rect 27755 32184 27896 32212
rect 27755 32181 27767 32184
rect 27709 32175 27767 32181
rect 27890 32172 27896 32184
rect 27948 32172 27954 32224
rect 28000 32212 28028 32252
rect 31726 32212 31754 32252
rect 34977 32249 34989 32283
rect 35023 32280 35035 32283
rect 38010 32280 38016 32292
rect 35023 32252 38016 32280
rect 35023 32249 35035 32252
rect 34977 32243 35035 32249
rect 38010 32240 38016 32252
rect 38068 32280 38074 32292
rect 38396 32280 38424 32379
rect 39022 32376 39028 32388
rect 39080 32376 39086 32428
rect 39206 32416 39212 32428
rect 39167 32388 39212 32416
rect 39206 32376 39212 32388
rect 39264 32376 39270 32428
rect 41322 32416 41328 32428
rect 41283 32388 41328 32416
rect 41322 32376 41328 32388
rect 41380 32376 41386 32428
rect 43346 32416 43352 32428
rect 43307 32388 43352 32416
rect 43346 32376 43352 32388
rect 43404 32376 43410 32428
rect 44910 32376 44916 32428
rect 44968 32416 44974 32428
rect 45281 32419 45339 32425
rect 45281 32416 45293 32419
rect 44968 32388 45293 32416
rect 44968 32376 44974 32388
rect 45281 32385 45293 32388
rect 45327 32385 45339 32419
rect 45646 32416 45652 32428
rect 45607 32388 45652 32416
rect 45281 32379 45339 32385
rect 45646 32376 45652 32388
rect 45704 32376 45710 32428
rect 47946 32376 47952 32428
rect 48004 32416 48010 32428
rect 48685 32419 48743 32425
rect 48685 32416 48697 32419
rect 48004 32388 48697 32416
rect 48004 32376 48010 32388
rect 48685 32385 48697 32388
rect 48731 32385 48743 32419
rect 48685 32379 48743 32385
rect 49145 32419 49203 32425
rect 49145 32385 49157 32419
rect 49191 32416 49203 32419
rect 49786 32416 49792 32428
rect 49191 32388 49792 32416
rect 49191 32385 49203 32388
rect 49145 32379 49203 32385
rect 49786 32376 49792 32388
rect 49844 32376 49850 32428
rect 52914 32416 52920 32428
rect 52875 32388 52920 32416
rect 52914 32376 52920 32388
rect 52972 32376 52978 32428
rect 41230 32348 41236 32360
rect 41191 32320 41236 32348
rect 41230 32308 41236 32320
rect 41288 32308 41294 32360
rect 41693 32351 41751 32357
rect 41693 32317 41705 32351
rect 41739 32348 41751 32351
rect 41782 32348 41788 32360
rect 41739 32320 41788 32348
rect 41739 32317 41751 32320
rect 41693 32311 41751 32317
rect 41782 32308 41788 32320
rect 41840 32308 41846 32360
rect 43441 32351 43499 32357
rect 43441 32317 43453 32351
rect 43487 32348 43499 32351
rect 45094 32348 45100 32360
rect 43487 32320 43668 32348
rect 45007 32320 45100 32348
rect 43487 32317 43499 32320
rect 43441 32311 43499 32317
rect 38068 32252 38424 32280
rect 38068 32240 38074 32252
rect 28000 32184 31754 32212
rect 43640 32212 43668 32320
rect 45094 32308 45100 32320
rect 45152 32308 45158 32360
rect 53101 32351 53159 32357
rect 53101 32317 53113 32351
rect 53147 32348 53159 32351
rect 53282 32348 53288 32360
rect 53147 32320 53288 32348
rect 53147 32317 53159 32320
rect 53101 32311 53159 32317
rect 53282 32308 53288 32320
rect 53340 32308 53346 32360
rect 43717 32283 43775 32289
rect 43717 32249 43729 32283
rect 43763 32280 43775 32283
rect 45112 32280 45140 32308
rect 43763 32252 45140 32280
rect 43763 32249 43775 32252
rect 43717 32243 43775 32249
rect 45186 32212 45192 32224
rect 43640 32184 45192 32212
rect 45186 32172 45192 32184
rect 45244 32172 45250 32224
rect 52730 32212 52736 32224
rect 52691 32184 52736 32212
rect 52730 32172 52736 32184
rect 52788 32172 52794 32224
rect 1104 32122 58880 32144
rect 1104 32070 4214 32122
rect 4266 32070 4278 32122
rect 4330 32070 4342 32122
rect 4394 32070 4406 32122
rect 4458 32070 4470 32122
rect 4522 32070 34934 32122
rect 34986 32070 34998 32122
rect 35050 32070 35062 32122
rect 35114 32070 35126 32122
rect 35178 32070 35190 32122
rect 35242 32070 58880 32122
rect 1104 32048 58880 32070
rect 1670 31968 1676 32020
rect 1728 32008 1734 32020
rect 2501 32011 2559 32017
rect 2501 32008 2513 32011
rect 1728 31980 2513 32008
rect 1728 31968 1734 31980
rect 2501 31977 2513 31980
rect 2547 31977 2559 32011
rect 8386 32008 8392 32020
rect 8347 31980 8392 32008
rect 2501 31971 2559 31977
rect 8386 31968 8392 31980
rect 8444 31968 8450 32020
rect 8754 31968 8760 32020
rect 8812 32008 8818 32020
rect 9306 32008 9312 32020
rect 8812 31980 9312 32008
rect 8812 31968 8818 31980
rect 9306 31968 9312 31980
rect 9364 31968 9370 32020
rect 10042 31968 10048 32020
rect 10100 32008 10106 32020
rect 10410 32008 10416 32020
rect 10100 31980 10416 32008
rect 10100 31968 10106 31980
rect 10410 31968 10416 31980
rect 10468 32008 10474 32020
rect 10597 32011 10655 32017
rect 10597 32008 10609 32011
rect 10468 31980 10609 32008
rect 10468 31968 10474 31980
rect 10597 31977 10609 31980
rect 10643 31977 10655 32011
rect 13265 32011 13323 32017
rect 10597 31971 10655 31977
rect 10888 31980 12434 32008
rect 10137 31943 10195 31949
rect 10137 31909 10149 31943
rect 10183 31940 10195 31943
rect 10888 31940 10916 31980
rect 10183 31912 10916 31940
rect 10965 31943 11023 31949
rect 10183 31909 10195 31912
rect 10137 31903 10195 31909
rect 10965 31909 10977 31943
rect 11011 31909 11023 31943
rect 12406 31940 12434 31980
rect 13265 31977 13277 32011
rect 13311 32008 13323 32011
rect 15194 32008 15200 32020
rect 13311 31980 15200 32008
rect 13311 31977 13323 31980
rect 13265 31971 13323 31977
rect 15194 31968 15200 31980
rect 15252 31968 15258 32020
rect 15654 32008 15660 32020
rect 15615 31980 15660 32008
rect 15654 31968 15660 31980
rect 15712 31968 15718 32020
rect 16301 32011 16359 32017
rect 16301 31977 16313 32011
rect 16347 31977 16359 32011
rect 16482 32008 16488 32020
rect 16443 31980 16488 32008
rect 16301 31971 16359 31977
rect 14182 31940 14188 31952
rect 12406 31912 14188 31940
rect 10965 31903 11023 31909
rect 9401 31875 9459 31881
rect 9401 31841 9413 31875
rect 9447 31872 9459 31875
rect 9766 31872 9772 31884
rect 9447 31844 9772 31872
rect 9447 31841 9459 31844
rect 9401 31835 9459 31841
rect 9766 31832 9772 31844
rect 9824 31832 9830 31884
rect 9861 31875 9919 31881
rect 9861 31841 9873 31875
rect 9907 31872 9919 31875
rect 9950 31872 9956 31884
rect 9907 31844 9956 31872
rect 9907 31841 9919 31844
rect 9861 31835 9919 31841
rect 9950 31832 9956 31844
rect 10008 31872 10014 31884
rect 10686 31872 10692 31884
rect 10008 31844 10692 31872
rect 10008 31832 10014 31844
rect 10686 31832 10692 31844
rect 10744 31832 10750 31884
rect 10980 31872 11008 31903
rect 14182 31900 14188 31912
rect 14240 31900 14246 31952
rect 14274 31900 14280 31952
rect 14332 31940 14338 31952
rect 16316 31940 16344 31971
rect 16482 31968 16488 31980
rect 16540 31968 16546 32020
rect 16574 31968 16580 32020
rect 16632 32008 16638 32020
rect 17034 32008 17040 32020
rect 16632 31980 17040 32008
rect 16632 31968 16638 31980
rect 17034 31968 17040 31980
rect 17092 31968 17098 32020
rect 18230 31968 18236 32020
rect 18288 32008 18294 32020
rect 18417 32011 18475 32017
rect 18417 32008 18429 32011
rect 18288 31980 18429 32008
rect 18288 31968 18294 31980
rect 18417 31977 18429 31980
rect 18463 31977 18475 32011
rect 22557 32011 22615 32017
rect 22557 32008 22569 32011
rect 18417 31971 18475 31977
rect 22066 31980 22569 32008
rect 14332 31912 16344 31940
rect 14332 31900 14338 31912
rect 10980 31844 15056 31872
rect 1946 31764 1952 31816
rect 2004 31804 2010 31816
rect 2041 31807 2099 31813
rect 2041 31804 2053 31807
rect 2004 31776 2053 31804
rect 2004 31764 2010 31776
rect 2041 31773 2053 31776
rect 2087 31773 2099 31807
rect 2041 31767 2099 31773
rect 2685 31807 2743 31813
rect 2685 31773 2697 31807
rect 2731 31804 2743 31807
rect 3145 31807 3203 31813
rect 3145 31804 3157 31807
rect 2731 31776 3157 31804
rect 2731 31773 2743 31776
rect 2685 31767 2743 31773
rect 3145 31773 3157 31776
rect 3191 31804 3203 31807
rect 3234 31804 3240 31816
rect 3191 31776 3240 31804
rect 3191 31773 3203 31776
rect 3145 31767 3203 31773
rect 3234 31764 3240 31776
rect 3292 31764 3298 31816
rect 7101 31807 7159 31813
rect 7101 31773 7113 31807
rect 7147 31773 7159 31807
rect 7101 31767 7159 31773
rect 1578 31696 1584 31748
rect 1636 31736 1642 31748
rect 1857 31739 1915 31745
rect 1857 31736 1869 31739
rect 1636 31708 1869 31736
rect 1636 31696 1642 31708
rect 1857 31705 1869 31708
rect 1903 31705 1915 31739
rect 7116 31736 7144 31767
rect 7190 31764 7196 31816
rect 7248 31804 7254 31816
rect 7561 31807 7619 31813
rect 7561 31804 7573 31807
rect 7248 31776 7573 31804
rect 7248 31764 7254 31776
rect 7561 31773 7573 31776
rect 7607 31773 7619 31807
rect 7561 31767 7619 31773
rect 8202 31764 8208 31816
rect 8260 31804 8266 31816
rect 9125 31807 9183 31813
rect 9125 31804 9137 31807
rect 8260 31776 9137 31804
rect 8260 31764 8266 31776
rect 9125 31773 9137 31776
rect 9171 31773 9183 31807
rect 10042 31804 10048 31816
rect 10003 31776 10048 31804
rect 9125 31767 9183 31773
rect 10042 31764 10048 31776
rect 10100 31764 10106 31816
rect 10134 31764 10140 31816
rect 10192 31804 10198 31816
rect 10502 31804 10508 31816
rect 10192 31776 10508 31804
rect 10192 31764 10198 31776
rect 10502 31764 10508 31776
rect 10560 31804 10566 31816
rect 10597 31807 10655 31813
rect 10597 31804 10609 31807
rect 10560 31776 10609 31804
rect 10560 31764 10566 31776
rect 10597 31773 10609 31776
rect 10643 31773 10655 31807
rect 13538 31804 13544 31816
rect 13499 31776 13544 31804
rect 10597 31767 10655 31773
rect 13538 31764 13544 31776
rect 13596 31764 13602 31816
rect 7282 31736 7288 31748
rect 7116 31708 7288 31736
rect 1857 31699 1915 31705
rect 7282 31696 7288 31708
rect 7340 31696 7346 31748
rect 13265 31739 13323 31745
rect 13265 31705 13277 31739
rect 13311 31736 13323 31739
rect 13354 31736 13360 31748
rect 13311 31708 13360 31736
rect 13311 31705 13323 31708
rect 13265 31699 13323 31705
rect 13354 31696 13360 31708
rect 13412 31696 13418 31748
rect 15028 31736 15056 31844
rect 15212 31813 15240 31912
rect 17218 31900 17224 31952
rect 17276 31940 17282 31952
rect 20165 31943 20223 31949
rect 20165 31940 20177 31943
rect 17276 31912 20177 31940
rect 17276 31900 17282 31912
rect 20165 31909 20177 31912
rect 20211 31909 20223 31943
rect 22066 31940 22094 31980
rect 22557 31977 22569 31980
rect 22603 32008 22615 32011
rect 23293 32011 23351 32017
rect 23293 32008 23305 32011
rect 22603 31980 23305 32008
rect 22603 31977 22615 31980
rect 22557 31971 22615 31977
rect 23293 31977 23305 31980
rect 23339 31977 23351 32011
rect 23293 31971 23351 31977
rect 26789 32011 26847 32017
rect 26789 31977 26801 32011
rect 26835 32008 26847 32011
rect 27062 32008 27068 32020
rect 26835 31980 27068 32008
rect 26835 31977 26847 31980
rect 26789 31971 26847 31977
rect 27062 31968 27068 31980
rect 27120 32008 27126 32020
rect 27522 32008 27528 32020
rect 27120 31980 27528 32008
rect 27120 31968 27126 31980
rect 27522 31968 27528 31980
rect 27580 31968 27586 32020
rect 32585 32011 32643 32017
rect 32585 31977 32597 32011
rect 32631 32008 32643 32011
rect 33962 32008 33968 32020
rect 32631 31980 33968 32008
rect 32631 31977 32643 31980
rect 32585 31971 32643 31977
rect 33962 31968 33968 31980
rect 34020 31968 34026 32020
rect 34146 32008 34152 32020
rect 34107 31980 34152 32008
rect 34146 31968 34152 31980
rect 34204 31968 34210 32020
rect 41785 32011 41843 32017
rect 41785 31977 41797 32011
rect 41831 32008 41843 32011
rect 43346 32008 43352 32020
rect 41831 31980 43352 32008
rect 41831 31977 41843 31980
rect 41785 31971 41843 31977
rect 43346 31968 43352 31980
rect 43404 32008 43410 32020
rect 45002 32008 45008 32020
rect 43404 31980 45008 32008
rect 43404 31968 43410 31980
rect 45002 31968 45008 31980
rect 45060 31968 45066 32020
rect 47946 32008 47952 32020
rect 47907 31980 47952 32008
rect 47946 31968 47952 31980
rect 48004 31968 48010 32020
rect 49050 32008 49056 32020
rect 49011 31980 49056 32008
rect 49050 31968 49056 31980
rect 49108 31968 49114 32020
rect 53282 31968 53288 32020
rect 53340 32008 53346 32020
rect 53340 31980 55214 32008
rect 53340 31968 53346 31980
rect 20165 31903 20223 31909
rect 20824 31912 22094 31940
rect 22741 31943 22799 31949
rect 15197 31807 15255 31813
rect 15197 31773 15209 31807
rect 15243 31773 15255 31807
rect 15197 31767 15255 31773
rect 15473 31807 15531 31813
rect 15473 31773 15485 31807
rect 15519 31804 15531 31807
rect 16206 31804 16212 31816
rect 15519 31776 16212 31804
rect 15519 31773 15531 31776
rect 15473 31767 15531 31773
rect 16206 31764 16212 31776
rect 16264 31764 16270 31816
rect 17954 31804 17960 31816
rect 17915 31776 17960 31804
rect 17954 31764 17960 31776
rect 18012 31764 18018 31816
rect 18046 31764 18052 31816
rect 18104 31804 18110 31816
rect 18233 31807 18291 31813
rect 18233 31804 18245 31807
rect 18104 31776 18245 31804
rect 18104 31764 18110 31776
rect 18233 31773 18245 31776
rect 18279 31773 18291 31807
rect 20180 31804 20208 31903
rect 20824 31813 20852 31912
rect 22741 31909 22753 31943
rect 22787 31940 22799 31943
rect 30466 31940 30472 31952
rect 22787 31912 30472 31940
rect 22787 31909 22799 31912
rect 22741 31903 22799 31909
rect 30466 31900 30472 31912
rect 30524 31900 30530 31952
rect 32122 31900 32128 31952
rect 32180 31940 32186 31952
rect 32401 31943 32459 31949
rect 32401 31940 32413 31943
rect 32180 31912 32413 31940
rect 32180 31900 32186 31912
rect 32401 31909 32413 31912
rect 32447 31909 32459 31943
rect 33980 31940 34008 31968
rect 33980 31912 38792 31940
rect 32401 31903 32459 31909
rect 20990 31832 20996 31884
rect 21048 31872 21054 31884
rect 21821 31875 21879 31881
rect 21048 31844 21496 31872
rect 21048 31832 21054 31844
rect 20809 31807 20867 31813
rect 20809 31804 20821 31807
rect 20180 31776 20821 31804
rect 18233 31767 18291 31773
rect 20809 31773 20821 31776
rect 20855 31773 20867 31807
rect 21468 31804 21496 31844
rect 21821 31841 21833 31875
rect 21867 31872 21879 31875
rect 22002 31872 22008 31884
rect 21867 31844 22008 31872
rect 21867 31841 21879 31844
rect 21821 31835 21879 31841
rect 22002 31832 22008 31844
rect 22060 31832 22066 31884
rect 24210 31832 24216 31884
rect 24268 31872 24274 31884
rect 24489 31875 24547 31881
rect 24489 31872 24501 31875
rect 24268 31844 24501 31872
rect 24268 31832 24274 31844
rect 24489 31841 24501 31844
rect 24535 31841 24547 31875
rect 24489 31835 24547 31841
rect 24949 31875 25007 31881
rect 24949 31841 24961 31875
rect 24995 31872 25007 31875
rect 26878 31872 26884 31884
rect 24995 31844 26884 31872
rect 24995 31841 25007 31844
rect 24949 31835 25007 31841
rect 26878 31832 26884 31844
rect 26936 31832 26942 31884
rect 28626 31872 28632 31884
rect 26988 31844 28632 31872
rect 26988 31816 27016 31844
rect 28626 31832 28632 31844
rect 28684 31832 28690 31884
rect 30650 31872 30656 31884
rect 30611 31844 30656 31872
rect 30650 31832 30656 31844
rect 30708 31832 30714 31884
rect 35710 31872 35716 31884
rect 34164 31844 34928 31872
rect 35671 31844 35716 31872
rect 29736 31816 29788 31822
rect 34164 31816 34192 31844
rect 22281 31807 22339 31813
rect 22281 31804 22293 31807
rect 21468 31790 22293 31804
rect 21482 31776 22293 31790
rect 20809 31767 20867 31773
rect 22281 31773 22293 31776
rect 22327 31773 22339 31807
rect 22281 31767 22339 31773
rect 24394 31764 24400 31816
rect 24452 31804 24458 31816
rect 24581 31807 24639 31813
rect 24581 31804 24593 31807
rect 24452 31776 24593 31804
rect 24452 31764 24458 31776
rect 24581 31773 24593 31776
rect 24627 31773 24639 31807
rect 26970 31804 26976 31816
rect 26931 31776 26976 31804
rect 24581 31767 24639 31773
rect 26970 31764 26976 31776
rect 27028 31764 27034 31816
rect 27249 31807 27307 31813
rect 27249 31773 27261 31807
rect 27295 31804 27307 31807
rect 27433 31807 27491 31813
rect 27295 31776 27384 31804
rect 27295 31773 27307 31776
rect 27249 31767 27307 31773
rect 15289 31739 15347 31745
rect 15289 31736 15301 31739
rect 15028 31708 15301 31736
rect 15289 31705 15301 31708
rect 15335 31736 15347 31739
rect 16117 31739 16175 31745
rect 16117 31736 16129 31739
rect 15335 31708 16129 31736
rect 15335 31705 15347 31708
rect 15289 31699 15347 31705
rect 16117 31705 16129 31708
rect 16163 31705 16175 31739
rect 16224 31736 16252 31764
rect 16317 31739 16375 31745
rect 16317 31736 16329 31739
rect 16224 31708 16329 31736
rect 16117 31699 16175 31705
rect 16317 31705 16329 31708
rect 16363 31705 16375 31739
rect 27356 31736 27384 31776
rect 27433 31773 27445 31807
rect 27479 31804 27491 31807
rect 27798 31804 27804 31816
rect 27479 31776 27804 31804
rect 27479 31773 27491 31776
rect 27433 31767 27491 31773
rect 27798 31764 27804 31776
rect 27856 31764 27862 31816
rect 29641 31807 29699 31813
rect 29641 31804 29653 31807
rect 29104 31776 29653 31804
rect 28350 31736 28356 31748
rect 27356 31708 28356 31736
rect 16317 31699 16375 31705
rect 28350 31696 28356 31708
rect 28408 31696 28414 31748
rect 29104 31680 29132 31776
rect 29641 31773 29653 31776
rect 29687 31773 29699 31807
rect 29641 31767 29699 31773
rect 33962 31804 33968 31816
rect 33875 31776 33968 31804
rect 33962 31764 33968 31776
rect 34020 31804 34026 31816
rect 34020 31776 34045 31804
rect 34020 31764 34026 31776
rect 34146 31764 34152 31816
rect 34204 31804 34210 31816
rect 34793 31807 34851 31813
rect 34793 31804 34805 31807
rect 34204 31776 34297 31804
rect 34348 31776 34805 31804
rect 34204 31764 34210 31776
rect 29736 31758 29788 31764
rect 32125 31739 32183 31745
rect 32125 31705 32137 31739
rect 32171 31736 32183 31739
rect 32214 31736 32220 31748
rect 32171 31708 32220 31736
rect 32171 31705 32183 31708
rect 32125 31699 32183 31705
rect 32214 31696 32220 31708
rect 32272 31696 32278 31748
rect 33980 31736 34008 31764
rect 34348 31736 34376 31776
rect 34793 31773 34805 31776
rect 34839 31773 34851 31807
rect 34900 31790 34928 31844
rect 35710 31832 35716 31844
rect 35768 31832 35774 31884
rect 38105 31875 38163 31881
rect 38105 31841 38117 31875
rect 38151 31872 38163 31875
rect 38654 31872 38660 31884
rect 38151 31844 38660 31872
rect 38151 31841 38163 31844
rect 38105 31835 38163 31841
rect 38654 31832 38660 31844
rect 38712 31832 38718 31884
rect 38010 31804 38016 31816
rect 37971 31776 38016 31804
rect 34793 31767 34851 31773
rect 38010 31764 38016 31776
rect 38068 31764 38074 31816
rect 38194 31804 38200 31816
rect 38155 31776 38200 31804
rect 38194 31764 38200 31776
rect 38252 31764 38258 31816
rect 38764 31804 38792 31912
rect 39022 31900 39028 31952
rect 39080 31940 39086 31952
rect 39080 31912 39160 31940
rect 39080 31900 39086 31912
rect 39132 31881 39160 31912
rect 41046 31900 41052 31952
rect 41104 31940 41110 31952
rect 55186 31940 55214 31980
rect 57885 31943 57943 31949
rect 57885 31940 57897 31943
rect 41104 31912 53512 31940
rect 55186 31912 57897 31940
rect 41104 31900 41110 31912
rect 39117 31875 39175 31881
rect 39117 31841 39129 31875
rect 39163 31841 39175 31875
rect 39117 31835 39175 31841
rect 41230 31832 41236 31884
rect 41288 31832 41294 31884
rect 41322 31832 41328 31884
rect 41380 31872 41386 31884
rect 41380 31844 41920 31872
rect 41380 31832 41386 31844
rect 39025 31807 39083 31813
rect 39025 31804 39037 31807
rect 38764 31776 39037 31804
rect 39025 31773 39037 31776
rect 39071 31804 39083 31807
rect 39206 31804 39212 31816
rect 39071 31776 39212 31804
rect 39071 31773 39083 31776
rect 39025 31767 39083 31773
rect 39206 31764 39212 31776
rect 39264 31764 39270 31816
rect 39301 31807 39359 31813
rect 39301 31773 39313 31807
rect 39347 31804 39359 31807
rect 41248 31804 41276 31832
rect 41892 31813 41920 31844
rect 45646 31832 45652 31884
rect 45704 31872 45710 31884
rect 48222 31872 48228 31884
rect 45704 31844 45784 31872
rect 45704 31832 45710 31844
rect 41693 31807 41751 31813
rect 41693 31804 41705 31807
rect 39347 31776 41705 31804
rect 39347 31773 39359 31776
rect 39301 31767 39359 31773
rect 41693 31773 41705 31776
rect 41739 31773 41751 31807
rect 41693 31767 41751 31773
rect 41877 31807 41935 31813
rect 41877 31773 41889 31807
rect 41923 31773 41935 31807
rect 45094 31804 45100 31816
rect 45055 31776 45100 31804
rect 41877 31767 41935 31773
rect 45094 31764 45100 31776
rect 45152 31764 45158 31816
rect 45554 31764 45560 31816
rect 45612 31804 45618 31816
rect 45756 31813 45784 31844
rect 47872 31844 48228 31872
rect 47872 31813 47900 31844
rect 48222 31832 48228 31844
rect 48280 31832 48286 31884
rect 48406 31832 48412 31884
rect 48464 31872 48470 31884
rect 48593 31875 48651 31881
rect 48593 31872 48605 31875
rect 48464 31844 48605 31872
rect 48464 31832 48470 31844
rect 48593 31841 48605 31844
rect 48639 31841 48651 31875
rect 48593 31835 48651 31841
rect 45741 31807 45799 31813
rect 45612 31776 45657 31804
rect 45612 31764 45618 31776
rect 45741 31773 45753 31807
rect 45787 31773 45799 31807
rect 45741 31767 45799 31773
rect 47857 31807 47915 31813
rect 47857 31773 47869 31807
rect 47903 31773 47915 31807
rect 47857 31767 47915 31773
rect 48041 31807 48099 31813
rect 48041 31773 48053 31807
rect 48087 31773 48099 31807
rect 48682 31804 48688 31816
rect 48643 31776 48688 31804
rect 48041 31767 48099 31773
rect 45370 31736 45376 31748
rect 33980 31708 34376 31736
rect 45331 31708 45376 31736
rect 45370 31696 45376 31708
rect 45428 31736 45434 31748
rect 48056 31736 48084 31767
rect 48682 31764 48688 31776
rect 48740 31764 48746 31816
rect 52914 31804 52920 31816
rect 52875 31776 52920 31804
rect 52914 31764 52920 31776
rect 52972 31764 52978 31816
rect 53282 31804 53288 31816
rect 53243 31776 53288 31804
rect 53282 31764 53288 31776
rect 53340 31764 53346 31816
rect 53484 31804 53512 31912
rect 57885 31909 57897 31912
rect 57931 31909 57943 31943
rect 57885 31903 57943 31909
rect 55309 31807 55367 31813
rect 55309 31804 55321 31807
rect 53484 31776 53604 31804
rect 48590 31736 48596 31748
rect 45428 31708 48596 31736
rect 45428 31696 45434 31708
rect 48590 31696 48596 31708
rect 48648 31696 48654 31748
rect 52270 31696 52276 31748
rect 52328 31696 52334 31748
rect 53576 31736 53604 31776
rect 53760 31776 55321 31804
rect 53760 31736 53788 31776
rect 55309 31773 55321 31776
rect 55355 31773 55367 31807
rect 55309 31767 55367 31773
rect 55490 31764 55496 31816
rect 55548 31804 55554 31816
rect 55548 31776 55706 31804
rect 55548 31764 55554 31776
rect 56318 31764 56324 31816
rect 56376 31804 56382 31816
rect 57425 31807 57483 31813
rect 56376 31776 56421 31804
rect 56376 31764 56382 31776
rect 57425 31773 57437 31807
rect 57471 31804 57483 31807
rect 57882 31804 57888 31816
rect 57471 31776 57888 31804
rect 57471 31773 57483 31776
rect 57425 31767 57483 31773
rect 57882 31764 57888 31776
rect 57940 31804 57946 31816
rect 58069 31807 58127 31813
rect 58069 31804 58081 31807
rect 57940 31776 58081 31804
rect 57940 31764 57946 31776
rect 58069 31773 58081 31776
rect 58115 31773 58127 31807
rect 58069 31767 58127 31773
rect 53576 31708 53788 31736
rect 8938 31668 8944 31680
rect 8899 31640 8944 31668
rect 8938 31628 8944 31640
rect 8996 31628 9002 31680
rect 13170 31628 13176 31680
rect 13228 31668 13234 31680
rect 13449 31671 13507 31677
rect 13449 31668 13461 31671
rect 13228 31640 13461 31668
rect 13228 31628 13234 31640
rect 13449 31637 13461 31640
rect 13495 31637 13507 31671
rect 13449 31631 13507 31637
rect 18049 31671 18107 31677
rect 18049 31637 18061 31671
rect 18095 31668 18107 31671
rect 18230 31668 18236 31680
rect 18095 31640 18236 31668
rect 18095 31637 18107 31640
rect 18049 31631 18107 31637
rect 18230 31628 18236 31640
rect 18288 31628 18294 31680
rect 28997 31671 29055 31677
rect 28997 31637 29009 31671
rect 29043 31668 29055 31671
rect 29086 31668 29092 31680
rect 29043 31640 29092 31668
rect 29043 31637 29055 31640
rect 28997 31631 29055 31637
rect 29086 31628 29092 31640
rect 29144 31628 29150 31680
rect 1104 31578 58880 31600
rect 1104 31526 19574 31578
rect 19626 31526 19638 31578
rect 19690 31526 19702 31578
rect 19754 31526 19766 31578
rect 19818 31526 19830 31578
rect 19882 31526 50294 31578
rect 50346 31526 50358 31578
rect 50410 31526 50422 31578
rect 50474 31526 50486 31578
rect 50538 31526 50550 31578
rect 50602 31526 58880 31578
rect 1104 31504 58880 31526
rect 10042 31464 10048 31476
rect 10003 31436 10048 31464
rect 10042 31424 10048 31436
rect 10100 31424 10106 31476
rect 13725 31467 13783 31473
rect 13725 31433 13737 31467
rect 13771 31464 13783 31467
rect 15102 31464 15108 31476
rect 13771 31436 15108 31464
rect 13771 31433 13783 31436
rect 13725 31427 13783 31433
rect 15102 31424 15108 31436
rect 15160 31424 15166 31476
rect 32585 31467 32643 31473
rect 19536 31436 28994 31464
rect 19536 31408 19564 31436
rect 1578 31396 1584 31408
rect 1539 31368 1584 31396
rect 1578 31356 1584 31368
rect 1636 31356 1642 31408
rect 7098 31356 7104 31408
rect 7156 31396 7162 31408
rect 7285 31399 7343 31405
rect 7285 31396 7297 31399
rect 7156 31368 7297 31396
rect 7156 31356 7162 31368
rect 7285 31365 7297 31368
rect 7331 31365 7343 31399
rect 7285 31359 7343 31365
rect 7653 31399 7711 31405
rect 7653 31365 7665 31399
rect 7699 31396 7711 31399
rect 8938 31396 8944 31408
rect 7699 31368 8944 31396
rect 7699 31365 7711 31368
rect 7653 31359 7711 31365
rect 8938 31356 8944 31368
rect 8996 31356 9002 31408
rect 13354 31396 13360 31408
rect 13315 31368 13360 31396
rect 13354 31356 13360 31368
rect 13412 31356 13418 31408
rect 13538 31356 13544 31408
rect 13596 31405 13602 31408
rect 13596 31399 13615 31405
rect 13603 31365 13615 31399
rect 13596 31359 13615 31365
rect 13596 31356 13602 31359
rect 17954 31356 17960 31408
rect 18012 31396 18018 31408
rect 18012 31368 18552 31396
rect 18012 31356 18018 31368
rect 18524 31340 18552 31368
rect 19518 31356 19524 31408
rect 19576 31356 19582 31408
rect 22830 31396 22836 31408
rect 22112 31368 22836 31396
rect 7190 31328 7196 31340
rect 7151 31300 7196 31328
rect 7190 31288 7196 31300
rect 7248 31288 7254 31340
rect 8110 31328 8116 31340
rect 7392 31300 8116 31328
rect 7392 31269 7420 31300
rect 8110 31288 8116 31300
rect 8168 31288 8174 31340
rect 10042 31288 10048 31340
rect 10100 31328 10106 31340
rect 10137 31331 10195 31337
rect 10137 31328 10149 31331
rect 10100 31300 10149 31328
rect 10100 31288 10106 31300
rect 10137 31297 10149 31300
rect 10183 31297 10195 31331
rect 18046 31328 18052 31340
rect 18007 31300 18052 31328
rect 10137 31291 10195 31297
rect 18046 31288 18052 31300
rect 18104 31288 18110 31340
rect 18230 31328 18236 31340
rect 18191 31300 18236 31328
rect 18230 31288 18236 31300
rect 18288 31288 18294 31340
rect 18506 31328 18512 31340
rect 18467 31300 18512 31328
rect 18506 31288 18512 31300
rect 18564 31288 18570 31340
rect 21821 31331 21879 31337
rect 21821 31297 21833 31331
rect 21867 31297 21879 31331
rect 21821 31291 21879 31297
rect 7377 31263 7435 31269
rect 7377 31229 7389 31263
rect 7423 31229 7435 31263
rect 7377 31223 7435 31229
rect 9490 31220 9496 31272
rect 9548 31260 9554 31272
rect 9769 31263 9827 31269
rect 9769 31260 9781 31263
rect 9548 31232 9781 31260
rect 9548 31220 9554 31232
rect 9769 31229 9781 31232
rect 9815 31260 9827 31263
rect 10594 31260 10600 31272
rect 9815 31232 10600 31260
rect 9815 31229 9827 31232
rect 9769 31223 9827 31229
rect 10594 31220 10600 31232
rect 10652 31220 10658 31272
rect 18322 31220 18328 31272
rect 18380 31260 18386 31272
rect 18417 31263 18475 31269
rect 18417 31260 18429 31263
rect 18380 31232 18429 31260
rect 18380 31220 18386 31232
rect 18417 31229 18429 31232
rect 18463 31260 18475 31263
rect 21836 31260 21864 31291
rect 22112 31269 22140 31368
rect 22830 31356 22836 31368
rect 22888 31356 22894 31408
rect 27062 31396 27068 31408
rect 27023 31368 27068 31396
rect 27062 31356 27068 31368
rect 27120 31356 27126 31408
rect 27798 31356 27804 31408
rect 27856 31396 27862 31408
rect 27856 31368 28304 31396
rect 27856 31356 27862 31368
rect 28276 31337 28304 31368
rect 22189 31331 22247 31337
rect 22189 31297 22201 31331
rect 22235 31328 22247 31331
rect 27525 31331 27583 31337
rect 22235 31300 22416 31328
rect 22235 31297 22247 31300
rect 22189 31291 22247 31297
rect 18463 31232 21864 31260
rect 22097 31263 22155 31269
rect 18463 31229 18475 31232
rect 18417 31223 18475 31229
rect 22097 31229 22109 31263
rect 22143 31229 22155 31263
rect 22097 31223 22155 31229
rect 7558 31152 7564 31204
rect 7616 31192 7622 31204
rect 7837 31195 7895 31201
rect 7837 31192 7849 31195
rect 7616 31164 7849 31192
rect 7616 31152 7622 31164
rect 7837 31161 7849 31164
rect 7883 31161 7895 31195
rect 7837 31155 7895 31161
rect 22189 31195 22247 31201
rect 22189 31161 22201 31195
rect 22235 31192 22247 31195
rect 22278 31192 22284 31204
rect 22235 31164 22284 31192
rect 22235 31161 22247 31164
rect 22189 31155 22247 31161
rect 22278 31152 22284 31164
rect 22336 31152 22342 31204
rect 9858 31124 9864 31136
rect 9819 31096 9864 31124
rect 9858 31084 9864 31096
rect 9916 31084 9922 31136
rect 9953 31127 10011 31133
rect 9953 31093 9965 31127
rect 9999 31124 10011 31127
rect 10318 31124 10324 31136
rect 9999 31096 10324 31124
rect 9999 31093 10011 31096
rect 9953 31087 10011 31093
rect 10318 31084 10324 31096
rect 10376 31084 10382 31136
rect 13170 31084 13176 31136
rect 13228 31124 13234 31136
rect 13541 31127 13599 31133
rect 13541 31124 13553 31127
rect 13228 31096 13553 31124
rect 13228 31084 13234 31096
rect 13541 31093 13553 31096
rect 13587 31093 13599 31127
rect 13541 31087 13599 31093
rect 18322 31084 18328 31136
rect 18380 31124 18386 31136
rect 21177 31127 21235 31133
rect 21177 31124 21189 31127
rect 18380 31096 21189 31124
rect 18380 31084 18386 31096
rect 21177 31093 21189 31096
rect 21223 31124 21235 31127
rect 22388 31124 22416 31300
rect 27525 31297 27537 31331
rect 27571 31328 27583 31331
rect 28261 31331 28319 31337
rect 27571 31300 28120 31328
rect 27571 31297 27583 31300
rect 27525 31291 27583 31297
rect 26694 31220 26700 31272
rect 26752 31260 26758 31272
rect 27157 31263 27215 31269
rect 27157 31260 27169 31263
rect 26752 31232 27169 31260
rect 26752 31220 26758 31232
rect 27157 31229 27169 31232
rect 27203 31229 27215 31263
rect 27157 31223 27215 31229
rect 28092 31201 28120 31300
rect 28261 31297 28273 31331
rect 28307 31297 28319 31331
rect 28626 31328 28632 31340
rect 28587 31300 28632 31328
rect 28261 31291 28319 31297
rect 28626 31288 28632 31300
rect 28684 31288 28690 31340
rect 28966 31260 28994 31436
rect 32585 31433 32597 31467
rect 32631 31464 32643 31467
rect 33778 31464 33784 31476
rect 32631 31436 33784 31464
rect 32631 31433 32643 31436
rect 32585 31427 32643 31433
rect 33778 31424 33784 31436
rect 33836 31424 33842 31476
rect 37829 31467 37887 31473
rect 37829 31433 37841 31467
rect 37875 31464 37887 31467
rect 38194 31464 38200 31476
rect 37875 31436 38200 31464
rect 37875 31433 37887 31436
rect 37829 31427 37887 31433
rect 38194 31424 38200 31436
rect 38252 31424 38258 31476
rect 48590 31424 48596 31476
rect 48648 31424 48654 31476
rect 48682 31424 48688 31476
rect 48740 31464 48746 31476
rect 48869 31467 48927 31473
rect 48869 31464 48881 31467
rect 48740 31436 48881 31464
rect 48740 31424 48746 31436
rect 48869 31433 48881 31436
rect 48915 31433 48927 31467
rect 49786 31464 49792 31476
rect 49747 31436 49792 31464
rect 48869 31427 48927 31433
rect 49786 31424 49792 31436
rect 49844 31424 49850 31476
rect 32122 31396 32128 31408
rect 32083 31368 32128 31396
rect 32122 31356 32128 31368
rect 32180 31356 32186 31408
rect 29641 31331 29699 31337
rect 29641 31297 29653 31331
rect 29687 31328 29699 31331
rect 29730 31328 29736 31340
rect 29687 31300 29736 31328
rect 29687 31297 29699 31300
rect 29641 31291 29699 31297
rect 29656 31260 29684 31291
rect 29730 31288 29736 31300
rect 29788 31288 29794 31340
rect 33962 31328 33968 31340
rect 31726 31300 33968 31328
rect 28966 31232 29684 31260
rect 30101 31263 30159 31269
rect 30101 31229 30113 31263
rect 30147 31260 30159 31263
rect 31726 31260 31754 31300
rect 33962 31288 33968 31300
rect 34020 31288 34026 31340
rect 37461 31331 37519 31337
rect 37461 31297 37473 31331
rect 37507 31328 37519 31331
rect 37550 31328 37556 31340
rect 37507 31300 37556 31328
rect 37507 31297 37519 31300
rect 37461 31291 37519 31297
rect 37550 31288 37556 31300
rect 37608 31288 37614 31340
rect 40494 31288 40500 31340
rect 40552 31328 40558 31340
rect 40773 31331 40831 31337
rect 40773 31328 40785 31331
rect 40552 31300 40785 31328
rect 40552 31288 40558 31300
rect 40773 31297 40785 31300
rect 40819 31297 40831 31331
rect 40773 31291 40831 31297
rect 45370 31288 45376 31340
rect 45428 31328 45434 31340
rect 45465 31331 45523 31337
rect 45465 31328 45477 31331
rect 45428 31300 45477 31328
rect 45428 31288 45434 31300
rect 45465 31297 45477 31300
rect 45511 31297 45523 31331
rect 45465 31291 45523 31297
rect 45646 31288 45652 31340
rect 45704 31328 45710 31340
rect 45741 31331 45799 31337
rect 45741 31328 45753 31331
rect 45704 31300 45753 31328
rect 45704 31288 45710 31300
rect 45741 31297 45753 31300
rect 45787 31297 45799 31331
rect 45741 31291 45799 31297
rect 48314 31288 48320 31340
rect 48372 31328 48378 31340
rect 48409 31331 48467 31337
rect 48409 31328 48421 31331
rect 48372 31300 48421 31328
rect 48372 31288 48378 31300
rect 48409 31297 48421 31300
rect 48455 31297 48467 31331
rect 48409 31291 48467 31297
rect 48501 31331 48559 31337
rect 48501 31297 48513 31331
rect 48547 31328 48559 31331
rect 48608 31328 48636 31424
rect 52730 31396 52736 31408
rect 51920 31368 52736 31396
rect 51920 31337 51948 31368
rect 52730 31356 52736 31368
rect 52788 31356 52794 31408
rect 54938 31396 54944 31408
rect 54899 31368 54944 31396
rect 54938 31356 54944 31368
rect 54996 31356 55002 31408
rect 49329 31331 49387 31337
rect 49329 31328 49341 31331
rect 48547 31300 48636 31328
rect 48792 31300 49341 31328
rect 48547 31297 48559 31300
rect 48501 31291 48559 31297
rect 48792 31272 48820 31300
rect 49329 31297 49341 31300
rect 49375 31297 49387 31331
rect 49329 31291 49387 31297
rect 51905 31331 51963 31337
rect 51905 31297 51917 31331
rect 51951 31297 51963 31331
rect 51905 31291 51963 31297
rect 52089 31331 52147 31337
rect 52089 31297 52101 31331
rect 52135 31297 52147 31331
rect 52089 31291 52147 31297
rect 52181 31331 52239 31337
rect 52181 31297 52193 31331
rect 52227 31328 52239 31331
rect 52362 31328 52368 31340
rect 52227 31300 52368 31328
rect 52227 31297 52239 31300
rect 52181 31291 52239 31297
rect 37366 31260 37372 31272
rect 30147 31232 31754 31260
rect 37327 31232 37372 31260
rect 30147 31229 30159 31232
rect 30101 31223 30159 31229
rect 37366 31220 37372 31232
rect 37424 31220 37430 31272
rect 40678 31260 40684 31272
rect 40639 31232 40684 31260
rect 40678 31220 40684 31232
rect 40736 31220 40742 31272
rect 41141 31263 41199 31269
rect 41141 31229 41153 31263
rect 41187 31260 41199 31263
rect 41322 31260 41328 31272
rect 41187 31232 41328 31260
rect 41187 31229 41199 31232
rect 41141 31223 41199 31229
rect 41322 31220 41328 31232
rect 41380 31220 41386 31272
rect 44453 31263 44511 31269
rect 44453 31229 44465 31263
rect 44499 31260 44511 31263
rect 45094 31260 45100 31272
rect 44499 31232 45100 31260
rect 44499 31229 44511 31232
rect 44453 31223 44511 31229
rect 45094 31220 45100 31232
rect 45152 31260 45158 31272
rect 45278 31260 45284 31272
rect 45152 31232 45284 31260
rect 45152 31220 45158 31232
rect 45278 31220 45284 31232
rect 45336 31220 45342 31272
rect 48222 31220 48228 31272
rect 48280 31260 48286 31272
rect 48593 31263 48651 31269
rect 48593 31260 48605 31263
rect 48280 31232 48605 31260
rect 48280 31220 48286 31232
rect 48593 31229 48605 31232
rect 48639 31229 48651 31263
rect 48593 31223 48651 31229
rect 48685 31263 48743 31269
rect 48685 31229 48697 31263
rect 48731 31260 48743 31263
rect 48774 31260 48780 31272
rect 48731 31232 48780 31260
rect 48731 31229 48743 31232
rect 48685 31223 48743 31229
rect 48774 31220 48780 31232
rect 48832 31220 48838 31272
rect 52104 31260 52132 31291
rect 52362 31288 52368 31300
rect 52420 31288 52426 31340
rect 55398 31328 55404 31340
rect 55359 31300 55404 31328
rect 55398 31288 55404 31300
rect 55456 31288 55462 31340
rect 52270 31260 52276 31272
rect 52104 31232 52276 31260
rect 52270 31220 52276 31232
rect 52328 31220 52334 31272
rect 55306 31220 55312 31272
rect 55364 31260 55370 31272
rect 55493 31263 55551 31269
rect 55493 31260 55505 31263
rect 55364 31232 55505 31260
rect 55364 31220 55370 31232
rect 55493 31229 55505 31232
rect 55539 31229 55551 31263
rect 55493 31223 55551 31229
rect 28077 31195 28135 31201
rect 28077 31161 28089 31195
rect 28123 31161 28135 31195
rect 28077 31155 28135 31161
rect 32214 31152 32220 31204
rect 32272 31192 32278 31204
rect 32401 31195 32459 31201
rect 32401 31192 32413 31195
rect 32272 31164 32413 31192
rect 32272 31152 32278 31164
rect 32401 31161 32413 31164
rect 32447 31161 32459 31195
rect 44818 31192 44824 31204
rect 44779 31164 44824 31192
rect 32401 31155 32459 31161
rect 44818 31152 44824 31164
rect 44876 31152 44882 31204
rect 44913 31195 44971 31201
rect 44913 31161 44925 31195
rect 44959 31192 44971 31195
rect 45557 31195 45615 31201
rect 45557 31192 45569 31195
rect 44959 31164 45569 31192
rect 44959 31161 44971 31164
rect 44913 31155 44971 31161
rect 45557 31161 45569 31164
rect 45603 31161 45615 31195
rect 45557 31155 45615 31161
rect 45646 31152 45652 31204
rect 45704 31192 45710 31204
rect 45925 31195 45983 31201
rect 45704 31164 45749 31192
rect 45704 31152 45710 31164
rect 45925 31161 45937 31195
rect 45971 31192 45983 31195
rect 49970 31192 49976 31204
rect 45971 31164 49976 31192
rect 45971 31161 45983 31164
rect 45925 31155 45983 31161
rect 49970 31152 49976 31164
rect 50028 31152 50034 31204
rect 50062 31152 50068 31204
rect 50120 31192 50126 31204
rect 52362 31192 52368 31204
rect 50120 31164 52368 31192
rect 50120 31152 50126 31164
rect 52362 31152 52368 31164
rect 52420 31152 52426 31204
rect 28350 31124 28356 31136
rect 21223 31096 22416 31124
rect 28311 31096 28356 31124
rect 21223 31093 21235 31096
rect 21177 31087 21235 31093
rect 28350 31084 28356 31096
rect 28408 31084 28414 31136
rect 29086 31124 29092 31136
rect 29047 31096 29092 31124
rect 29086 31084 29092 31096
rect 29144 31124 29150 31136
rect 29733 31127 29791 31133
rect 29733 31124 29745 31127
rect 29144 31096 29745 31124
rect 29144 31084 29150 31096
rect 29733 31093 29745 31096
rect 29779 31093 29791 31127
rect 29733 31087 29791 31093
rect 48314 31084 48320 31136
rect 48372 31124 48378 31136
rect 49421 31127 49479 31133
rect 49421 31124 49433 31127
rect 48372 31096 49433 31124
rect 48372 31084 48378 31096
rect 49421 31093 49433 31096
rect 49467 31093 49479 31127
rect 49421 31087 49479 31093
rect 51721 31127 51779 31133
rect 51721 31093 51733 31127
rect 51767 31124 51779 31127
rect 51994 31124 52000 31136
rect 51767 31096 52000 31124
rect 51767 31093 51779 31096
rect 51721 31087 51779 31093
rect 51994 31084 52000 31096
rect 52052 31084 52058 31136
rect 1104 31034 58880 31056
rect 1104 30982 4214 31034
rect 4266 30982 4278 31034
rect 4330 30982 4342 31034
rect 4394 30982 4406 31034
rect 4458 30982 4470 31034
rect 4522 30982 34934 31034
rect 34986 30982 34998 31034
rect 35050 30982 35062 31034
rect 35114 30982 35126 31034
rect 35178 30982 35190 31034
rect 35242 30982 58880 31034
rect 1104 30960 58880 30982
rect 10045 30923 10103 30929
rect 10045 30889 10057 30923
rect 10091 30920 10103 30923
rect 10134 30920 10140 30932
rect 10091 30892 10140 30920
rect 10091 30889 10103 30892
rect 10045 30883 10103 30889
rect 10134 30880 10140 30892
rect 10192 30880 10198 30932
rect 12894 30880 12900 30932
rect 12952 30920 12958 30932
rect 12989 30923 13047 30929
rect 12989 30920 13001 30923
rect 12952 30892 13001 30920
rect 12952 30880 12958 30892
rect 12989 30889 13001 30892
rect 13035 30889 13047 30923
rect 12989 30883 13047 30889
rect 19334 30880 19340 30932
rect 19392 30920 19398 30932
rect 19392 30892 19437 30920
rect 19392 30880 19398 30892
rect 22094 30880 22100 30932
rect 22152 30920 22158 30932
rect 22649 30923 22707 30929
rect 22649 30920 22661 30923
rect 22152 30892 22661 30920
rect 22152 30880 22158 30892
rect 22649 30889 22661 30892
rect 22695 30889 22707 30923
rect 27798 30920 27804 30932
rect 27759 30892 27804 30920
rect 22649 30883 22707 30889
rect 27798 30880 27804 30892
rect 27856 30880 27862 30932
rect 37366 30920 37372 30932
rect 37327 30892 37372 30920
rect 37366 30880 37372 30892
rect 37424 30880 37430 30932
rect 45097 30923 45155 30929
rect 45097 30889 45109 30923
rect 45143 30920 45155 30923
rect 45186 30920 45192 30932
rect 45143 30892 45192 30920
rect 45143 30889 45155 30892
rect 45097 30883 45155 30889
rect 45186 30880 45192 30892
rect 45244 30880 45250 30932
rect 45278 30880 45284 30932
rect 45336 30920 45342 30932
rect 45649 30923 45707 30929
rect 45649 30920 45661 30923
rect 45336 30892 45661 30920
rect 45336 30880 45342 30892
rect 45649 30889 45661 30892
rect 45695 30889 45707 30923
rect 55490 30920 55496 30932
rect 55451 30892 55496 30920
rect 45649 30883 45707 30889
rect 55490 30880 55496 30892
rect 55548 30880 55554 30932
rect 10318 30852 10324 30864
rect 10279 30824 10324 30852
rect 10318 30812 10324 30824
rect 10376 30812 10382 30864
rect 13354 30852 13360 30864
rect 10428 30824 13360 30852
rect 10428 30784 10456 30824
rect 13354 30812 13360 30824
rect 13412 30812 13418 30864
rect 16942 30852 16948 30864
rect 14200 30824 16948 30852
rect 10336 30756 10456 30784
rect 7282 30716 7288 30728
rect 7243 30688 7288 30716
rect 7282 30676 7288 30688
rect 7340 30676 7346 30728
rect 9858 30676 9864 30728
rect 9916 30716 9922 30728
rect 10229 30719 10287 30725
rect 10229 30718 10241 30719
rect 10152 30716 10241 30718
rect 9916 30690 10241 30716
rect 9916 30688 10180 30690
rect 9916 30676 9922 30688
rect 10229 30685 10241 30690
rect 10275 30685 10287 30719
rect 10229 30679 10287 30685
rect 7377 30651 7435 30657
rect 7377 30617 7389 30651
rect 7423 30648 7435 30651
rect 10336 30648 10364 30756
rect 10594 30744 10600 30796
rect 10652 30784 10658 30796
rect 12710 30784 12716 30796
rect 10652 30756 12716 30784
rect 10652 30744 10658 30756
rect 12710 30744 12716 30756
rect 12768 30744 12774 30796
rect 13262 30784 13268 30796
rect 12820 30756 13268 30784
rect 10413 30719 10471 30725
rect 10413 30685 10425 30719
rect 10459 30685 10471 30719
rect 10413 30679 10471 30685
rect 10505 30719 10563 30725
rect 10505 30685 10517 30719
rect 10551 30716 10563 30719
rect 12820 30716 12848 30756
rect 13262 30744 13268 30756
rect 13320 30744 13326 30796
rect 12986 30716 12992 30728
rect 10551 30688 12848 30716
rect 12947 30688 12992 30716
rect 10551 30685 10563 30688
rect 10505 30679 10563 30685
rect 7423 30620 10364 30648
rect 7423 30617 7435 30620
rect 7377 30611 7435 30617
rect 10042 30540 10048 30592
rect 10100 30580 10106 30592
rect 10428 30580 10456 30679
rect 12986 30676 12992 30688
rect 13044 30676 13050 30728
rect 13078 30676 13084 30728
rect 13136 30716 13142 30728
rect 14200 30716 14228 30824
rect 16942 30812 16948 30824
rect 17000 30812 17006 30864
rect 18046 30852 18052 30864
rect 18007 30824 18052 30852
rect 18046 30812 18052 30824
rect 18104 30812 18110 30864
rect 22830 30812 22836 30864
rect 22888 30852 22894 30864
rect 30929 30855 30987 30861
rect 22888 30824 30604 30852
rect 22888 30812 22894 30824
rect 18322 30784 18328 30796
rect 18235 30756 18328 30784
rect 18322 30744 18328 30756
rect 18380 30744 18386 30796
rect 26878 30784 26884 30796
rect 26839 30756 26884 30784
rect 26878 30744 26884 30756
rect 26936 30784 26942 30796
rect 30466 30784 30472 30796
rect 26936 30756 28028 30784
rect 30427 30756 30472 30784
rect 26936 30744 26942 30756
rect 14366 30716 14372 30728
rect 13136 30688 14228 30716
rect 14327 30688 14372 30716
rect 13136 30676 13142 30688
rect 14366 30676 14372 30688
rect 14424 30676 14430 30728
rect 14550 30716 14556 30728
rect 14511 30688 14556 30716
rect 14550 30676 14556 30688
rect 14608 30716 14614 30728
rect 15838 30716 15844 30728
rect 14608 30688 15844 30716
rect 14608 30676 14614 30688
rect 15838 30676 15844 30688
rect 15896 30676 15902 30728
rect 17497 30719 17555 30725
rect 17497 30716 17509 30719
rect 15948 30688 17509 30716
rect 11238 30608 11244 30660
rect 11296 30648 11302 30660
rect 15948 30648 15976 30688
rect 17497 30685 17509 30688
rect 17543 30716 17555 30719
rect 18340 30716 18368 30744
rect 17543 30688 18368 30716
rect 18417 30719 18475 30725
rect 17543 30685 17555 30688
rect 17497 30679 17555 30685
rect 18417 30685 18429 30719
rect 18463 30716 18475 30719
rect 19334 30716 19340 30728
rect 18463 30688 19340 30716
rect 18463 30685 18475 30688
rect 18417 30679 18475 30685
rect 19334 30676 19340 30688
rect 19392 30676 19398 30728
rect 19426 30676 19432 30728
rect 19484 30716 19490 30728
rect 22830 30716 22836 30728
rect 19484 30688 22692 30716
rect 22791 30688 22836 30716
rect 19484 30676 19490 30688
rect 11296 30620 15976 30648
rect 16025 30651 16083 30657
rect 11296 30608 11302 30620
rect 16025 30617 16037 30651
rect 16071 30648 16083 30651
rect 19518 30648 19524 30660
rect 16071 30620 19524 30648
rect 16071 30617 16083 30620
rect 16025 30611 16083 30617
rect 19518 30608 19524 30620
rect 19576 30608 19582 30660
rect 22664 30648 22692 30688
rect 22830 30676 22836 30688
rect 22888 30676 22894 30728
rect 23106 30716 23112 30728
rect 23067 30688 23112 30716
rect 23106 30676 23112 30688
rect 23164 30676 23170 30728
rect 26970 30716 26976 30728
rect 26931 30688 26976 30716
rect 26970 30676 26976 30688
rect 27028 30676 27034 30728
rect 28000 30725 28028 30756
rect 30466 30744 30472 30756
rect 30524 30744 30530 30796
rect 30576 30784 30604 30824
rect 30929 30821 30941 30855
rect 30975 30852 30987 30855
rect 32122 30852 32128 30864
rect 30975 30824 32128 30852
rect 30975 30821 30987 30824
rect 30929 30815 30987 30821
rect 32122 30812 32128 30824
rect 32180 30812 32186 30864
rect 48961 30855 49019 30861
rect 48961 30821 48973 30855
rect 49007 30852 49019 30855
rect 51350 30852 51356 30864
rect 49007 30824 51356 30852
rect 49007 30821 49019 30824
rect 48961 30815 49019 30821
rect 51350 30812 51356 30824
rect 51408 30812 51414 30864
rect 31389 30787 31447 30793
rect 31389 30784 31401 30787
rect 30576 30756 31401 30784
rect 27985 30719 28043 30725
rect 27985 30685 27997 30719
rect 28031 30685 28043 30719
rect 27985 30679 28043 30685
rect 28169 30719 28227 30725
rect 28169 30685 28181 30719
rect 28215 30716 28227 30719
rect 28718 30716 28724 30728
rect 28215 30688 28724 30716
rect 28215 30685 28227 30688
rect 28169 30679 28227 30685
rect 28718 30676 28724 30688
rect 28776 30676 28782 30728
rect 30576 30725 30604 30756
rect 31389 30753 31401 30756
rect 31435 30784 31447 30787
rect 45002 30784 45008 30796
rect 31435 30756 31754 30784
rect 44963 30756 45008 30784
rect 31435 30753 31447 30756
rect 31389 30747 31447 30753
rect 30561 30719 30619 30725
rect 30561 30685 30573 30719
rect 30607 30685 30619 30719
rect 31726 30716 31754 30756
rect 45002 30744 45008 30756
rect 45060 30744 45066 30796
rect 55306 30784 55312 30796
rect 55267 30756 55312 30784
rect 55306 30744 55312 30756
rect 55364 30744 55370 30796
rect 34514 30716 34520 30728
rect 31726 30688 34520 30716
rect 30561 30679 30619 30685
rect 34514 30676 34520 30688
rect 34572 30676 34578 30728
rect 37182 30716 37188 30728
rect 37143 30688 37188 30716
rect 37182 30676 37188 30688
rect 37240 30676 37246 30728
rect 37369 30719 37427 30725
rect 37369 30685 37381 30719
rect 37415 30716 37427 30719
rect 37458 30716 37464 30728
rect 37415 30688 37464 30716
rect 37415 30685 37427 30688
rect 37369 30679 37427 30685
rect 37458 30676 37464 30688
rect 37516 30676 37522 30728
rect 44358 30676 44364 30728
rect 44416 30716 44422 30728
rect 45370 30716 45376 30728
rect 44416 30688 45376 30716
rect 44416 30676 44422 30688
rect 45370 30676 45376 30688
rect 45428 30716 45434 30728
rect 45468 30719 45526 30725
rect 45468 30716 45480 30719
rect 45428 30688 45480 30716
rect 45428 30676 45434 30688
rect 45468 30685 45480 30688
rect 45514 30685 45526 30719
rect 48314 30716 48320 30728
rect 48275 30688 48320 30716
rect 45468 30679 45526 30685
rect 48314 30676 48320 30688
rect 48372 30676 48378 30728
rect 48406 30676 48412 30728
rect 48464 30716 48470 30728
rect 48464 30688 48509 30716
rect 48464 30676 48470 30688
rect 48590 30676 48596 30728
rect 48648 30716 48654 30728
rect 48774 30716 48780 30728
rect 48648 30688 48693 30716
rect 48735 30688 48780 30716
rect 48648 30676 48654 30688
rect 48774 30676 48780 30688
rect 48832 30676 48838 30728
rect 49970 30676 49976 30728
rect 50028 30716 50034 30728
rect 50890 30716 50896 30728
rect 50028 30688 50896 30716
rect 50028 30676 50034 30688
rect 50890 30676 50896 30688
rect 50948 30676 50954 30728
rect 52270 30716 52276 30728
rect 52231 30688 52276 30716
rect 52270 30676 52276 30688
rect 52328 30676 52334 30728
rect 52362 30676 52368 30728
rect 52420 30716 52426 30728
rect 52733 30719 52791 30725
rect 52733 30716 52745 30719
rect 52420 30688 52745 30716
rect 52420 30676 52426 30688
rect 52733 30685 52745 30688
rect 52779 30685 52791 30719
rect 55766 30716 55772 30728
rect 55727 30688 55772 30716
rect 52733 30679 52791 30685
rect 55766 30676 55772 30688
rect 55824 30676 55830 30728
rect 29086 30648 29092 30660
rect 22664 30620 29092 30648
rect 29086 30608 29092 30620
rect 29144 30608 29150 30660
rect 44818 30608 44824 30660
rect 44876 30648 44882 30660
rect 48222 30648 48228 30660
rect 44876 30620 48228 30648
rect 44876 30608 44882 30620
rect 48222 30608 48228 30620
rect 48280 30648 48286 30660
rect 48685 30651 48743 30657
rect 48685 30648 48697 30651
rect 48280 30620 48697 30648
rect 48280 30608 48286 30620
rect 48685 30617 48697 30620
rect 48731 30617 48743 30651
rect 48685 30611 48743 30617
rect 51074 30608 51080 30660
rect 51132 30648 51138 30660
rect 51132 30620 51177 30648
rect 51132 30608 51138 30620
rect 52178 30608 52184 30660
rect 52236 30608 52242 30660
rect 10100 30552 10456 30580
rect 10100 30540 10106 30552
rect 12710 30540 12716 30592
rect 12768 30580 12774 30592
rect 13078 30580 13084 30592
rect 12768 30552 13084 30580
rect 12768 30540 12774 30552
rect 13078 30540 13084 30552
rect 13136 30540 13142 30592
rect 13357 30583 13415 30589
rect 13357 30549 13369 30583
rect 13403 30580 13415 30583
rect 13538 30580 13544 30592
rect 13403 30552 13544 30580
rect 13403 30549 13415 30552
rect 13357 30543 13415 30549
rect 13538 30540 13544 30552
rect 13596 30540 13602 30592
rect 17494 30540 17500 30592
rect 17552 30580 17558 30592
rect 19426 30580 19432 30592
rect 17552 30552 19432 30580
rect 17552 30540 17558 30552
rect 19426 30540 19432 30552
rect 19484 30540 19490 30592
rect 19889 30583 19947 30589
rect 19889 30549 19901 30583
rect 19935 30580 19947 30583
rect 19978 30580 19984 30592
rect 19935 30552 19984 30580
rect 19935 30549 19947 30552
rect 19889 30543 19947 30549
rect 19978 30540 19984 30552
rect 20036 30540 20042 30592
rect 22186 30580 22192 30592
rect 22099 30552 22192 30580
rect 22186 30540 22192 30552
rect 22244 30580 22250 30592
rect 23014 30580 23020 30592
rect 22244 30552 23020 30580
rect 22244 30540 22250 30552
rect 23014 30540 23020 30552
rect 23072 30540 23078 30592
rect 24489 30583 24547 30589
rect 24489 30549 24501 30583
rect 24535 30580 24547 30583
rect 24762 30580 24768 30592
rect 24535 30552 24768 30580
rect 24535 30549 24547 30552
rect 24489 30543 24547 30549
rect 24762 30540 24768 30552
rect 24820 30540 24826 30592
rect 27341 30583 27399 30589
rect 27341 30549 27353 30583
rect 27387 30580 27399 30583
rect 27706 30580 27712 30592
rect 27387 30552 27712 30580
rect 27387 30549 27399 30552
rect 27341 30543 27399 30549
rect 27706 30540 27712 30552
rect 27764 30540 27770 30592
rect 28718 30580 28724 30592
rect 28679 30552 28724 30580
rect 28718 30540 28724 30552
rect 28776 30540 28782 30592
rect 45462 30580 45468 30592
rect 45423 30552 45468 30580
rect 45462 30540 45468 30552
rect 45520 30540 45526 30592
rect 51261 30583 51319 30589
rect 51261 30549 51273 30583
rect 51307 30580 51319 30583
rect 51626 30580 51632 30592
rect 51307 30552 51632 30580
rect 51307 30549 51319 30552
rect 51261 30543 51319 30549
rect 51626 30540 51632 30552
rect 51684 30540 51690 30592
rect 55677 30583 55735 30589
rect 55677 30549 55689 30583
rect 55723 30580 55735 30583
rect 56042 30580 56048 30592
rect 55723 30552 56048 30580
rect 55723 30549 55735 30552
rect 55677 30543 55735 30549
rect 56042 30540 56048 30552
rect 56100 30580 56106 30592
rect 56229 30583 56287 30589
rect 56229 30580 56241 30583
rect 56100 30552 56241 30580
rect 56100 30540 56106 30552
rect 56229 30549 56241 30552
rect 56275 30549 56287 30583
rect 56229 30543 56287 30549
rect 1104 30490 58880 30512
rect 1104 30438 19574 30490
rect 19626 30438 19638 30490
rect 19690 30438 19702 30490
rect 19754 30438 19766 30490
rect 19818 30438 19830 30490
rect 19882 30438 50294 30490
rect 50346 30438 50358 30490
rect 50410 30438 50422 30490
rect 50474 30438 50486 30490
rect 50538 30438 50550 30490
rect 50602 30438 58880 30490
rect 1104 30416 58880 30438
rect 10318 30336 10324 30388
rect 10376 30376 10382 30388
rect 10778 30376 10784 30388
rect 10376 30348 10784 30376
rect 10376 30336 10382 30348
rect 10778 30336 10784 30348
rect 10836 30336 10842 30388
rect 10962 30336 10968 30388
rect 11020 30376 11026 30388
rect 11020 30348 22508 30376
rect 11020 30336 11026 30348
rect 7009 30311 7067 30317
rect 7009 30277 7021 30311
rect 7055 30308 7067 30311
rect 9490 30308 9496 30320
rect 7055 30280 9496 30308
rect 7055 30277 7067 30280
rect 7009 30271 7067 30277
rect 9490 30268 9496 30280
rect 9548 30268 9554 30320
rect 9585 30311 9643 30317
rect 9585 30277 9597 30311
rect 9631 30308 9643 30311
rect 10042 30308 10048 30320
rect 9631 30280 10048 30308
rect 9631 30277 9643 30280
rect 9585 30271 9643 30277
rect 10042 30268 10048 30280
rect 10100 30268 10106 30320
rect 13170 30308 13176 30320
rect 13131 30280 13176 30308
rect 13170 30268 13176 30280
rect 13228 30268 13234 30320
rect 16022 30268 16028 30320
rect 16080 30308 16086 30320
rect 16669 30311 16727 30317
rect 16669 30308 16681 30311
rect 16080 30280 16681 30308
rect 16080 30268 16086 30280
rect 16669 30277 16681 30280
rect 16715 30277 16727 30311
rect 19978 30308 19984 30320
rect 19891 30280 19984 30308
rect 16669 30271 16727 30277
rect 5442 30200 5448 30252
rect 5500 30240 5506 30252
rect 6825 30243 6883 30249
rect 6825 30240 6837 30243
rect 5500 30212 6837 30240
rect 5500 30200 5506 30212
rect 6825 30209 6837 30212
rect 6871 30209 6883 30243
rect 6825 30203 6883 30209
rect 6914 30200 6920 30252
rect 6972 30240 6978 30252
rect 7469 30243 7527 30249
rect 7469 30240 7481 30243
rect 6972 30212 7481 30240
rect 6972 30200 6978 30212
rect 7469 30209 7481 30212
rect 7515 30209 7527 30243
rect 7650 30240 7656 30252
rect 7611 30212 7656 30240
rect 7469 30203 7527 30209
rect 7650 30200 7656 30212
rect 7708 30200 7714 30252
rect 9861 30243 9919 30249
rect 9861 30209 9873 30243
rect 9907 30240 9919 30243
rect 10686 30240 10692 30252
rect 9907 30212 10692 30240
rect 9907 30209 9919 30212
rect 9861 30203 9919 30209
rect 10686 30200 10692 30212
rect 10744 30200 10750 30252
rect 12894 30240 12900 30252
rect 12807 30212 12900 30240
rect 12894 30200 12900 30212
rect 12952 30200 12958 30252
rect 12986 30200 12992 30252
rect 13044 30240 13050 30252
rect 15381 30243 15439 30249
rect 13044 30212 13089 30240
rect 13044 30200 13050 30212
rect 15381 30209 15393 30243
rect 15427 30209 15439 30243
rect 15381 30203 15439 30209
rect 9122 30132 9128 30184
rect 9180 30172 9186 30184
rect 9769 30175 9827 30181
rect 9769 30172 9781 30175
rect 9180 30144 9781 30172
rect 9180 30132 9186 30144
rect 9769 30141 9781 30144
rect 9815 30141 9827 30175
rect 9769 30135 9827 30141
rect 9953 30175 10011 30181
rect 9953 30141 9965 30175
rect 9999 30172 10011 30175
rect 12434 30172 12440 30184
rect 9999 30144 12440 30172
rect 9999 30141 10011 30144
rect 9953 30135 10011 30141
rect 12434 30132 12440 30144
rect 12492 30132 12498 30184
rect 12912 30104 12940 30200
rect 13173 30175 13231 30181
rect 13173 30141 13185 30175
rect 13219 30172 13231 30175
rect 13262 30172 13268 30184
rect 13219 30144 13268 30172
rect 13219 30141 13231 30144
rect 13173 30135 13231 30141
rect 13262 30132 13268 30144
rect 13320 30172 13326 30184
rect 14550 30172 14556 30184
rect 13320 30144 14556 30172
rect 13320 30132 13326 30144
rect 14550 30132 14556 30144
rect 14608 30132 14614 30184
rect 13814 30104 13820 30116
rect 12912 30076 13820 30104
rect 13814 30064 13820 30076
rect 13872 30064 13878 30116
rect 15396 30048 15424 30203
rect 15562 30200 15568 30252
rect 15620 30240 15626 30252
rect 15838 30240 15844 30252
rect 15620 30212 15665 30240
rect 15799 30212 15844 30240
rect 15620 30200 15626 30212
rect 15838 30200 15844 30212
rect 15896 30200 15902 30252
rect 15930 30200 15936 30252
rect 15988 30240 15994 30252
rect 16117 30243 16175 30249
rect 16117 30240 16129 30243
rect 15988 30212 16129 30240
rect 15988 30200 15994 30212
rect 16117 30209 16129 30212
rect 16163 30240 16175 30243
rect 16163 30212 16896 30240
rect 16163 30209 16175 30212
rect 16117 30203 16175 30209
rect 15580 30172 15608 30200
rect 16761 30175 16819 30181
rect 16761 30172 16773 30175
rect 15580 30164 15976 30172
rect 16040 30164 16773 30172
rect 15580 30144 16773 30164
rect 15948 30136 16068 30144
rect 16761 30141 16773 30144
rect 16807 30141 16819 30175
rect 16868 30172 16896 30212
rect 16942 30200 16948 30252
rect 17000 30240 17006 30252
rect 17862 30240 17868 30252
rect 17000 30212 17868 30240
rect 17000 30200 17006 30212
rect 17862 30200 17868 30212
rect 17920 30240 17926 30252
rect 19904 30249 19932 30280
rect 19978 30268 19984 30280
rect 20036 30308 20042 30320
rect 22480 30317 22508 30348
rect 22830 30336 22836 30388
rect 22888 30376 22894 30388
rect 23109 30379 23167 30385
rect 23109 30376 23121 30379
rect 22888 30348 23121 30376
rect 22888 30336 22894 30348
rect 23109 30345 23121 30348
rect 23155 30345 23167 30379
rect 23109 30339 23167 30345
rect 24394 30336 24400 30388
rect 24452 30376 24458 30388
rect 24489 30379 24547 30385
rect 24489 30376 24501 30379
rect 24452 30348 24501 30376
rect 24452 30336 24458 30348
rect 24489 30345 24501 30348
rect 24535 30345 24547 30379
rect 24489 30339 24547 30345
rect 26970 30336 26976 30388
rect 27028 30376 27034 30388
rect 27525 30379 27583 30385
rect 27525 30376 27537 30379
rect 27028 30348 27537 30376
rect 27028 30336 27034 30348
rect 27525 30345 27537 30348
rect 27571 30376 27583 30379
rect 28718 30376 28724 30388
rect 27571 30348 28724 30376
rect 27571 30345 27583 30348
rect 27525 30339 27583 30345
rect 28718 30336 28724 30348
rect 28776 30336 28782 30388
rect 40129 30379 40187 30385
rect 40129 30345 40141 30379
rect 40175 30376 40187 30379
rect 40402 30376 40408 30388
rect 40175 30348 40408 30376
rect 40175 30345 40187 30348
rect 40129 30339 40187 30345
rect 40402 30336 40408 30348
rect 40460 30376 40466 30388
rect 40678 30376 40684 30388
rect 40460 30348 40684 30376
rect 40460 30336 40466 30348
rect 40678 30336 40684 30348
rect 40736 30336 40742 30388
rect 44358 30376 44364 30388
rect 44319 30348 44364 30376
rect 44358 30336 44364 30348
rect 44416 30336 44422 30388
rect 44818 30336 44824 30388
rect 44876 30376 44882 30388
rect 45097 30379 45155 30385
rect 45097 30376 45109 30379
rect 44876 30348 45109 30376
rect 44876 30336 44882 30348
rect 45097 30345 45109 30348
rect 45143 30345 45155 30379
rect 45097 30339 45155 30345
rect 48593 30379 48651 30385
rect 48593 30345 48605 30379
rect 48639 30376 48651 30379
rect 48774 30376 48780 30388
rect 48639 30348 48780 30376
rect 48639 30345 48651 30348
rect 48593 30339 48651 30345
rect 48774 30336 48780 30348
rect 48832 30336 48838 30388
rect 55306 30336 55312 30388
rect 55364 30336 55370 30388
rect 55398 30336 55404 30388
rect 55456 30376 55462 30388
rect 55953 30379 56011 30385
rect 55953 30376 55965 30379
rect 55456 30348 55965 30376
rect 55456 30336 55462 30348
rect 55953 30345 55965 30348
rect 55999 30345 56011 30379
rect 55953 30339 56011 30345
rect 22465 30311 22523 30317
rect 20036 30280 22094 30308
rect 20036 30268 20042 30280
rect 18417 30243 18475 30249
rect 18417 30240 18429 30243
rect 17920 30212 18429 30240
rect 17920 30200 17926 30212
rect 18417 30209 18429 30212
rect 18463 30209 18475 30243
rect 18417 30203 18475 30209
rect 19889 30243 19947 30249
rect 19889 30209 19901 30243
rect 19935 30209 19947 30243
rect 19889 30203 19947 30209
rect 20717 30243 20775 30249
rect 20717 30209 20729 30243
rect 20763 30209 20775 30243
rect 20717 30203 20775 30209
rect 18693 30175 18751 30181
rect 18693 30172 18705 30175
rect 16868 30144 18705 30172
rect 16761 30135 16819 30141
rect 18693 30141 18705 30144
rect 18739 30172 18751 30175
rect 19794 30172 19800 30184
rect 18739 30144 19334 30172
rect 19755 30144 19800 30172
rect 18739 30141 18751 30144
rect 18693 30135 18751 30141
rect 16117 30107 16175 30113
rect 16117 30073 16129 30107
rect 16163 30104 16175 30107
rect 18230 30104 18236 30116
rect 16163 30076 18236 30104
rect 16163 30073 16175 30076
rect 16117 30067 16175 30073
rect 18230 30064 18236 30076
rect 18288 30064 18294 30116
rect 19306 30104 19334 30144
rect 19794 30132 19800 30144
rect 19852 30132 19858 30184
rect 20732 30172 20760 30203
rect 19904 30144 20760 30172
rect 22066 30172 22094 30280
rect 22465 30277 22477 30311
rect 22511 30277 22523 30311
rect 30374 30308 30380 30320
rect 22465 30271 22523 30277
rect 24044 30280 30380 30308
rect 22480 30240 22508 30271
rect 22922 30240 22928 30252
rect 22480 30212 22928 30240
rect 22922 30200 22928 30212
rect 22980 30240 22986 30252
rect 23017 30243 23075 30249
rect 23017 30240 23029 30243
rect 22980 30212 23029 30240
rect 22980 30200 22986 30212
rect 23017 30209 23029 30212
rect 23063 30209 23075 30243
rect 23017 30203 23075 30209
rect 23106 30200 23112 30252
rect 23164 30240 23170 30252
rect 23201 30243 23259 30249
rect 23201 30240 23213 30243
rect 23164 30212 23213 30240
rect 23164 30200 23170 30212
rect 23201 30209 23213 30212
rect 23247 30209 23259 30243
rect 23201 30203 23259 30209
rect 24044 30172 24072 30280
rect 30374 30268 30380 30280
rect 30432 30268 30438 30320
rect 33689 30311 33747 30317
rect 33689 30277 33701 30311
rect 33735 30308 33747 30311
rect 34146 30308 34152 30320
rect 33735 30280 34152 30308
rect 33735 30277 33747 30280
rect 33689 30271 33747 30277
rect 34146 30268 34152 30280
rect 34204 30268 34210 30320
rect 37182 30268 37188 30320
rect 37240 30308 37246 30320
rect 40494 30308 40500 30320
rect 37240 30280 40500 30308
rect 37240 30268 37246 30280
rect 24121 30243 24179 30249
rect 24121 30209 24133 30243
rect 24167 30240 24179 30243
rect 24854 30240 24860 30252
rect 24167 30212 24860 30240
rect 24167 30209 24179 30212
rect 24121 30203 24179 30209
rect 24854 30200 24860 30212
rect 24912 30200 24918 30252
rect 32674 30200 32680 30252
rect 32732 30240 32738 30252
rect 32861 30243 32919 30249
rect 32861 30240 32873 30243
rect 32732 30212 32873 30240
rect 32732 30200 32738 30212
rect 32861 30209 32873 30212
rect 32907 30209 32919 30243
rect 32861 30203 32919 30209
rect 34422 30200 34428 30252
rect 34480 30240 34486 30252
rect 35161 30243 35219 30249
rect 35161 30240 35173 30243
rect 34480 30212 35173 30240
rect 34480 30200 34486 30212
rect 35161 30209 35173 30212
rect 35207 30209 35219 30243
rect 35161 30203 35219 30209
rect 35989 30243 36047 30249
rect 35989 30209 36001 30243
rect 36035 30209 36047 30243
rect 37277 30243 37335 30249
rect 37277 30240 37289 30243
rect 35989 30203 36047 30209
rect 36464 30212 37289 30240
rect 22066 30144 24072 30172
rect 24213 30175 24271 30181
rect 19904 30104 19932 30144
rect 24213 30141 24225 30175
rect 24259 30172 24271 30175
rect 24302 30172 24308 30184
rect 24259 30144 24308 30172
rect 24259 30141 24271 30144
rect 24213 30135 24271 30141
rect 24302 30132 24308 30144
rect 24360 30132 24366 30184
rect 32766 30172 32772 30184
rect 32727 30144 32772 30172
rect 32766 30132 32772 30144
rect 32824 30132 32830 30184
rect 32950 30132 32956 30184
rect 33008 30172 33014 30184
rect 35069 30175 35127 30181
rect 35069 30172 35081 30175
rect 33008 30144 35081 30172
rect 33008 30132 33014 30144
rect 35069 30141 35081 30144
rect 35115 30172 35127 30175
rect 36004 30172 36032 30203
rect 36464 30181 36492 30212
rect 37277 30209 37289 30212
rect 37323 30209 37335 30243
rect 37277 30203 37335 30209
rect 37458 30200 37464 30252
rect 37516 30240 37522 30252
rect 37844 30249 37872 30280
rect 40494 30268 40500 30280
rect 40552 30268 40558 30320
rect 42613 30311 42671 30317
rect 42613 30277 42625 30311
rect 42659 30308 42671 30311
rect 43070 30308 43076 30320
rect 42659 30280 43076 30308
rect 42659 30277 42671 30280
rect 42613 30271 42671 30277
rect 43070 30268 43076 30280
rect 43128 30268 43134 30320
rect 55125 30311 55183 30317
rect 55125 30277 55137 30311
rect 55171 30308 55183 30311
rect 55324 30308 55352 30336
rect 55171 30280 55352 30308
rect 55692 30280 56180 30308
rect 55171 30277 55183 30280
rect 55125 30271 55183 30277
rect 55692 30252 55720 30280
rect 37553 30243 37611 30249
rect 37553 30240 37565 30243
rect 37516 30212 37565 30240
rect 37516 30200 37522 30212
rect 37553 30209 37565 30212
rect 37599 30209 37611 30243
rect 37553 30203 37611 30209
rect 37829 30243 37887 30249
rect 37829 30209 37841 30243
rect 37875 30209 37887 30243
rect 37829 30203 37887 30209
rect 37921 30243 37979 30249
rect 37921 30209 37933 30243
rect 37967 30209 37979 30243
rect 37921 30203 37979 30209
rect 39761 30243 39819 30249
rect 39761 30209 39773 30243
rect 39807 30209 39819 30243
rect 42426 30240 42432 30252
rect 42387 30212 42432 30240
rect 39761 30203 39819 30209
rect 35115 30144 36032 30172
rect 36449 30175 36507 30181
rect 35115 30141 35127 30144
rect 35069 30135 35127 30141
rect 36449 30141 36461 30175
rect 36495 30141 36507 30175
rect 37936 30172 37964 30203
rect 39666 30172 39672 30184
rect 36449 30135 36507 30141
rect 37568 30144 37964 30172
rect 39627 30144 39672 30172
rect 37568 30116 37596 30144
rect 39666 30132 39672 30144
rect 39724 30132 39730 30184
rect 19306 30076 19932 30104
rect 20257 30107 20315 30113
rect 20257 30073 20269 30107
rect 20303 30104 20315 30107
rect 20990 30104 20996 30116
rect 20303 30076 20996 30104
rect 20303 30073 20315 30076
rect 20257 30067 20315 30073
rect 20990 30064 20996 30076
rect 21048 30064 21054 30116
rect 27062 30064 27068 30116
rect 27120 30104 27126 30116
rect 30377 30107 30435 30113
rect 30377 30104 30389 30107
rect 27120 30076 30389 30104
rect 27120 30064 27126 30076
rect 30377 30073 30389 30076
rect 30423 30104 30435 30107
rect 30926 30104 30932 30116
rect 30423 30076 30932 30104
rect 30423 30073 30435 30076
rect 30377 30067 30435 30073
rect 30926 30064 30932 30076
rect 30984 30064 30990 30116
rect 35529 30107 35587 30113
rect 35529 30073 35541 30107
rect 35575 30104 35587 30107
rect 37550 30104 37556 30116
rect 35575 30076 37556 30104
rect 35575 30073 35587 30076
rect 35529 30067 35587 30073
rect 37550 30064 37556 30076
rect 37608 30064 37614 30116
rect 37645 30107 37703 30113
rect 37645 30073 37657 30107
rect 37691 30104 37703 30107
rect 39776 30104 39804 30203
rect 42426 30200 42432 30212
rect 42484 30200 42490 30252
rect 42705 30243 42763 30249
rect 42705 30209 42717 30243
rect 42751 30209 42763 30243
rect 42705 30203 42763 30209
rect 43165 30243 43223 30249
rect 43165 30209 43177 30243
rect 43211 30209 43223 30243
rect 43165 30203 43223 30209
rect 43349 30243 43407 30249
rect 43349 30209 43361 30243
rect 43395 30240 43407 30243
rect 44266 30240 44272 30252
rect 43395 30212 44272 30240
rect 43395 30209 43407 30212
rect 43349 30203 43407 30209
rect 39850 30132 39856 30184
rect 39908 30172 39914 30184
rect 41049 30175 41107 30181
rect 41049 30172 41061 30175
rect 39908 30144 41061 30172
rect 39908 30132 39914 30144
rect 41049 30141 41061 30144
rect 41095 30141 41107 30175
rect 41049 30135 41107 30141
rect 42518 30132 42524 30184
rect 42576 30172 42582 30184
rect 42720 30172 42748 30203
rect 42576 30144 42748 30172
rect 42576 30132 42582 30144
rect 40681 30107 40739 30113
rect 40681 30104 40693 30107
rect 37691 30076 40693 30104
rect 37691 30073 37703 30076
rect 37645 30067 37703 30073
rect 40681 30073 40693 30076
rect 40727 30073 40739 30107
rect 40681 30067 40739 30073
rect 42429 30107 42487 30113
rect 42429 30073 42441 30107
rect 42475 30104 42487 30107
rect 43180 30104 43208 30203
rect 44266 30200 44272 30212
rect 44324 30200 44330 30252
rect 44453 30243 44511 30249
rect 44453 30209 44465 30243
rect 44499 30240 44511 30243
rect 44913 30243 44971 30249
rect 44913 30240 44925 30243
rect 44499 30212 44925 30240
rect 44499 30209 44511 30212
rect 44453 30203 44511 30209
rect 44913 30209 44925 30212
rect 44959 30240 44971 30243
rect 45002 30240 45008 30252
rect 44959 30212 45008 30240
rect 44959 30209 44971 30212
rect 44913 30203 44971 30209
rect 45002 30200 45008 30212
rect 45060 30200 45066 30252
rect 45094 30200 45100 30252
rect 45152 30240 45158 30252
rect 45281 30243 45339 30249
rect 45281 30240 45293 30243
rect 45152 30212 45293 30240
rect 45152 30200 45158 30212
rect 45281 30209 45293 30212
rect 45327 30209 45339 30243
rect 45281 30203 45339 30209
rect 48038 30200 48044 30252
rect 48096 30240 48102 30252
rect 48133 30243 48191 30249
rect 48133 30240 48145 30243
rect 48096 30212 48145 30240
rect 48096 30200 48102 30212
rect 48133 30209 48145 30212
rect 48179 30209 48191 30243
rect 48133 30203 48191 30209
rect 51261 30243 51319 30249
rect 51261 30209 51273 30243
rect 51307 30209 51319 30243
rect 51626 30240 51632 30252
rect 51587 30212 51632 30240
rect 51261 30203 51319 30209
rect 42475 30076 43208 30104
rect 43533 30107 43591 30113
rect 42475 30073 42487 30076
rect 42429 30067 42487 30073
rect 43533 30073 43545 30107
rect 43579 30104 43591 30107
rect 43579 30076 45232 30104
rect 43579 30073 43591 30076
rect 43533 30067 43591 30073
rect 45204 30048 45232 30076
rect 49510 30064 49516 30116
rect 49568 30104 49574 30116
rect 51169 30107 51227 30113
rect 51169 30104 51181 30107
rect 49568 30076 51181 30104
rect 49568 30064 49574 30076
rect 51169 30073 51181 30076
rect 51215 30073 51227 30107
rect 51276 30104 51304 30203
rect 51626 30200 51632 30212
rect 51684 30240 51690 30252
rect 52733 30243 52791 30249
rect 52733 30240 52745 30243
rect 51684 30212 52745 30240
rect 51684 30200 51690 30212
rect 52733 30209 52745 30212
rect 52779 30209 52791 30243
rect 55306 30240 55312 30252
rect 55267 30212 55312 30240
rect 52733 30203 52791 30209
rect 55306 30200 55312 30212
rect 55364 30200 55370 30252
rect 55493 30243 55551 30249
rect 55493 30209 55505 30243
rect 55539 30240 55551 30243
rect 55674 30240 55680 30252
rect 55539 30212 55680 30240
rect 55539 30209 55551 30212
rect 55493 30203 55551 30209
rect 55674 30200 55680 30212
rect 55732 30200 55738 30252
rect 56152 30249 56180 30280
rect 55953 30243 56011 30249
rect 55953 30209 55965 30243
rect 55999 30209 56011 30243
rect 55953 30203 56011 30209
rect 56137 30243 56195 30249
rect 56137 30209 56149 30243
rect 56183 30209 56195 30243
rect 56137 30203 56195 30209
rect 52086 30172 52092 30184
rect 52047 30144 52092 30172
rect 52086 30132 52092 30144
rect 52144 30132 52150 30184
rect 55324 30172 55352 30200
rect 55968 30172 55996 30203
rect 55324 30144 55996 30172
rect 51718 30104 51724 30116
rect 51276 30076 51724 30104
rect 51169 30067 51227 30073
rect 51718 30064 51724 30076
rect 51776 30104 51782 30116
rect 51776 30076 52868 30104
rect 51776 30064 51782 30076
rect 7653 30039 7711 30045
rect 7653 30005 7665 30039
rect 7699 30036 7711 30039
rect 10502 30036 10508 30048
rect 7699 30008 10508 30036
rect 7699 30005 7711 30008
rect 7653 29999 7711 30005
rect 10502 29996 10508 30008
rect 10560 29996 10566 30048
rect 10597 30039 10655 30045
rect 10597 30005 10609 30039
rect 10643 30036 10655 30039
rect 11054 30036 11060 30048
rect 10643 30008 11060 30036
rect 10643 30005 10655 30008
rect 10597 29999 10655 30005
rect 11054 29996 11060 30008
rect 11112 29996 11118 30048
rect 15378 30036 15384 30048
rect 15291 30008 15384 30036
rect 15378 29996 15384 30008
rect 15436 30036 15442 30048
rect 16669 30039 16727 30045
rect 16669 30036 16681 30039
rect 15436 30008 16681 30036
rect 15436 29996 15442 30008
rect 16669 30005 16681 30008
rect 16715 30005 16727 30039
rect 16669 29999 16727 30005
rect 17129 30039 17187 30045
rect 17129 30005 17141 30039
rect 17175 30036 17187 30039
rect 18414 30036 18420 30048
rect 17175 30008 18420 30036
rect 17175 30005 17187 30008
rect 17129 29999 17187 30005
rect 18414 29996 18420 30008
rect 18472 29996 18478 30048
rect 20901 30039 20959 30045
rect 20901 30005 20913 30039
rect 20947 30036 20959 30039
rect 22186 30036 22192 30048
rect 20947 30008 22192 30036
rect 20947 30005 20959 30008
rect 20901 29999 20959 30005
rect 22186 29996 22192 30008
rect 22244 29996 22250 30048
rect 22922 29996 22928 30048
rect 22980 30036 22986 30048
rect 24121 30039 24179 30045
rect 24121 30036 24133 30039
rect 22980 30008 24133 30036
rect 22980 29996 22986 30008
rect 24121 30005 24133 30008
rect 24167 30036 24179 30039
rect 24762 30036 24768 30048
rect 24167 30008 24768 30036
rect 24167 30005 24179 30008
rect 24121 29999 24179 30005
rect 24762 29996 24768 30008
rect 24820 30036 24826 30048
rect 24949 30039 25007 30045
rect 24949 30036 24961 30039
rect 24820 30008 24961 30036
rect 24820 29996 24826 30008
rect 24949 30005 24961 30008
rect 24995 30005 25007 30039
rect 24949 29999 25007 30005
rect 34422 29996 34428 30048
rect 34480 30036 34486 30048
rect 36081 30039 36139 30045
rect 36081 30036 36093 30039
rect 34480 30008 36093 30036
rect 34480 29996 34486 30008
rect 36081 30005 36093 30008
rect 36127 30005 36139 30039
rect 40586 30036 40592 30048
rect 40547 30008 40592 30036
rect 36081 29999 36139 30005
rect 40586 29996 40592 30008
rect 40644 29996 40650 30048
rect 45186 29996 45192 30048
rect 45244 30036 45250 30048
rect 45281 30039 45339 30045
rect 45281 30036 45293 30039
rect 45244 30008 45293 30036
rect 45244 29996 45250 30008
rect 45281 30005 45293 30008
rect 45327 30005 45339 30039
rect 45281 29999 45339 30005
rect 45370 29996 45376 30048
rect 45428 30036 45434 30048
rect 48317 30039 48375 30045
rect 48317 30036 48329 30039
rect 45428 30008 48329 30036
rect 45428 29996 45434 30008
rect 48317 30005 48329 30008
rect 48363 30036 48375 30039
rect 48498 30036 48504 30048
rect 48363 30008 48504 30036
rect 48363 30005 48375 30008
rect 48317 29999 48375 30005
rect 48498 29996 48504 30008
rect 48556 29996 48562 30048
rect 52840 30045 52868 30076
rect 52825 30039 52883 30045
rect 52825 30005 52837 30039
rect 52871 30005 52883 30039
rect 52825 29999 52883 30005
rect 53006 29996 53012 30048
rect 53064 30036 53070 30048
rect 53193 30039 53251 30045
rect 53193 30036 53205 30039
rect 53064 30008 53205 30036
rect 53064 29996 53070 30008
rect 53193 30005 53205 30008
rect 53239 30005 53251 30039
rect 53193 29999 53251 30005
rect 56042 29996 56048 30048
rect 56100 30036 56106 30048
rect 57057 30039 57115 30045
rect 57057 30036 57069 30039
rect 56100 30008 57069 30036
rect 56100 29996 56106 30008
rect 57057 30005 57069 30008
rect 57103 30005 57115 30039
rect 57057 29999 57115 30005
rect 1104 29946 58880 29968
rect 1104 29894 4214 29946
rect 4266 29894 4278 29946
rect 4330 29894 4342 29946
rect 4394 29894 4406 29946
rect 4458 29894 4470 29946
rect 4522 29894 34934 29946
rect 34986 29894 34998 29946
rect 35050 29894 35062 29946
rect 35114 29894 35126 29946
rect 35178 29894 35190 29946
rect 35242 29894 58880 29946
rect 1104 29872 58880 29894
rect 2222 29832 2228 29844
rect 2183 29804 2228 29832
rect 2222 29792 2228 29804
rect 2280 29792 2286 29844
rect 7374 29792 7380 29844
rect 7432 29832 7438 29844
rect 9674 29832 9680 29844
rect 7432 29804 9680 29832
rect 7432 29792 7438 29804
rect 9674 29792 9680 29804
rect 9732 29792 9738 29844
rect 9858 29832 9864 29844
rect 9819 29804 9864 29832
rect 9858 29792 9864 29804
rect 9916 29792 9922 29844
rect 10686 29832 10692 29844
rect 10647 29804 10692 29832
rect 10686 29792 10692 29804
rect 10744 29792 10750 29844
rect 10778 29792 10784 29844
rect 10836 29832 10842 29844
rect 10873 29835 10931 29841
rect 10873 29832 10885 29835
rect 10836 29804 10885 29832
rect 10836 29792 10842 29804
rect 10873 29801 10885 29804
rect 10919 29801 10931 29835
rect 12986 29832 12992 29844
rect 12947 29804 12992 29832
rect 10873 29795 10931 29801
rect 12986 29792 12992 29804
rect 13044 29792 13050 29844
rect 14458 29832 14464 29844
rect 14419 29804 14464 29832
rect 14458 29792 14464 29804
rect 14516 29832 14522 29844
rect 15102 29832 15108 29844
rect 14516 29804 15108 29832
rect 14516 29792 14522 29804
rect 15102 29792 15108 29804
rect 15160 29792 15166 29844
rect 15378 29832 15384 29844
rect 15339 29804 15384 29832
rect 15378 29792 15384 29804
rect 15436 29792 15442 29844
rect 15838 29832 15844 29844
rect 15799 29804 15844 29832
rect 15838 29792 15844 29804
rect 15896 29792 15902 29844
rect 19337 29835 19395 29841
rect 19337 29801 19349 29835
rect 19383 29832 19395 29835
rect 19978 29832 19984 29844
rect 19383 29804 19984 29832
rect 19383 29801 19395 29804
rect 19337 29795 19395 29801
rect 19978 29792 19984 29804
rect 20036 29792 20042 29844
rect 22922 29832 22928 29844
rect 22883 29804 22928 29832
rect 22922 29792 22928 29804
rect 22980 29792 22986 29844
rect 23014 29792 23020 29844
rect 23072 29832 23078 29844
rect 27525 29835 27583 29841
rect 23072 29804 25544 29832
rect 23072 29792 23078 29804
rect 9309 29767 9367 29773
rect 9309 29733 9321 29767
rect 9355 29764 9367 29767
rect 11054 29764 11060 29776
rect 9355 29736 11060 29764
rect 9355 29733 9367 29736
rect 9309 29727 9367 29733
rect 11054 29724 11060 29736
rect 11112 29724 11118 29776
rect 15120 29764 15148 29792
rect 19058 29764 19064 29776
rect 15120 29736 19064 29764
rect 19058 29724 19064 29736
rect 19116 29724 19122 29776
rect 19150 29724 19156 29776
rect 19208 29764 19214 29776
rect 19889 29767 19947 29773
rect 19889 29764 19901 29767
rect 19208 29736 19901 29764
rect 19208 29724 19214 29736
rect 19889 29733 19901 29736
rect 19935 29733 19947 29767
rect 19889 29727 19947 29733
rect 23661 29767 23719 29773
rect 23661 29733 23673 29767
rect 23707 29733 23719 29767
rect 23661 29727 23719 29733
rect 23753 29767 23811 29773
rect 23753 29733 23765 29767
rect 23799 29764 23811 29767
rect 24854 29764 24860 29776
rect 23799 29736 24860 29764
rect 23799 29733 23811 29736
rect 23753 29727 23811 29733
rect 3326 29656 3332 29708
rect 3384 29696 3390 29708
rect 3881 29699 3939 29705
rect 3881 29696 3893 29699
rect 3384 29668 3893 29696
rect 3384 29656 3390 29668
rect 3881 29665 3893 29668
rect 3927 29665 3939 29699
rect 5718 29696 5724 29708
rect 5679 29668 5724 29696
rect 3881 29659 3939 29665
rect 5718 29656 5724 29668
rect 5776 29656 5782 29708
rect 5997 29699 6055 29705
rect 5997 29665 6009 29699
rect 6043 29696 6055 29699
rect 7650 29696 7656 29708
rect 6043 29668 7656 29696
rect 6043 29665 6055 29668
rect 5997 29659 6055 29665
rect 7650 29656 7656 29668
rect 7708 29656 7714 29708
rect 19426 29696 19432 29708
rect 12452 29668 19432 29696
rect 12452 29640 12480 29668
rect 19426 29656 19432 29668
rect 19484 29696 19490 29708
rect 21637 29699 21695 29705
rect 21637 29696 21649 29699
rect 19484 29668 21649 29696
rect 19484 29656 19490 29668
rect 21637 29665 21649 29668
rect 21683 29696 21695 29699
rect 21683 29668 22094 29696
rect 21683 29665 21695 29668
rect 21637 29659 21695 29665
rect 1673 29631 1731 29637
rect 1673 29597 1685 29631
rect 1719 29628 1731 29631
rect 2222 29628 2228 29640
rect 1719 29600 2228 29628
rect 1719 29597 1731 29600
rect 1673 29591 1731 29597
rect 2222 29588 2228 29600
rect 2280 29588 2286 29640
rect 3973 29631 4031 29637
rect 3973 29597 3985 29631
rect 4019 29628 4031 29631
rect 4019 29600 4936 29628
rect 4019 29597 4031 29600
rect 3973 29591 4031 29597
rect 4908 29504 4936 29600
rect 5442 29588 5448 29640
rect 5500 29628 5506 29640
rect 5629 29631 5687 29637
rect 5629 29628 5641 29631
rect 5500 29600 5641 29628
rect 5500 29588 5506 29600
rect 5629 29597 5641 29600
rect 5675 29597 5687 29631
rect 7374 29628 7380 29640
rect 7335 29600 7380 29628
rect 5629 29591 5687 29597
rect 7374 29588 7380 29600
rect 7432 29588 7438 29640
rect 9674 29588 9680 29640
rect 9732 29628 9738 29640
rect 10321 29631 10379 29637
rect 10321 29628 10333 29631
rect 9732 29600 10333 29628
rect 9732 29588 9738 29600
rect 10321 29597 10333 29600
rect 10367 29597 10379 29631
rect 10321 29591 10379 29597
rect 12434 29588 12440 29640
rect 12492 29628 12498 29640
rect 12805 29631 12863 29637
rect 12492 29600 12537 29628
rect 12492 29588 12498 29600
rect 12805 29597 12817 29631
rect 12851 29628 12863 29631
rect 13630 29628 13636 29640
rect 12851 29600 13636 29628
rect 12851 29597 12863 29600
rect 12805 29591 12863 29597
rect 13630 29588 13636 29600
rect 13688 29588 13694 29640
rect 15010 29628 15016 29640
rect 14971 29600 15016 29628
rect 15010 29588 15016 29600
rect 15068 29588 15074 29640
rect 15102 29588 15108 29640
rect 15160 29628 15166 29640
rect 15197 29631 15255 29637
rect 15197 29628 15209 29631
rect 15160 29600 15209 29628
rect 15160 29588 15166 29600
rect 15197 29597 15209 29600
rect 15243 29597 15255 29631
rect 16022 29628 16028 29640
rect 15983 29600 16028 29628
rect 15197 29591 15255 29597
rect 16022 29588 16028 29600
rect 16080 29588 16086 29640
rect 16206 29628 16212 29640
rect 16167 29600 16212 29628
rect 16206 29588 16212 29600
rect 16264 29588 16270 29640
rect 17862 29588 17868 29640
rect 17920 29628 17926 29640
rect 19245 29631 19303 29637
rect 19245 29628 19257 29631
rect 17920 29600 19257 29628
rect 17920 29588 17926 29600
rect 19245 29597 19257 29600
rect 19291 29597 19303 29631
rect 19245 29591 19303 29597
rect 7466 29520 7472 29572
rect 7524 29560 7530 29572
rect 12618 29560 12624 29572
rect 7524 29532 12624 29560
rect 7524 29520 7530 29532
rect 12618 29520 12624 29532
rect 12676 29520 12682 29572
rect 12713 29563 12771 29569
rect 12713 29529 12725 29563
rect 12759 29529 12771 29563
rect 12713 29523 12771 29529
rect 1486 29492 1492 29504
rect 1447 29464 1492 29492
rect 1486 29452 1492 29464
rect 1544 29452 1550 29504
rect 4338 29492 4344 29504
rect 4299 29464 4344 29492
rect 4338 29452 4344 29464
rect 4396 29452 4402 29504
rect 4890 29492 4896 29504
rect 4851 29464 4896 29492
rect 4890 29452 4896 29464
rect 4948 29452 4954 29504
rect 9677 29495 9735 29501
rect 9677 29461 9689 29495
rect 9723 29492 9735 29495
rect 9858 29492 9864 29504
rect 9723 29464 9864 29492
rect 9723 29461 9735 29464
rect 9677 29455 9735 29461
rect 9858 29452 9864 29464
rect 9916 29452 9922 29504
rect 10689 29495 10747 29501
rect 10689 29461 10701 29495
rect 10735 29492 10747 29495
rect 12250 29492 12256 29504
rect 10735 29464 12256 29492
rect 10735 29461 10747 29464
rect 10689 29455 10747 29461
rect 12250 29452 12256 29464
rect 12308 29452 12314 29504
rect 12342 29452 12348 29504
rect 12400 29492 12406 29504
rect 12728 29492 12756 29523
rect 14182 29520 14188 29572
rect 14240 29560 14246 29572
rect 19794 29560 19800 29572
rect 14240 29532 19800 29560
rect 14240 29520 14246 29532
rect 19794 29520 19800 29532
rect 19852 29520 19858 29572
rect 21453 29563 21511 29569
rect 21453 29529 21465 29563
rect 21499 29529 21511 29563
rect 22066 29560 22094 29668
rect 23106 29656 23112 29708
rect 23164 29696 23170 29708
rect 23569 29699 23627 29705
rect 23569 29696 23581 29699
rect 23164 29668 23581 29696
rect 23164 29656 23170 29668
rect 23569 29665 23581 29668
rect 23615 29665 23627 29699
rect 23676 29696 23704 29727
rect 24854 29724 24860 29736
rect 24912 29764 24918 29776
rect 25406 29764 25412 29776
rect 24912 29736 25412 29764
rect 24912 29724 24918 29736
rect 25406 29724 25412 29736
rect 25464 29724 25470 29776
rect 25516 29764 25544 29804
rect 27525 29801 27537 29835
rect 27571 29832 27583 29835
rect 27798 29832 27804 29844
rect 27571 29804 27804 29832
rect 27571 29801 27583 29804
rect 27525 29795 27583 29801
rect 27798 29792 27804 29804
rect 27856 29832 27862 29844
rect 28350 29832 28356 29844
rect 27856 29804 28356 29832
rect 27856 29792 27862 29804
rect 28350 29792 28356 29804
rect 28408 29792 28414 29844
rect 30285 29835 30343 29841
rect 30285 29801 30297 29835
rect 30331 29832 30343 29835
rect 30374 29832 30380 29844
rect 30331 29804 30380 29832
rect 30331 29801 30343 29804
rect 30285 29795 30343 29801
rect 30374 29792 30380 29804
rect 30432 29792 30438 29844
rect 32950 29832 32956 29844
rect 32911 29804 32956 29832
rect 32950 29792 32956 29804
rect 33008 29792 33014 29844
rect 36817 29835 36875 29841
rect 36817 29801 36829 29835
rect 36863 29832 36875 29835
rect 37182 29832 37188 29844
rect 36863 29804 37188 29832
rect 36863 29801 36875 29804
rect 36817 29795 36875 29801
rect 37182 29792 37188 29804
rect 37240 29792 37246 29844
rect 37458 29832 37464 29844
rect 37419 29804 37464 29832
rect 37458 29792 37464 29804
rect 37516 29792 37522 29844
rect 42518 29792 42524 29844
rect 42576 29832 42582 29844
rect 42797 29835 42855 29841
rect 42797 29832 42809 29835
rect 42576 29804 42809 29832
rect 42576 29792 42582 29804
rect 42797 29801 42809 29804
rect 42843 29801 42855 29835
rect 42797 29795 42855 29801
rect 45373 29835 45431 29841
rect 45373 29801 45385 29835
rect 45419 29832 45431 29835
rect 45462 29832 45468 29844
rect 45419 29804 45468 29832
rect 45419 29801 45431 29804
rect 45373 29795 45431 29801
rect 45462 29792 45468 29804
rect 45520 29792 45526 29844
rect 48314 29832 48320 29844
rect 48275 29804 48320 29832
rect 48314 29792 48320 29804
rect 48372 29792 48378 29844
rect 30834 29764 30840 29776
rect 25516 29736 30840 29764
rect 30834 29724 30840 29736
rect 30892 29724 30898 29776
rect 42981 29767 43039 29773
rect 42981 29733 42993 29767
rect 43027 29764 43039 29767
rect 47857 29767 47915 29773
rect 43027 29736 44312 29764
rect 43027 29733 43039 29736
rect 42981 29727 43039 29733
rect 44284 29708 44312 29736
rect 47857 29733 47869 29767
rect 47903 29764 47915 29767
rect 48685 29767 48743 29773
rect 48685 29764 48697 29767
rect 47903 29736 48697 29764
rect 47903 29733 47915 29736
rect 47857 29727 47915 29733
rect 48685 29733 48697 29736
rect 48731 29733 48743 29767
rect 48685 29727 48743 29733
rect 30926 29696 30932 29708
rect 23676 29668 24624 29696
rect 30887 29668 30932 29696
rect 23569 29659 23627 29665
rect 22922 29588 22928 29640
rect 22980 29628 22986 29640
rect 23477 29631 23535 29637
rect 23477 29628 23489 29631
rect 22980 29600 23489 29628
rect 22980 29588 22986 29600
rect 23477 29597 23489 29600
rect 23523 29597 23535 29631
rect 23477 29591 23535 29597
rect 23584 29560 23612 29659
rect 23842 29628 23848 29640
rect 23803 29600 23848 29628
rect 23842 29588 23848 29600
rect 23900 29588 23906 29640
rect 24394 29628 24400 29640
rect 24355 29600 24400 29628
rect 24394 29588 24400 29600
rect 24452 29588 24458 29640
rect 24596 29637 24624 29668
rect 30926 29656 30932 29668
rect 30984 29656 30990 29708
rect 32674 29696 32680 29708
rect 32635 29668 32680 29696
rect 32674 29656 32680 29668
rect 32732 29656 32738 29708
rect 32766 29656 32772 29708
rect 32824 29696 32830 29708
rect 32824 29668 32869 29696
rect 36648 29668 37504 29696
rect 32824 29656 32830 29668
rect 24581 29631 24639 29637
rect 24581 29597 24593 29631
rect 24627 29597 24639 29631
rect 24581 29591 24639 29597
rect 24673 29631 24731 29637
rect 24673 29597 24685 29631
rect 24719 29597 24731 29631
rect 24673 29591 24731 29597
rect 24688 29560 24716 29591
rect 24762 29588 24768 29640
rect 24820 29628 24826 29640
rect 27706 29628 27712 29640
rect 24820 29600 24865 29628
rect 27667 29600 27712 29628
rect 24820 29588 24826 29600
rect 27706 29588 27712 29600
rect 27764 29588 27770 29640
rect 27890 29588 27896 29640
rect 27948 29628 27954 29640
rect 27985 29631 28043 29637
rect 27985 29628 27997 29631
rect 27948 29600 27997 29628
rect 27948 29588 27954 29600
rect 27985 29597 27997 29600
rect 28031 29597 28043 29631
rect 27985 29591 28043 29597
rect 28074 29588 28080 29640
rect 28132 29628 28138 29640
rect 28169 29631 28227 29637
rect 28169 29628 28181 29631
rect 28132 29600 28181 29628
rect 28132 29588 28138 29600
rect 28169 29597 28181 29600
rect 28215 29597 28227 29631
rect 28169 29591 28227 29597
rect 30374 29588 30380 29640
rect 30432 29628 30438 29640
rect 30650 29628 30656 29640
rect 30432 29600 30656 29628
rect 30432 29588 30438 29600
rect 30650 29588 30656 29600
rect 30708 29628 30714 29640
rect 31021 29631 31079 29637
rect 31021 29628 31033 29631
rect 30708 29600 31033 29628
rect 30708 29588 30714 29600
rect 31021 29597 31033 29600
rect 31067 29597 31079 29631
rect 31021 29591 31079 29597
rect 31849 29631 31907 29637
rect 31849 29597 31861 29631
rect 31895 29628 31907 29631
rect 32784 29628 32812 29656
rect 36648 29640 36676 29668
rect 36446 29628 36452 29640
rect 31895 29600 32812 29628
rect 36407 29600 36452 29628
rect 31895 29597 31907 29600
rect 31849 29591 31907 29597
rect 36446 29588 36452 29600
rect 36504 29588 36510 29640
rect 36630 29628 36636 29640
rect 36591 29600 36636 29628
rect 36630 29588 36636 29600
rect 36688 29588 36694 29640
rect 37476 29637 37504 29668
rect 44266 29656 44272 29708
rect 44324 29696 44330 29708
rect 44324 29668 45232 29696
rect 44324 29656 44330 29668
rect 37277 29631 37335 29637
rect 37277 29597 37289 29631
rect 37323 29597 37335 29631
rect 37277 29591 37335 29597
rect 37461 29631 37519 29637
rect 37461 29597 37473 29631
rect 37507 29597 37519 29631
rect 40402 29628 40408 29640
rect 40363 29600 40408 29628
rect 37461 29591 37519 29597
rect 22066 29532 23520 29560
rect 23584 29532 24716 29560
rect 21453 29523 21511 29529
rect 13722 29492 13728 29504
rect 12400 29464 13728 29492
rect 12400 29452 12406 29464
rect 13722 29452 13728 29464
rect 13780 29452 13786 29504
rect 14090 29452 14096 29504
rect 14148 29492 14154 29504
rect 15470 29492 15476 29504
rect 14148 29464 15476 29492
rect 14148 29452 14154 29464
rect 15470 29452 15476 29464
rect 15528 29452 15534 29504
rect 17586 29452 17592 29504
rect 17644 29492 17650 29504
rect 18601 29495 18659 29501
rect 18601 29492 18613 29495
rect 17644 29464 18613 29492
rect 17644 29452 17650 29464
rect 18601 29461 18613 29464
rect 18647 29492 18659 29495
rect 21468 29492 21496 29523
rect 22189 29495 22247 29501
rect 22189 29492 22201 29495
rect 18647 29464 22201 29492
rect 18647 29461 18659 29464
rect 18601 29455 18659 29461
rect 22189 29461 22201 29464
rect 22235 29492 22247 29495
rect 22370 29492 22376 29504
rect 22235 29464 22376 29492
rect 22235 29461 22247 29464
rect 22189 29455 22247 29461
rect 22370 29452 22376 29464
rect 22428 29452 22434 29504
rect 23492 29492 23520 29532
rect 24118 29492 24124 29504
rect 23492 29464 24124 29492
rect 24118 29452 24124 29464
rect 24176 29452 24182 29504
rect 25041 29495 25099 29501
rect 25041 29461 25053 29495
rect 25087 29492 25099 29495
rect 27154 29492 27160 29504
rect 25087 29464 27160 29492
rect 25087 29461 25099 29464
rect 25041 29455 25099 29461
rect 27154 29452 27160 29464
rect 27212 29452 27218 29504
rect 27724 29492 27752 29588
rect 36464 29560 36492 29588
rect 37292 29560 37320 29591
rect 40402 29588 40408 29600
rect 40460 29588 40466 29640
rect 40586 29588 40592 29640
rect 40644 29628 40650 29640
rect 40681 29631 40739 29637
rect 40681 29628 40693 29631
rect 40644 29600 40693 29628
rect 40644 29588 40650 29600
rect 40681 29597 40693 29600
rect 40727 29597 40739 29631
rect 45002 29628 45008 29640
rect 44963 29600 45008 29628
rect 40681 29591 40739 29597
rect 45002 29588 45008 29600
rect 45060 29588 45066 29640
rect 45204 29637 45232 29668
rect 55214 29656 55220 29708
rect 55272 29696 55278 29708
rect 56045 29699 56103 29705
rect 56045 29696 56057 29699
rect 55272 29668 56057 29696
rect 55272 29656 55278 29668
rect 56045 29665 56057 29668
rect 56091 29665 56103 29699
rect 57333 29699 57391 29705
rect 57333 29696 57345 29699
rect 56045 29659 56103 29665
rect 56796 29668 57345 29696
rect 45189 29631 45247 29637
rect 45189 29597 45201 29631
rect 45235 29597 45247 29631
rect 47670 29628 47676 29640
rect 47631 29600 47676 29628
rect 45189 29591 45247 29597
rect 47670 29588 47676 29600
rect 47728 29588 47734 29640
rect 47857 29631 47915 29637
rect 47857 29597 47869 29631
rect 47903 29628 47915 29631
rect 48038 29628 48044 29640
rect 47903 29600 48044 29628
rect 47903 29597 47915 29600
rect 47857 29591 47915 29597
rect 48038 29588 48044 29600
rect 48096 29588 48102 29640
rect 48498 29628 48504 29640
rect 48459 29600 48504 29628
rect 48498 29588 48504 29600
rect 48556 29588 48562 29640
rect 48774 29628 48780 29640
rect 48735 29600 48780 29628
rect 48774 29588 48780 29600
rect 48832 29588 48838 29640
rect 52086 29628 52092 29640
rect 52047 29600 52092 29628
rect 52086 29588 52092 29600
rect 52144 29588 52150 29640
rect 53006 29628 53012 29640
rect 52967 29600 53012 29628
rect 53006 29588 53012 29600
rect 53064 29588 53070 29640
rect 55306 29628 55312 29640
rect 55267 29600 55312 29628
rect 55306 29588 55312 29600
rect 55364 29588 55370 29640
rect 55674 29628 55680 29640
rect 55635 29600 55680 29628
rect 55674 29588 55680 29600
rect 55732 29588 55738 29640
rect 56318 29628 56324 29640
rect 56279 29600 56324 29628
rect 56318 29588 56324 29600
rect 56376 29588 56382 29640
rect 56796 29637 56824 29668
rect 57333 29665 57345 29668
rect 57379 29665 57391 29699
rect 57333 29659 57391 29665
rect 56781 29631 56839 29637
rect 56781 29597 56793 29631
rect 56827 29597 56839 29631
rect 56781 29591 56839 29597
rect 56962 29588 56968 29640
rect 57020 29628 57026 29640
rect 57241 29631 57299 29637
rect 57241 29628 57253 29631
rect 57020 29600 57253 29628
rect 57020 29588 57026 29600
rect 57241 29597 57253 29600
rect 57287 29597 57299 29631
rect 57241 29591 57299 29597
rect 57517 29631 57575 29637
rect 57517 29597 57529 29631
rect 57563 29597 57575 29631
rect 57517 29591 57575 29597
rect 36464 29532 37320 29560
rect 42613 29563 42671 29569
rect 42613 29529 42625 29563
rect 42659 29560 42671 29563
rect 43070 29560 43076 29572
rect 42659 29532 43076 29560
rect 42659 29529 42671 29532
rect 42613 29523 42671 29529
rect 43070 29520 43076 29532
rect 43128 29520 43134 29572
rect 51534 29560 51540 29572
rect 51495 29532 51540 29560
rect 51534 29520 51540 29532
rect 51592 29520 51598 29572
rect 56042 29520 56048 29572
rect 56100 29560 56106 29572
rect 57532 29560 57560 29591
rect 57698 29588 57704 29640
rect 57756 29628 57762 29640
rect 57793 29631 57851 29637
rect 57793 29628 57805 29631
rect 57756 29600 57805 29628
rect 57756 29588 57762 29600
rect 57793 29597 57805 29600
rect 57839 29597 57851 29631
rect 57793 29591 57851 29597
rect 57882 29588 57888 29640
rect 57940 29628 57946 29640
rect 57977 29631 58035 29637
rect 57977 29628 57989 29631
rect 57940 29600 57989 29628
rect 57940 29588 57946 29600
rect 57977 29597 57989 29600
rect 58023 29597 58035 29631
rect 57977 29591 58035 29597
rect 56100 29532 57560 29560
rect 56100 29520 56106 29532
rect 28166 29492 28172 29504
rect 27724 29464 28172 29492
rect 28166 29452 28172 29464
rect 28224 29452 28230 29504
rect 32306 29492 32312 29504
rect 32267 29464 32312 29492
rect 32306 29452 32312 29464
rect 32364 29452 32370 29504
rect 40494 29492 40500 29504
rect 40455 29464 40500 29492
rect 40494 29452 40500 29464
rect 40552 29452 40558 29504
rect 40865 29495 40923 29501
rect 40865 29461 40877 29495
rect 40911 29492 40923 29495
rect 42426 29492 42432 29504
rect 40911 29464 42432 29492
rect 40911 29461 40923 29464
rect 40865 29455 40923 29461
rect 42426 29452 42432 29464
rect 42484 29492 42490 29504
rect 42813 29495 42871 29501
rect 42813 29492 42825 29495
rect 42484 29464 42825 29492
rect 42484 29452 42490 29464
rect 42813 29461 42825 29464
rect 42859 29461 42871 29495
rect 42813 29455 42871 29461
rect 1104 29402 58880 29424
rect 1104 29350 19574 29402
rect 19626 29350 19638 29402
rect 19690 29350 19702 29402
rect 19754 29350 19766 29402
rect 19818 29350 19830 29402
rect 19882 29350 50294 29402
rect 50346 29350 50358 29402
rect 50410 29350 50422 29402
rect 50474 29350 50486 29402
rect 50538 29350 50550 29402
rect 50602 29350 58880 29402
rect 1104 29328 58880 29350
rect 5629 29291 5687 29297
rect 5629 29257 5641 29291
rect 5675 29288 5687 29291
rect 7285 29291 7343 29297
rect 5675 29260 7144 29288
rect 5675 29257 5687 29260
rect 5629 29251 5687 29257
rect 4338 29180 4344 29232
rect 4396 29220 4402 29232
rect 6914 29220 6920 29232
rect 4396 29192 6920 29220
rect 4396 29180 4402 29192
rect 6914 29180 6920 29192
rect 6972 29180 6978 29232
rect 7116 29229 7144 29260
rect 7285 29257 7297 29291
rect 7331 29288 7343 29291
rect 7466 29288 7472 29300
rect 7331 29260 7472 29288
rect 7331 29257 7343 29260
rect 7285 29251 7343 29257
rect 7466 29248 7472 29260
rect 7524 29248 7530 29300
rect 10965 29291 11023 29297
rect 10428 29260 10916 29288
rect 7101 29223 7159 29229
rect 7101 29189 7113 29223
rect 7147 29220 7159 29223
rect 9122 29220 9128 29232
rect 7147 29192 9128 29220
rect 7147 29189 7159 29192
rect 7101 29183 7159 29189
rect 9122 29180 9128 29192
rect 9180 29180 9186 29232
rect 3326 29112 3332 29164
rect 3384 29152 3390 29164
rect 5261 29155 5319 29161
rect 5261 29152 5273 29155
rect 3384 29124 5273 29152
rect 3384 29112 3390 29124
rect 5261 29121 5273 29124
rect 5307 29121 5319 29155
rect 5261 29115 5319 29121
rect 8938 29112 8944 29164
rect 8996 29152 9002 29164
rect 10428 29161 10456 29260
rect 10502 29180 10508 29232
rect 10560 29220 10566 29232
rect 10560 29192 10824 29220
rect 10560 29180 10566 29192
rect 9309 29155 9367 29161
rect 9309 29152 9321 29155
rect 8996 29124 9321 29152
rect 8996 29112 9002 29124
rect 9309 29121 9321 29124
rect 9355 29121 9367 29155
rect 9309 29115 9367 29121
rect 10413 29155 10471 29161
rect 10413 29121 10425 29155
rect 10459 29121 10471 29155
rect 10594 29152 10600 29164
rect 10555 29124 10600 29152
rect 10413 29115 10471 29121
rect 10594 29112 10600 29124
rect 10652 29112 10658 29164
rect 10796 29161 10824 29192
rect 10689 29155 10747 29161
rect 10689 29121 10701 29155
rect 10735 29121 10747 29155
rect 10689 29115 10747 29121
rect 10781 29155 10839 29161
rect 10781 29121 10793 29155
rect 10827 29121 10839 29155
rect 10888 29152 10916 29260
rect 10965 29257 10977 29291
rect 11011 29288 11023 29291
rect 11011 29260 12296 29288
rect 11011 29257 11023 29260
rect 10965 29251 11023 29257
rect 11146 29152 11152 29164
rect 10888 29124 11152 29152
rect 10781 29115 10839 29121
rect 5353 29087 5411 29093
rect 5353 29053 5365 29087
rect 5399 29084 5411 29087
rect 5718 29084 5724 29096
rect 5399 29056 5724 29084
rect 5399 29053 5411 29056
rect 5353 29047 5411 29053
rect 5718 29044 5724 29056
rect 5776 29044 5782 29096
rect 9766 29044 9772 29096
rect 9824 29084 9830 29096
rect 9824 29056 10456 29084
rect 9824 29044 9830 29056
rect 10428 29028 10456 29056
rect 9493 29019 9551 29025
rect 9493 28985 9505 29019
rect 9539 29016 9551 29019
rect 9858 29016 9864 29028
rect 9539 28988 9864 29016
rect 9539 28985 9551 28988
rect 9493 28979 9551 28985
rect 9858 28976 9864 28988
rect 9916 28976 9922 29028
rect 10410 28976 10416 29028
rect 10468 29016 10474 29028
rect 10704 29016 10732 29115
rect 10796 29084 10824 29115
rect 11146 29112 11152 29124
rect 11204 29112 11210 29164
rect 12268 29152 12296 29260
rect 12618 29248 12624 29300
rect 12676 29288 12682 29300
rect 13078 29288 13084 29300
rect 12676 29260 13084 29288
rect 12676 29248 12682 29260
rect 13078 29248 13084 29260
rect 13136 29248 13142 29300
rect 13446 29248 13452 29300
rect 13504 29288 13510 29300
rect 14090 29288 14096 29300
rect 13504 29260 13584 29288
rect 13504 29248 13510 29260
rect 13556 29161 13584 29260
rect 13648 29260 14096 29288
rect 13648 29161 13676 29260
rect 14090 29248 14096 29260
rect 14148 29248 14154 29300
rect 15013 29291 15071 29297
rect 15013 29257 15025 29291
rect 15059 29288 15071 29291
rect 15562 29288 15568 29300
rect 15059 29260 15568 29288
rect 15059 29257 15071 29260
rect 15013 29251 15071 29257
rect 15562 29248 15568 29260
rect 15620 29248 15626 29300
rect 20533 29291 20591 29297
rect 20533 29288 20545 29291
rect 19168 29260 20545 29288
rect 19168 29232 19196 29260
rect 20533 29257 20545 29260
rect 20579 29257 20591 29291
rect 21174 29288 21180 29300
rect 21135 29260 21180 29288
rect 20533 29251 20591 29257
rect 21174 29248 21180 29260
rect 21232 29248 21238 29300
rect 23106 29248 23112 29300
rect 23164 29288 23170 29300
rect 23569 29291 23627 29297
rect 23569 29288 23581 29291
rect 23164 29260 23581 29288
rect 23164 29248 23170 29260
rect 23569 29257 23581 29260
rect 23615 29257 23627 29291
rect 23569 29251 23627 29257
rect 24854 29248 24860 29300
rect 24912 29288 24918 29300
rect 30745 29291 30803 29297
rect 24912 29260 30328 29288
rect 24912 29248 24918 29260
rect 17034 29180 17040 29232
rect 17092 29220 17098 29232
rect 17954 29220 17960 29232
rect 17092 29192 17960 29220
rect 17092 29180 17098 29192
rect 13906 29161 13912 29164
rect 13364 29155 13422 29161
rect 13364 29152 13376 29155
rect 12268 29124 13376 29152
rect 13364 29121 13376 29124
rect 13410 29121 13422 29155
rect 13364 29115 13422 29121
rect 13505 29155 13584 29161
rect 13505 29121 13517 29155
rect 13551 29124 13584 29155
rect 13633 29155 13691 29161
rect 13551 29121 13563 29124
rect 13505 29115 13563 29121
rect 13633 29121 13645 29155
rect 13679 29121 13691 29155
rect 13633 29115 13691 29121
rect 13725 29155 13783 29161
rect 13725 29121 13737 29155
rect 13771 29121 13783 29155
rect 13725 29115 13783 29121
rect 13863 29155 13912 29161
rect 13863 29121 13875 29155
rect 13909 29121 13912 29155
rect 13863 29115 13912 29121
rect 12069 29087 12127 29093
rect 12069 29084 12081 29087
rect 10796 29056 12081 29084
rect 12069 29053 12081 29056
rect 12115 29053 12127 29087
rect 12069 29047 12127 29053
rect 12345 29087 12403 29093
rect 12345 29053 12357 29087
rect 12391 29053 12403 29087
rect 12345 29047 12403 29053
rect 10468 28988 10732 29016
rect 12360 29016 12388 29047
rect 13740 29028 13768 29115
rect 13906 29112 13912 29115
rect 13964 29112 13970 29164
rect 14461 29155 14519 29161
rect 14461 29121 14473 29155
rect 14507 29121 14519 29155
rect 14642 29152 14648 29164
rect 14603 29124 14648 29152
rect 14461 29115 14519 29121
rect 14476 29084 14504 29115
rect 14642 29112 14648 29124
rect 14700 29112 14706 29164
rect 14734 29112 14740 29164
rect 14792 29152 14798 29164
rect 14918 29161 14924 29164
rect 14875 29155 14924 29161
rect 14792 29124 14837 29152
rect 14792 29112 14798 29124
rect 14875 29121 14887 29155
rect 14921 29121 14924 29155
rect 14875 29115 14924 29121
rect 14918 29112 14924 29115
rect 14976 29112 14982 29164
rect 15470 29152 15476 29164
rect 15431 29124 15476 29152
rect 15470 29112 15476 29124
rect 15528 29112 15534 29164
rect 17512 29161 17540 29192
rect 17954 29180 17960 29192
rect 18012 29220 18018 29232
rect 19150 29220 19156 29232
rect 18012 29192 19156 29220
rect 18012 29180 18018 29192
rect 19150 29180 19156 29192
rect 19208 29180 19214 29232
rect 19426 29180 19432 29232
rect 19484 29220 19490 29232
rect 19889 29223 19947 29229
rect 19889 29220 19901 29223
rect 19484 29192 19901 29220
rect 19484 29180 19490 29192
rect 19889 29189 19901 29192
rect 19935 29189 19947 29223
rect 27062 29220 27068 29232
rect 19889 29183 19947 29189
rect 19996 29192 27068 29220
rect 17497 29155 17555 29161
rect 17497 29121 17509 29155
rect 17543 29121 17555 29155
rect 17497 29115 17555 29121
rect 17586 29112 17592 29164
rect 17644 29152 17650 29164
rect 17773 29155 17831 29161
rect 17773 29152 17785 29155
rect 17644 29124 17785 29152
rect 17644 29112 17650 29124
rect 17773 29121 17785 29124
rect 17819 29121 17831 29155
rect 17773 29115 17831 29121
rect 19242 29112 19248 29164
rect 19300 29152 19306 29164
rect 19996 29152 20024 29192
rect 27062 29180 27068 29192
rect 27120 29180 27126 29232
rect 27172 29192 28856 29220
rect 27172 29164 27200 29192
rect 19300 29124 20024 29152
rect 19300 29112 19306 29124
rect 22738 29112 22744 29164
rect 22796 29152 22802 29164
rect 23477 29155 23535 29161
rect 23477 29152 23489 29155
rect 22796 29124 23489 29152
rect 22796 29112 22802 29124
rect 23477 29121 23489 29124
rect 23523 29121 23535 29155
rect 23477 29115 23535 29121
rect 23661 29155 23719 29161
rect 23661 29121 23673 29155
rect 23707 29152 23719 29155
rect 26973 29155 27031 29161
rect 23707 29124 24440 29152
rect 23707 29121 23719 29124
rect 23661 29115 23719 29121
rect 13832 29056 14596 29084
rect 13630 29016 13636 29028
rect 12360 28988 13636 29016
rect 10468 28976 10474 28988
rect 13630 28976 13636 28988
rect 13688 28976 13694 29028
rect 13722 28976 13728 29028
rect 13780 28976 13786 29028
rect 7101 28951 7159 28957
rect 7101 28917 7113 28951
rect 7147 28948 7159 28951
rect 7374 28948 7380 28960
rect 7147 28920 7380 28948
rect 7147 28917 7159 28920
rect 7101 28911 7159 28917
rect 7374 28908 7380 28920
rect 7432 28908 7438 28960
rect 11974 28908 11980 28960
rect 12032 28948 12038 28960
rect 13832 28948 13860 29056
rect 14001 29019 14059 29025
rect 14001 28985 14013 29019
rect 14047 29016 14059 29019
rect 14182 29016 14188 29028
rect 14047 28988 14188 29016
rect 14047 28985 14059 28988
rect 14001 28979 14059 28985
rect 14182 28976 14188 28988
rect 14240 28976 14246 29028
rect 14568 29016 14596 29056
rect 18598 29044 18604 29096
rect 18656 29084 18662 29096
rect 20073 29087 20131 29093
rect 20073 29084 20085 29087
rect 18656 29056 20085 29084
rect 18656 29044 18662 29056
rect 20073 29053 20085 29056
rect 20119 29084 20131 29087
rect 24118 29084 24124 29096
rect 20119 29056 22094 29084
rect 24079 29056 24124 29084
rect 20119 29053 20131 29056
rect 20073 29047 20131 29053
rect 17218 29016 17224 29028
rect 14568 28988 17224 29016
rect 17218 28976 17224 28988
rect 17276 28976 17282 29028
rect 18046 29016 18052 29028
rect 18007 28988 18052 29016
rect 18046 28976 18052 28988
rect 18104 29016 18110 29028
rect 18506 29016 18512 29028
rect 18104 28988 18512 29016
rect 18104 28976 18110 28988
rect 18506 28976 18512 28988
rect 18564 28976 18570 29028
rect 19334 29016 19340 29028
rect 19295 28988 19340 29016
rect 19334 28976 19340 28988
rect 19392 28976 19398 29028
rect 22066 29016 22094 29056
rect 24118 29044 24124 29056
rect 24176 29044 24182 29096
rect 24412 29093 24440 29124
rect 26973 29121 26985 29155
rect 27019 29121 27031 29155
rect 27154 29152 27160 29164
rect 27115 29124 27160 29152
rect 26973 29115 27031 29121
rect 24397 29087 24455 29093
rect 24397 29053 24409 29087
rect 24443 29084 24455 29087
rect 24578 29084 24584 29096
rect 24443 29056 24584 29084
rect 24443 29053 24455 29056
rect 24397 29047 24455 29053
rect 24578 29044 24584 29056
rect 24636 29044 24642 29096
rect 26421 29087 26479 29093
rect 26421 29053 26433 29087
rect 26467 29084 26479 29087
rect 26988 29084 27016 29115
rect 27154 29112 27160 29124
rect 27212 29112 27218 29164
rect 27893 29155 27951 29161
rect 27893 29121 27905 29155
rect 27939 29152 27951 29155
rect 28074 29152 28080 29164
rect 27939 29124 28080 29152
rect 27939 29121 27951 29124
rect 27893 29115 27951 29121
rect 28074 29112 28080 29124
rect 28132 29112 28138 29164
rect 28166 29112 28172 29164
rect 28224 29152 28230 29164
rect 28828 29161 28856 29192
rect 28813 29155 28871 29161
rect 28224 29124 28269 29152
rect 28224 29112 28230 29124
rect 28813 29121 28825 29155
rect 28859 29121 28871 29155
rect 28813 29115 28871 29121
rect 26467 29056 28120 29084
rect 26467 29053 26479 29056
rect 26421 29047 26479 29053
rect 24302 29016 24308 29028
rect 22066 28988 24308 29016
rect 24302 28976 24308 28988
rect 24360 28976 24366 29028
rect 27157 29019 27215 29025
rect 27157 28985 27169 29019
rect 27203 29016 27215 29019
rect 27706 29016 27712 29028
rect 27203 28988 27712 29016
rect 27203 28985 27215 28988
rect 27157 28979 27215 28985
rect 27706 28976 27712 28988
rect 27764 28976 27770 29028
rect 28092 29016 28120 29056
rect 28258 29044 28264 29096
rect 28316 29084 28322 29096
rect 30300 29093 30328 29260
rect 30745 29257 30757 29291
rect 30791 29288 30803 29291
rect 32214 29288 32220 29300
rect 30791 29260 32220 29288
rect 30791 29257 30803 29260
rect 30745 29251 30803 29257
rect 32214 29248 32220 29260
rect 32272 29248 32278 29300
rect 32309 29291 32367 29297
rect 32309 29257 32321 29291
rect 32355 29288 32367 29291
rect 32674 29288 32680 29300
rect 32355 29260 32680 29288
rect 32355 29257 32367 29260
rect 32309 29251 32367 29257
rect 32674 29248 32680 29260
rect 32732 29248 32738 29300
rect 34425 29291 34483 29297
rect 34425 29257 34437 29291
rect 34471 29288 34483 29291
rect 36446 29288 36452 29300
rect 34471 29260 36452 29288
rect 34471 29257 34483 29260
rect 34425 29251 34483 29257
rect 36446 29248 36452 29260
rect 36504 29248 36510 29300
rect 48774 29248 48780 29300
rect 48832 29288 48838 29300
rect 49602 29288 49608 29300
rect 48832 29260 49608 29288
rect 48832 29248 48838 29260
rect 49602 29248 49608 29260
rect 49660 29248 49666 29300
rect 51718 29288 51724 29300
rect 51679 29260 51724 29288
rect 51718 29248 51724 29260
rect 51776 29248 51782 29300
rect 54941 29291 54999 29297
rect 54941 29257 54953 29291
rect 54987 29288 54999 29291
rect 55306 29288 55312 29300
rect 54987 29260 55312 29288
rect 54987 29257 54999 29260
rect 54941 29251 54999 29257
rect 55306 29248 55312 29260
rect 55364 29248 55370 29300
rect 56318 29248 56324 29300
rect 56376 29288 56382 29300
rect 56873 29291 56931 29297
rect 56873 29288 56885 29291
rect 56376 29260 56885 29288
rect 56376 29248 56382 29260
rect 56873 29257 56885 29260
rect 56919 29257 56931 29291
rect 56873 29251 56931 29257
rect 45002 29220 45008 29232
rect 44744 29192 45008 29220
rect 30377 29155 30435 29161
rect 30377 29121 30389 29155
rect 30423 29152 30435 29155
rect 30926 29152 30932 29164
rect 30423 29124 30932 29152
rect 30423 29121 30435 29124
rect 30377 29115 30435 29121
rect 30926 29112 30932 29124
rect 30984 29112 30990 29164
rect 32214 29152 32220 29164
rect 32175 29124 32220 29152
rect 32214 29112 32220 29124
rect 32272 29112 32278 29164
rect 34057 29155 34115 29161
rect 34057 29121 34069 29155
rect 34103 29152 34115 29155
rect 34514 29152 34520 29164
rect 34103 29124 34520 29152
rect 34103 29121 34115 29124
rect 34057 29115 34115 29121
rect 34514 29112 34520 29124
rect 34572 29152 34578 29164
rect 34885 29155 34943 29161
rect 34885 29152 34897 29155
rect 34572 29124 34897 29152
rect 34572 29112 34578 29124
rect 34885 29121 34897 29124
rect 34931 29121 34943 29155
rect 43070 29152 43076 29164
rect 43031 29124 43076 29152
rect 34885 29115 34943 29121
rect 43070 29112 43076 29124
rect 43128 29112 43134 29164
rect 28629 29087 28687 29093
rect 28629 29084 28641 29087
rect 28316 29056 28641 29084
rect 28316 29044 28322 29056
rect 28629 29053 28641 29056
rect 28675 29053 28687 29087
rect 28629 29047 28687 29053
rect 28997 29087 29055 29093
rect 28997 29053 29009 29087
rect 29043 29053 29055 29087
rect 28997 29047 29055 29053
rect 30285 29087 30343 29093
rect 30285 29053 30297 29087
rect 30331 29053 30343 29087
rect 30285 29047 30343 29053
rect 29012 29016 29040 29047
rect 33134 29044 33140 29096
rect 33192 29084 33198 29096
rect 33965 29087 34023 29093
rect 33965 29084 33977 29087
rect 33192 29056 33977 29084
rect 33192 29044 33198 29056
rect 33965 29053 33977 29056
rect 34011 29053 34023 29087
rect 42886 29084 42892 29096
rect 42847 29056 42892 29084
rect 33965 29047 34023 29053
rect 42886 29044 42892 29056
rect 42944 29044 42950 29096
rect 44744 29093 44772 29192
rect 45002 29180 45008 29192
rect 45060 29180 45066 29232
rect 47670 29180 47676 29232
rect 47728 29220 47734 29232
rect 47728 29192 49280 29220
rect 47728 29180 47734 29192
rect 45097 29155 45155 29161
rect 45097 29121 45109 29155
rect 45143 29152 45155 29155
rect 45462 29152 45468 29164
rect 45143 29124 45468 29152
rect 45143 29121 45155 29124
rect 45097 29115 45155 29121
rect 45462 29112 45468 29124
rect 45520 29112 45526 29164
rect 48409 29155 48467 29161
rect 48409 29121 48421 29155
rect 48455 29152 48467 29155
rect 49142 29152 49148 29164
rect 48455 29124 49148 29152
rect 48455 29121 48467 29124
rect 48409 29115 48467 29121
rect 49142 29112 49148 29124
rect 49200 29112 49206 29164
rect 44729 29087 44787 29093
rect 44729 29053 44741 29087
rect 44775 29053 44787 29087
rect 44729 29047 44787 29053
rect 45005 29087 45063 29093
rect 45005 29053 45017 29087
rect 45051 29084 45063 29087
rect 45186 29084 45192 29096
rect 45051 29056 45192 29084
rect 45051 29053 45063 29056
rect 45005 29047 45063 29053
rect 29270 29016 29276 29028
rect 28092 28988 29276 29016
rect 29270 28976 29276 28988
rect 29328 29016 29334 29028
rect 29457 29019 29515 29025
rect 29457 29016 29469 29019
rect 29328 28988 29469 29016
rect 29328 28976 29334 28988
rect 29457 28985 29469 28988
rect 29503 28985 29515 29019
rect 29457 28979 29515 28985
rect 43257 29019 43315 29025
rect 43257 28985 43269 29019
rect 43303 29016 43315 29019
rect 45020 29016 45048 29047
rect 45186 29044 45192 29056
rect 45244 29044 45250 29096
rect 48498 29084 48504 29096
rect 48459 29056 48504 29084
rect 48498 29044 48504 29056
rect 48556 29044 48562 29096
rect 49252 29093 49280 29192
rect 51074 29180 51080 29232
rect 51132 29220 51138 29232
rect 57606 29220 57612 29232
rect 51132 29192 57612 29220
rect 51132 29180 51138 29192
rect 49421 29155 49479 29161
rect 49421 29121 49433 29155
rect 49467 29121 49479 29155
rect 49421 29115 49479 29121
rect 49237 29087 49295 29093
rect 49237 29053 49249 29087
rect 49283 29053 49295 29087
rect 49237 29047 49295 29053
rect 43303 28988 45048 29016
rect 43303 28985 43315 28988
rect 43257 28979 43315 28985
rect 48406 28976 48412 29028
rect 48464 29016 48470 29028
rect 48777 29019 48835 29025
rect 48777 29016 48789 29019
rect 48464 28988 48789 29016
rect 48464 28976 48470 28988
rect 48777 28985 48789 28988
rect 48823 28985 48835 29019
rect 49436 29016 49464 29115
rect 50890 29112 50896 29164
rect 50948 29152 50954 29164
rect 52104 29161 52132 29192
rect 57606 29180 57612 29192
rect 57664 29180 57670 29232
rect 51905 29155 51963 29161
rect 51905 29152 51917 29155
rect 50948 29124 51917 29152
rect 50948 29112 50954 29124
rect 51905 29121 51917 29124
rect 51951 29121 51963 29155
rect 51905 29115 51963 29121
rect 52089 29155 52147 29161
rect 52089 29121 52101 29155
rect 52135 29121 52147 29155
rect 52089 29115 52147 29121
rect 55677 29155 55735 29161
rect 55677 29121 55689 29155
rect 55723 29152 55735 29155
rect 56042 29152 56048 29164
rect 55723 29124 56048 29152
rect 55723 29121 55735 29124
rect 55677 29115 55735 29121
rect 56042 29112 56048 29124
rect 56100 29112 56106 29164
rect 57333 29155 57391 29161
rect 57333 29121 57345 29155
rect 57379 29152 57391 29155
rect 57882 29152 57888 29164
rect 57379 29124 57888 29152
rect 57379 29121 57391 29124
rect 57333 29115 57391 29121
rect 57882 29112 57888 29124
rect 57940 29112 57946 29164
rect 58158 29152 58164 29164
rect 58119 29124 58164 29152
rect 58158 29112 58164 29124
rect 58216 29112 58222 29164
rect 55766 29044 55772 29096
rect 55824 29084 55830 29096
rect 55861 29087 55919 29093
rect 55861 29084 55873 29087
rect 55824 29056 55873 29084
rect 55824 29044 55830 29056
rect 55861 29053 55873 29056
rect 55907 29084 55919 29087
rect 57698 29084 57704 29096
rect 55907 29056 57704 29084
rect 55907 29053 55919 29056
rect 55861 29047 55919 29053
rect 57698 29044 57704 29056
rect 57756 29044 57762 29096
rect 48777 28979 48835 28985
rect 48884 28988 49464 29016
rect 12032 28920 13860 28948
rect 22189 28951 22247 28957
rect 12032 28908 12038 28920
rect 22189 28917 22201 28951
rect 22235 28948 22247 28951
rect 22462 28948 22468 28960
rect 22235 28920 22468 28948
rect 22235 28917 22247 28920
rect 22189 28911 22247 28917
rect 22462 28908 22468 28920
rect 22520 28948 22526 28960
rect 22649 28951 22707 28957
rect 22649 28948 22661 28951
rect 22520 28920 22661 28948
rect 22520 28908 22526 28920
rect 22649 28917 22661 28920
rect 22695 28917 22707 28951
rect 27614 28948 27620 28960
rect 27575 28920 27620 28948
rect 22649 28911 22707 28917
rect 27614 28908 27620 28920
rect 27672 28908 27678 28960
rect 27890 28908 27896 28960
rect 27948 28948 27954 28960
rect 28077 28951 28135 28957
rect 28077 28948 28089 28951
rect 27948 28920 28089 28948
rect 27948 28908 27954 28920
rect 28077 28917 28089 28920
rect 28123 28948 28135 28951
rect 28626 28948 28632 28960
rect 28123 28920 28632 28948
rect 28123 28917 28135 28920
rect 28077 28911 28135 28917
rect 28626 28908 28632 28920
rect 28684 28908 28690 28960
rect 48038 28908 48044 28960
rect 48096 28948 48102 28960
rect 48884 28948 48912 28988
rect 57422 28976 57428 29028
rect 57480 29016 57486 29028
rect 57977 29019 58035 29025
rect 57977 29016 57989 29019
rect 57480 28988 57989 29016
rect 57480 28976 57486 28988
rect 57977 28985 57989 28988
rect 58023 28985 58035 29019
rect 57977 28979 58035 28985
rect 48096 28920 48912 28948
rect 48096 28908 48102 28920
rect 56962 28908 56968 28960
rect 57020 28948 57026 28960
rect 57057 28951 57115 28957
rect 57057 28948 57069 28951
rect 57020 28920 57069 28948
rect 57020 28908 57026 28920
rect 57057 28917 57069 28920
rect 57103 28917 57115 28951
rect 57057 28911 57115 28917
rect 1104 28858 58880 28880
rect 1104 28806 4214 28858
rect 4266 28806 4278 28858
rect 4330 28806 4342 28858
rect 4394 28806 4406 28858
rect 4458 28806 4470 28858
rect 4522 28806 34934 28858
rect 34986 28806 34998 28858
rect 35050 28806 35062 28858
rect 35114 28806 35126 28858
rect 35178 28806 35190 28858
rect 35242 28806 58880 28858
rect 1104 28784 58880 28806
rect 9125 28747 9183 28753
rect 9125 28713 9137 28747
rect 9171 28744 9183 28747
rect 10594 28744 10600 28756
rect 9171 28716 10600 28744
rect 9171 28713 9183 28716
rect 9125 28707 9183 28713
rect 10594 28704 10600 28716
rect 10652 28744 10658 28756
rect 10778 28744 10784 28756
rect 10652 28716 10784 28744
rect 10652 28704 10658 28716
rect 10778 28704 10784 28716
rect 10836 28704 10842 28756
rect 12158 28704 12164 28756
rect 12216 28744 12222 28756
rect 12342 28744 12348 28756
rect 12216 28716 12348 28744
rect 12216 28704 12222 28716
rect 12342 28704 12348 28716
rect 12400 28704 12406 28756
rect 18601 28747 18659 28753
rect 18601 28713 18613 28747
rect 18647 28744 18659 28747
rect 18782 28744 18788 28756
rect 18647 28716 18788 28744
rect 18647 28713 18659 28716
rect 18601 28707 18659 28713
rect 18782 28704 18788 28716
rect 18840 28704 18846 28756
rect 23753 28747 23811 28753
rect 23753 28713 23765 28747
rect 23799 28744 23811 28747
rect 24854 28744 24860 28756
rect 23799 28716 24860 28744
rect 23799 28713 23811 28716
rect 23753 28707 23811 28713
rect 24854 28704 24860 28716
rect 24912 28704 24918 28756
rect 25225 28747 25283 28753
rect 25225 28713 25237 28747
rect 25271 28744 25283 28747
rect 42518 28744 42524 28756
rect 25271 28716 41414 28744
rect 42479 28716 42524 28744
rect 25271 28713 25283 28716
rect 25225 28707 25283 28713
rect 9858 28676 9864 28688
rect 9771 28648 9864 28676
rect 9858 28636 9864 28648
rect 9916 28676 9922 28688
rect 10686 28676 10692 28688
rect 9916 28648 10692 28676
rect 9916 28636 9922 28648
rect 10686 28636 10692 28648
rect 10744 28676 10750 28688
rect 22738 28676 22744 28688
rect 10744 28648 22744 28676
rect 10744 28636 10750 28648
rect 22738 28636 22744 28648
rect 22796 28636 22802 28688
rect 23842 28636 23848 28688
rect 23900 28676 23906 28688
rect 24581 28679 24639 28685
rect 24581 28676 24593 28679
rect 23900 28648 24593 28676
rect 23900 28636 23906 28648
rect 24581 28645 24593 28648
rect 24627 28676 24639 28679
rect 24762 28676 24768 28688
rect 24627 28648 24768 28676
rect 24627 28645 24639 28648
rect 24581 28639 24639 28645
rect 24762 28636 24768 28648
rect 24820 28636 24826 28688
rect 8938 28540 8944 28552
rect 8899 28512 8944 28540
rect 8938 28500 8944 28512
rect 8996 28500 9002 28552
rect 9122 28540 9128 28552
rect 9083 28512 9128 28540
rect 9122 28500 9128 28512
rect 9180 28500 9186 28552
rect 9674 28540 9680 28552
rect 9635 28512 9680 28540
rect 9674 28500 9680 28512
rect 9732 28500 9738 28552
rect 9876 28549 9904 28636
rect 11974 28608 11980 28620
rect 11935 28580 11980 28608
rect 11974 28568 11980 28580
rect 12032 28568 12038 28620
rect 17126 28608 17132 28620
rect 12406 28580 17132 28608
rect 9861 28543 9919 28549
rect 9861 28509 9873 28543
rect 9907 28509 9919 28543
rect 11146 28540 11152 28552
rect 11107 28512 11152 28540
rect 9861 28503 9919 28509
rect 11146 28500 11152 28512
rect 11204 28500 11210 28552
rect 11422 28500 11428 28552
rect 11480 28540 11486 28552
rect 12158 28540 12164 28552
rect 11480 28512 12164 28540
rect 11480 28500 11486 28512
rect 12158 28500 12164 28512
rect 12216 28540 12222 28552
rect 12253 28543 12311 28549
rect 12253 28540 12265 28543
rect 12216 28512 12265 28540
rect 12216 28500 12222 28512
rect 12253 28509 12265 28512
rect 12299 28509 12311 28543
rect 12253 28503 12311 28509
rect 6730 28432 6736 28484
rect 6788 28472 6794 28484
rect 9953 28475 10011 28481
rect 6788 28444 7696 28472
rect 6788 28432 6794 28444
rect 7006 28404 7012 28416
rect 6967 28376 7012 28404
rect 7006 28364 7012 28376
rect 7064 28364 7070 28416
rect 7668 28413 7696 28444
rect 9953 28441 9965 28475
rect 9999 28472 10011 28475
rect 10502 28472 10508 28484
rect 9999 28444 10508 28472
rect 9999 28441 10011 28444
rect 9953 28435 10011 28441
rect 10502 28432 10508 28444
rect 10560 28432 10566 28484
rect 10686 28432 10692 28484
rect 10744 28472 10750 28484
rect 10965 28475 11023 28481
rect 10965 28472 10977 28475
rect 10744 28444 10977 28472
rect 10744 28432 10750 28444
rect 10965 28441 10977 28444
rect 11011 28441 11023 28475
rect 10965 28435 11023 28441
rect 7653 28407 7711 28413
rect 7653 28373 7665 28407
rect 7699 28404 7711 28407
rect 12406 28404 12434 28580
rect 17126 28568 17132 28580
rect 17184 28568 17190 28620
rect 21082 28608 21088 28620
rect 19628 28580 21088 28608
rect 13446 28500 13452 28552
rect 13504 28540 13510 28552
rect 13722 28540 13728 28552
rect 13504 28512 13728 28540
rect 13504 28500 13510 28512
rect 13722 28500 13728 28512
rect 13780 28540 13786 28552
rect 14645 28543 14703 28549
rect 14645 28540 14657 28543
rect 13780 28512 14657 28540
rect 13780 28500 13786 28512
rect 14645 28509 14657 28512
rect 14691 28540 14703 28543
rect 15010 28540 15016 28552
rect 14691 28512 15016 28540
rect 14691 28509 14703 28512
rect 14645 28503 14703 28509
rect 15010 28500 15016 28512
rect 15068 28500 15074 28552
rect 18509 28543 18567 28549
rect 18509 28509 18521 28543
rect 18555 28509 18567 28543
rect 18509 28503 18567 28509
rect 14550 28404 14556 28416
rect 7699 28376 12434 28404
rect 14511 28376 14556 28404
rect 7699 28373 7711 28376
rect 7653 28367 7711 28373
rect 14550 28364 14556 28376
rect 14608 28364 14614 28416
rect 18524 28404 18552 28503
rect 18598 28500 18604 28552
rect 18656 28540 18662 28552
rect 18693 28543 18751 28549
rect 18693 28540 18705 28543
rect 18656 28512 18705 28540
rect 18656 28500 18662 28512
rect 18693 28509 18705 28512
rect 18739 28509 18751 28543
rect 18693 28503 18751 28509
rect 19334 28500 19340 28552
rect 19392 28540 19398 28552
rect 19628 28540 19656 28580
rect 21082 28568 21088 28580
rect 21140 28568 21146 28620
rect 21545 28611 21603 28617
rect 21545 28577 21557 28611
rect 21591 28577 21603 28611
rect 21545 28571 21603 28577
rect 21821 28611 21879 28617
rect 21821 28577 21833 28611
rect 21867 28608 21879 28611
rect 22278 28608 22284 28620
rect 21867 28580 22284 28608
rect 21867 28577 21879 28580
rect 21821 28571 21879 28577
rect 19392 28526 19656 28540
rect 20257 28543 20315 28549
rect 19392 28512 19642 28526
rect 19392 28500 19398 28512
rect 20257 28509 20269 28543
rect 20303 28540 20315 28543
rect 21453 28543 21511 28549
rect 21453 28540 21465 28543
rect 20303 28512 21465 28540
rect 20303 28509 20315 28512
rect 20257 28503 20315 28509
rect 21453 28509 21465 28512
rect 21499 28509 21511 28543
rect 21560 28540 21588 28571
rect 22278 28568 22284 28580
rect 22336 28568 22342 28620
rect 22557 28611 22615 28617
rect 22557 28577 22569 28611
rect 22603 28577 22615 28611
rect 22557 28571 22615 28577
rect 22462 28540 22468 28552
rect 21560 28512 22468 28540
rect 21453 28503 21511 28509
rect 19426 28432 19432 28484
rect 19484 28472 19490 28484
rect 19521 28475 19579 28481
rect 19521 28472 19533 28475
rect 19484 28444 19533 28472
rect 19484 28432 19490 28444
rect 19521 28441 19533 28444
rect 19567 28441 19579 28475
rect 21468 28472 21496 28503
rect 22462 28500 22468 28512
rect 22520 28500 22526 28552
rect 22572 28484 22600 28571
rect 23658 28540 23664 28552
rect 23619 28512 23664 28540
rect 23658 28500 23664 28512
rect 23716 28500 23722 28552
rect 23845 28543 23903 28549
rect 23845 28509 23857 28543
rect 23891 28540 23903 28543
rect 24302 28540 24308 28552
rect 23891 28512 24308 28540
rect 23891 28509 23903 28512
rect 23845 28503 23903 28509
rect 24302 28500 24308 28512
rect 24360 28500 24366 28552
rect 24397 28543 24455 28549
rect 24397 28509 24409 28543
rect 24443 28540 24455 28543
rect 24578 28540 24584 28552
rect 24443 28512 24584 28540
rect 24443 28509 24455 28512
rect 24397 28503 24455 28509
rect 24578 28500 24584 28512
rect 24636 28500 24642 28552
rect 22002 28472 22008 28484
rect 21468 28444 22008 28472
rect 19521 28435 19579 28441
rect 22002 28432 22008 28444
rect 22060 28432 22066 28484
rect 22094 28432 22100 28484
rect 22152 28472 22158 28484
rect 22554 28472 22560 28484
rect 22152 28444 22560 28472
rect 22152 28432 22158 28444
rect 22554 28432 22560 28444
rect 22612 28472 22618 28484
rect 25240 28472 25268 28707
rect 27433 28679 27491 28685
rect 27433 28645 27445 28679
rect 27479 28676 27491 28679
rect 27614 28676 27620 28688
rect 27479 28648 27620 28676
rect 27479 28645 27491 28648
rect 27433 28639 27491 28645
rect 27614 28636 27620 28648
rect 27672 28636 27678 28688
rect 31573 28679 31631 28685
rect 31573 28645 31585 28679
rect 31619 28676 31631 28679
rect 32306 28676 32312 28688
rect 31619 28648 32312 28676
rect 31619 28645 31631 28648
rect 31573 28639 31631 28645
rect 32306 28636 32312 28648
rect 32364 28636 32370 28688
rect 35253 28679 35311 28685
rect 35253 28645 35265 28679
rect 35299 28676 35311 28679
rect 36630 28676 36636 28688
rect 35299 28648 36636 28676
rect 35299 28645 35311 28648
rect 35253 28639 35311 28645
rect 36630 28636 36636 28648
rect 36688 28636 36694 28688
rect 39209 28679 39267 28685
rect 39209 28645 39221 28679
rect 39255 28676 39267 28679
rect 39666 28676 39672 28688
rect 39255 28648 39672 28676
rect 39255 28645 39267 28648
rect 39209 28639 39267 28645
rect 39666 28636 39672 28648
rect 39724 28636 39730 28688
rect 41386 28676 41414 28716
rect 42518 28704 42524 28716
rect 42576 28704 42582 28756
rect 48498 28744 48504 28756
rect 48459 28716 48504 28744
rect 48498 28704 48504 28716
rect 48556 28704 48562 28756
rect 51258 28704 51264 28756
rect 51316 28744 51322 28756
rect 51353 28747 51411 28753
rect 51353 28744 51365 28747
rect 51316 28716 51365 28744
rect 51316 28704 51322 28716
rect 51353 28713 51365 28716
rect 51399 28713 51411 28747
rect 51353 28707 51411 28713
rect 57609 28747 57667 28753
rect 57609 28713 57621 28747
rect 57655 28744 57667 28747
rect 57882 28744 57888 28756
rect 57655 28716 57888 28744
rect 57655 28713 57667 28716
rect 57609 28707 57667 28713
rect 57882 28704 57888 28716
rect 57940 28704 57946 28756
rect 58158 28744 58164 28756
rect 58119 28716 58164 28744
rect 58158 28704 58164 28716
rect 58216 28704 58222 28756
rect 57790 28676 57796 28688
rect 41386 28648 57796 28676
rect 57790 28636 57796 28648
rect 57848 28636 57854 28688
rect 27709 28611 27767 28617
rect 27709 28577 27721 28611
rect 27755 28608 27767 28611
rect 27798 28608 27804 28620
rect 27755 28580 27804 28608
rect 27755 28577 27767 28580
rect 27709 28571 27767 28577
rect 27798 28568 27804 28580
rect 27856 28568 27862 28620
rect 34606 28568 34612 28620
rect 34664 28608 34670 28620
rect 34793 28611 34851 28617
rect 34793 28608 34805 28611
rect 34664 28580 34805 28608
rect 34664 28568 34670 28580
rect 34793 28577 34805 28580
rect 34839 28577 34851 28611
rect 37550 28608 37556 28620
rect 37463 28580 37556 28608
rect 34793 28571 34851 28577
rect 37550 28568 37556 28580
rect 37608 28608 37614 28620
rect 37921 28611 37979 28617
rect 37608 28580 37872 28608
rect 37608 28568 37614 28580
rect 28169 28543 28227 28549
rect 28169 28509 28181 28543
rect 28215 28509 28227 28543
rect 28169 28503 28227 28509
rect 22612 28444 25268 28472
rect 22612 28432 22618 28444
rect 20070 28404 20076 28416
rect 18524 28376 20076 28404
rect 20070 28364 20076 28376
rect 20128 28364 20134 28416
rect 22830 28404 22836 28416
rect 22791 28376 22836 28404
rect 22830 28364 22836 28376
rect 22888 28364 22894 28416
rect 27246 28404 27252 28416
rect 27207 28376 27252 28404
rect 27246 28364 27252 28376
rect 27304 28364 27310 28416
rect 27706 28364 27712 28416
rect 27764 28404 27770 28416
rect 28184 28404 28212 28503
rect 28258 28500 28264 28552
rect 28316 28540 28322 28552
rect 28353 28543 28411 28549
rect 28353 28540 28365 28543
rect 28316 28512 28365 28540
rect 28316 28500 28322 28512
rect 28353 28509 28365 28512
rect 28399 28509 28411 28543
rect 28353 28503 28411 28509
rect 34885 28543 34943 28549
rect 34885 28509 34897 28543
rect 34931 28540 34943 28543
rect 35342 28540 35348 28552
rect 34931 28512 35348 28540
rect 34931 28509 34943 28512
rect 34885 28503 34943 28509
rect 35342 28500 35348 28512
rect 35400 28500 35406 28552
rect 37734 28540 37740 28552
rect 37695 28512 37740 28540
rect 37734 28500 37740 28512
rect 37792 28500 37798 28552
rect 31205 28475 31263 28481
rect 31205 28472 31217 28475
rect 30668 28444 31217 28472
rect 28534 28404 28540 28416
rect 27764 28376 28212 28404
rect 28495 28376 28540 28404
rect 27764 28364 27770 28376
rect 28534 28364 28540 28376
rect 28592 28364 28598 28416
rect 30374 28364 30380 28416
rect 30432 28404 30438 28416
rect 30668 28413 30696 28444
rect 31205 28441 31217 28444
rect 31251 28441 31263 28475
rect 31386 28472 31392 28484
rect 31347 28444 31392 28472
rect 31205 28435 31263 28441
rect 31386 28432 31392 28444
rect 31444 28432 31450 28484
rect 37844 28472 37872 28580
rect 37921 28577 37933 28611
rect 37967 28608 37979 28611
rect 38749 28611 38807 28617
rect 38749 28608 38761 28611
rect 37967 28580 38761 28608
rect 37967 28577 37979 28580
rect 37921 28571 37979 28577
rect 38749 28577 38761 28580
rect 38795 28608 38807 28611
rect 39114 28608 39120 28620
rect 38795 28580 39120 28608
rect 38795 28577 38807 28580
rect 38749 28571 38807 28577
rect 39114 28568 39120 28580
rect 39172 28568 39178 28620
rect 42245 28611 42303 28617
rect 42245 28577 42257 28611
rect 42291 28608 42303 28611
rect 42886 28608 42892 28620
rect 42291 28580 42892 28608
rect 42291 28577 42303 28580
rect 42245 28571 42303 28577
rect 42886 28568 42892 28580
rect 42944 28568 42950 28620
rect 45186 28568 45192 28620
rect 45244 28608 45250 28620
rect 45244 28580 45692 28608
rect 45244 28568 45250 28580
rect 38841 28543 38899 28549
rect 38841 28509 38853 28543
rect 38887 28540 38899 28543
rect 39298 28540 39304 28552
rect 38887 28512 39304 28540
rect 38887 28509 38899 28512
rect 38841 28503 38899 28509
rect 39298 28500 39304 28512
rect 39356 28500 39362 28552
rect 42334 28540 42340 28552
rect 42295 28512 42340 28540
rect 42334 28500 42340 28512
rect 42392 28500 42398 28552
rect 45462 28540 45468 28552
rect 45423 28512 45468 28540
rect 45462 28500 45468 28512
rect 45520 28500 45526 28552
rect 45664 28549 45692 28580
rect 51350 28568 51356 28620
rect 51408 28608 51414 28620
rect 51408 28580 51580 28608
rect 51408 28568 51414 28580
rect 45649 28543 45707 28549
rect 45649 28509 45661 28543
rect 45695 28509 45707 28543
rect 48038 28540 48044 28552
rect 47999 28512 48044 28540
rect 45649 28503 45707 28509
rect 48038 28500 48044 28512
rect 48096 28500 48102 28552
rect 48314 28540 48320 28552
rect 48275 28512 48320 28540
rect 48314 28500 48320 28512
rect 48372 28500 48378 28552
rect 49326 28500 49332 28552
rect 49384 28540 49390 28552
rect 49421 28543 49479 28549
rect 49421 28540 49433 28543
rect 49384 28512 49433 28540
rect 49384 28500 49390 28512
rect 49421 28509 49433 28512
rect 49467 28509 49479 28543
rect 49602 28540 49608 28552
rect 49563 28512 49608 28540
rect 49421 28503 49479 28509
rect 49602 28500 49608 28512
rect 49660 28500 49666 28552
rect 51552 28549 51580 28580
rect 51537 28543 51595 28549
rect 51537 28509 51549 28543
rect 51583 28509 51595 28543
rect 51537 28503 51595 28509
rect 57149 28543 57207 28549
rect 57149 28509 57161 28543
rect 57195 28540 57207 28543
rect 57238 28540 57244 28552
rect 57195 28512 57244 28540
rect 57195 28509 57207 28512
rect 57149 28503 57207 28509
rect 57238 28500 57244 28512
rect 57296 28500 57302 28552
rect 57422 28540 57428 28552
rect 57383 28512 57428 28540
rect 57422 28500 57428 28512
rect 57480 28500 57486 28552
rect 45557 28475 45615 28481
rect 37844 28444 41414 28472
rect 30653 28407 30711 28413
rect 30653 28404 30665 28407
rect 30432 28376 30665 28404
rect 30432 28364 30438 28376
rect 30653 28373 30665 28376
rect 30699 28373 30711 28407
rect 41386 28404 41414 28444
rect 45557 28441 45569 28475
rect 45603 28472 45615 28475
rect 47670 28472 47676 28484
rect 45603 28444 47676 28472
rect 45603 28441 45615 28444
rect 45557 28435 45615 28441
rect 47670 28432 47676 28444
rect 47728 28472 47734 28484
rect 48133 28475 48191 28481
rect 48133 28472 48145 28475
rect 47728 28444 48145 28472
rect 47728 28432 47734 28444
rect 48133 28441 48145 28444
rect 48179 28441 48191 28475
rect 51258 28472 51264 28484
rect 51219 28444 51264 28472
rect 48133 28435 48191 28441
rect 51258 28432 51264 28444
rect 51316 28432 51322 28484
rect 51445 28475 51503 28481
rect 51445 28441 51457 28475
rect 51491 28441 51503 28475
rect 51445 28435 51503 28441
rect 41874 28404 41880 28416
rect 41386 28376 41880 28404
rect 30653 28367 30711 28373
rect 41874 28364 41880 28376
rect 41932 28364 41938 28416
rect 49605 28407 49663 28413
rect 49605 28373 49617 28407
rect 49651 28404 49663 28407
rect 51460 28404 51488 28435
rect 51626 28404 51632 28416
rect 49651 28376 51632 28404
rect 49651 28373 49663 28376
rect 49605 28367 49663 28373
rect 51626 28364 51632 28376
rect 51684 28364 51690 28416
rect 56042 28364 56048 28416
rect 56100 28404 56106 28416
rect 56137 28407 56195 28413
rect 56137 28404 56149 28407
rect 56100 28376 56149 28404
rect 56100 28364 56106 28376
rect 56137 28373 56149 28376
rect 56183 28373 56195 28407
rect 56137 28367 56195 28373
rect 57241 28407 57299 28413
rect 57241 28373 57253 28407
rect 57287 28404 57299 28407
rect 57974 28404 57980 28416
rect 57287 28376 57980 28404
rect 57287 28373 57299 28376
rect 57241 28367 57299 28373
rect 57974 28364 57980 28376
rect 58032 28364 58038 28416
rect 1104 28314 58880 28336
rect 1104 28262 19574 28314
rect 19626 28262 19638 28314
rect 19690 28262 19702 28314
rect 19754 28262 19766 28314
rect 19818 28262 19830 28314
rect 19882 28262 50294 28314
rect 50346 28262 50358 28314
rect 50410 28262 50422 28314
rect 50474 28262 50486 28314
rect 50538 28262 50550 28314
rect 50602 28262 58880 28314
rect 1104 28240 58880 28262
rect 6717 28203 6775 28209
rect 6717 28169 6729 28203
rect 6763 28200 6775 28203
rect 9769 28203 9827 28209
rect 6763 28172 7604 28200
rect 6763 28169 6775 28172
rect 6717 28163 6775 28169
rect 6917 28135 6975 28141
rect 6917 28101 6929 28135
rect 6963 28132 6975 28135
rect 7006 28132 7012 28144
rect 6963 28104 7012 28132
rect 6963 28101 6975 28104
rect 6917 28095 6975 28101
rect 3697 28067 3755 28073
rect 3697 28033 3709 28067
rect 3743 28033 3755 28067
rect 6932 28064 6960 28095
rect 7006 28092 7012 28104
rect 7064 28092 7070 28144
rect 7576 28141 7604 28172
rect 9769 28169 9781 28203
rect 9815 28200 9827 28203
rect 13722 28200 13728 28212
rect 9815 28172 13728 28200
rect 9815 28169 9827 28172
rect 9769 28163 9827 28169
rect 13722 28160 13728 28172
rect 13780 28160 13786 28212
rect 13814 28160 13820 28212
rect 13872 28200 13878 28212
rect 14369 28203 14427 28209
rect 14369 28200 14381 28203
rect 13872 28172 14381 28200
rect 13872 28160 13878 28172
rect 14369 28169 14381 28172
rect 14415 28169 14427 28203
rect 25406 28200 25412 28212
rect 25367 28172 25412 28200
rect 14369 28163 14427 28169
rect 25406 28160 25412 28172
rect 25464 28160 25470 28212
rect 31389 28203 31447 28209
rect 31389 28169 31401 28203
rect 31435 28200 31447 28203
rect 32214 28200 32220 28212
rect 31435 28172 32220 28200
rect 31435 28169 31447 28172
rect 31389 28163 31447 28169
rect 32214 28160 32220 28172
rect 32272 28160 32278 28212
rect 36725 28203 36783 28209
rect 36725 28169 36737 28203
rect 36771 28200 36783 28203
rect 37734 28200 37740 28212
rect 36771 28172 37740 28200
rect 36771 28169 36783 28172
rect 36725 28163 36783 28169
rect 37734 28160 37740 28172
rect 37792 28160 37798 28212
rect 42889 28203 42947 28209
rect 42889 28169 42901 28203
rect 42935 28200 42947 28203
rect 43070 28200 43076 28212
rect 42935 28172 43076 28200
rect 42935 28169 42947 28172
rect 42889 28163 42947 28169
rect 43070 28160 43076 28172
rect 43128 28160 43134 28212
rect 51350 28160 51356 28212
rect 51408 28160 51414 28212
rect 55309 28203 55367 28209
rect 55309 28169 55321 28203
rect 55355 28200 55367 28203
rect 55674 28200 55680 28212
rect 55355 28172 55680 28200
rect 55355 28169 55367 28172
rect 55309 28163 55367 28169
rect 55674 28160 55680 28172
rect 55732 28160 55738 28212
rect 56962 28200 56968 28212
rect 56923 28172 56968 28200
rect 56962 28160 56968 28172
rect 57020 28160 57026 28212
rect 7561 28135 7619 28141
rect 7561 28101 7573 28135
rect 7607 28132 7619 28135
rect 8202 28132 8208 28144
rect 7607 28104 8208 28132
rect 7607 28101 7619 28104
rect 7561 28095 7619 28101
rect 8202 28092 8208 28104
rect 8260 28092 8266 28144
rect 8389 28135 8447 28141
rect 8389 28101 8401 28135
rect 8435 28132 8447 28135
rect 10410 28132 10416 28144
rect 8435 28104 10416 28132
rect 8435 28101 8447 28104
rect 8389 28095 8447 28101
rect 10410 28092 10416 28104
rect 10468 28092 10474 28144
rect 15013 28135 15071 28141
rect 15013 28132 15025 28135
rect 13740 28104 15025 28132
rect 8478 28064 8484 28076
rect 6932 28036 8484 28064
rect 3697 28027 3755 28033
rect 2777 27999 2835 28005
rect 2777 27965 2789 27999
rect 2823 27996 2835 27999
rect 2958 27996 2964 28008
rect 2823 27968 2964 27996
rect 2823 27965 2835 27968
rect 2777 27959 2835 27965
rect 2958 27956 2964 27968
rect 3016 27956 3022 28008
rect 3050 27956 3056 28008
rect 3108 27996 3114 28008
rect 3108 27968 3153 27996
rect 3108 27956 3114 27968
rect 3326 27956 3332 28008
rect 3384 27996 3390 28008
rect 3605 27999 3663 28005
rect 3605 27996 3617 27999
rect 3384 27968 3617 27996
rect 3384 27956 3390 27968
rect 3605 27965 3617 27968
rect 3651 27965 3663 27999
rect 3605 27959 3663 27965
rect 3712 27928 3740 28027
rect 8478 28024 8484 28036
rect 8536 28024 8542 28076
rect 9585 28067 9643 28073
rect 9585 28033 9597 28067
rect 9631 28064 9643 28067
rect 9674 28064 9680 28076
rect 9631 28036 9680 28064
rect 9631 28033 9643 28036
rect 9585 28027 9643 28033
rect 9674 28024 9680 28036
rect 9732 28024 9738 28076
rect 13740 28008 13768 28104
rect 15013 28101 15025 28104
rect 15059 28101 15071 28135
rect 15013 28095 15071 28101
rect 15102 28092 15108 28144
rect 15160 28132 15166 28144
rect 19242 28132 19248 28144
rect 15160 28104 19248 28132
rect 15160 28092 15166 28104
rect 19242 28092 19248 28104
rect 19300 28092 19306 28144
rect 24762 28092 24768 28144
rect 24820 28132 24826 28144
rect 27798 28132 27804 28144
rect 24820 28104 27804 28132
rect 24820 28092 24826 28104
rect 27798 28092 27804 28104
rect 27856 28092 27862 28144
rect 41601 28135 41659 28141
rect 41601 28101 41613 28135
rect 41647 28132 41659 28135
rect 51368 28132 51396 28160
rect 51445 28135 51503 28141
rect 51445 28132 51457 28135
rect 41647 28104 42748 28132
rect 51368 28104 51457 28132
rect 41647 28101 41659 28104
rect 41601 28095 41659 28101
rect 13909 28067 13967 28073
rect 13909 28033 13921 28067
rect 13955 28064 13967 28067
rect 13998 28064 14004 28076
rect 13955 28036 14004 28064
rect 13955 28033 13967 28036
rect 13909 28027 13967 28033
rect 13998 28024 14004 28036
rect 14056 28024 14062 28076
rect 14645 28067 14703 28073
rect 14645 28033 14657 28067
rect 14691 28033 14703 28067
rect 14645 28027 14703 28033
rect 14921 28067 14979 28073
rect 14921 28033 14933 28067
rect 14967 28064 14979 28067
rect 15194 28064 15200 28076
rect 14967 28036 15200 28064
rect 14967 28033 14979 28036
rect 14921 28027 14979 28033
rect 4065 27999 4123 28005
rect 4065 27965 4077 27999
rect 4111 27996 4123 27999
rect 8938 27996 8944 28008
rect 4111 27968 8944 27996
rect 4111 27965 4123 27968
rect 4065 27959 4123 27965
rect 8938 27956 8944 27968
rect 8996 27996 9002 28008
rect 9401 27999 9459 28005
rect 9401 27996 9413 27999
rect 8996 27968 9413 27996
rect 8996 27956 9002 27968
rect 9401 27965 9413 27968
rect 9447 27965 9459 27999
rect 9401 27959 9459 27965
rect 13633 27999 13691 28005
rect 13633 27965 13645 27999
rect 13679 27996 13691 27999
rect 13722 27996 13728 28008
rect 13679 27968 13728 27996
rect 13679 27965 13691 27968
rect 13633 27959 13691 27965
rect 13722 27956 13728 27968
rect 13780 27956 13786 28008
rect 14553 27999 14611 28005
rect 14553 27965 14565 27999
rect 14599 27965 14611 27999
rect 14660 27996 14688 28027
rect 15194 28024 15200 28036
rect 15252 28064 15258 28076
rect 16206 28064 16212 28076
rect 15252 28036 16212 28064
rect 15252 28024 15258 28036
rect 16206 28024 16212 28036
rect 16264 28024 16270 28076
rect 16945 28067 17003 28073
rect 16945 28033 16957 28067
rect 16991 28064 17003 28067
rect 17034 28064 17040 28076
rect 16991 28036 17040 28064
rect 16991 28033 17003 28036
rect 16945 28027 17003 28033
rect 17034 28024 17040 28036
rect 17092 28024 17098 28076
rect 17218 28064 17224 28076
rect 17179 28036 17224 28064
rect 17218 28024 17224 28036
rect 17276 28024 17282 28076
rect 22278 28024 22284 28076
rect 22336 28064 22342 28076
rect 22465 28067 22523 28073
rect 22465 28064 22477 28067
rect 22336 28036 22477 28064
rect 22336 28024 22342 28036
rect 22465 28033 22477 28036
rect 22511 28033 22523 28067
rect 22465 28027 22523 28033
rect 24118 28024 24124 28076
rect 24176 28064 24182 28076
rect 24673 28067 24731 28073
rect 24673 28064 24685 28067
rect 24176 28036 24685 28064
rect 24176 28024 24182 28036
rect 24673 28033 24685 28036
rect 24719 28033 24731 28067
rect 24673 28027 24731 28033
rect 24857 28067 24915 28073
rect 24857 28033 24869 28067
rect 24903 28033 24915 28067
rect 24857 28027 24915 28033
rect 20717 27999 20775 28005
rect 14660 27968 15608 27996
rect 14553 27959 14611 27965
rect 4617 27931 4675 27937
rect 4617 27928 4629 27931
rect 3712 27900 4629 27928
rect 4617 27897 4629 27900
rect 4663 27928 4675 27931
rect 4890 27928 4896 27940
rect 4663 27900 4896 27928
rect 4663 27897 4675 27900
rect 4617 27891 4675 27897
rect 4890 27888 4896 27900
rect 4948 27928 4954 27940
rect 4948 27900 6776 27928
rect 4948 27888 4954 27900
rect 6748 27872 6776 27900
rect 8018 27888 8024 27940
rect 8076 27928 8082 27940
rect 8205 27931 8263 27937
rect 8205 27928 8217 27931
rect 8076 27900 8217 27928
rect 8076 27888 8082 27900
rect 8205 27897 8217 27900
rect 8251 27897 8263 27931
rect 8205 27891 8263 27897
rect 10502 27888 10508 27940
rect 10560 27928 10566 27940
rect 14458 27928 14464 27940
rect 10560 27900 14464 27928
rect 10560 27888 10566 27900
rect 14458 27888 14464 27900
rect 14516 27928 14522 27940
rect 14568 27928 14596 27959
rect 14516 27900 14596 27928
rect 14516 27888 14522 27900
rect 6454 27820 6460 27872
rect 6512 27860 6518 27872
rect 6549 27863 6607 27869
rect 6549 27860 6561 27863
rect 6512 27832 6561 27860
rect 6512 27820 6518 27832
rect 6549 27829 6561 27832
rect 6595 27829 6607 27863
rect 6730 27860 6736 27872
rect 6691 27832 6736 27860
rect 6549 27823 6607 27829
rect 6730 27820 6736 27832
rect 6788 27820 6794 27872
rect 7466 27860 7472 27872
rect 7427 27832 7472 27860
rect 7466 27820 7472 27832
rect 7524 27820 7530 27872
rect 12250 27820 12256 27872
rect 12308 27860 12314 27872
rect 15194 27860 15200 27872
rect 12308 27832 15200 27860
rect 12308 27820 12314 27832
rect 15194 27820 15200 27832
rect 15252 27820 15258 27872
rect 15580 27869 15608 27968
rect 20717 27965 20729 27999
rect 20763 27996 20775 27999
rect 22002 27996 22008 28008
rect 20763 27968 22008 27996
rect 20763 27965 20775 27968
rect 20717 27959 20775 27965
rect 22002 27956 22008 27968
rect 22060 27956 22066 28008
rect 22741 27999 22799 28005
rect 22741 27965 22753 27999
rect 22787 27996 22799 27999
rect 23658 27996 23664 28008
rect 22787 27968 23664 27996
rect 22787 27965 22799 27968
rect 22741 27959 22799 27965
rect 23658 27956 23664 27968
rect 23716 27956 23722 28008
rect 24210 27956 24216 28008
rect 24268 27996 24274 28008
rect 24872 27996 24900 28027
rect 25130 28024 25136 28076
rect 25188 28064 25194 28076
rect 25317 28067 25375 28073
rect 25317 28064 25329 28067
rect 25188 28036 25329 28064
rect 25188 28024 25194 28036
rect 25317 28033 25329 28036
rect 25363 28033 25375 28067
rect 25317 28027 25375 28033
rect 25501 28067 25559 28073
rect 25501 28033 25513 28067
rect 25547 28033 25559 28067
rect 25501 28027 25559 28033
rect 25516 27996 25544 28027
rect 30742 28024 30748 28076
rect 30800 28064 30806 28076
rect 31021 28067 31079 28073
rect 31021 28064 31033 28067
rect 30800 28036 31033 28064
rect 30800 28024 30806 28036
rect 31021 28033 31033 28036
rect 31067 28064 31079 28067
rect 31386 28064 31392 28076
rect 31067 28036 31392 28064
rect 31067 28033 31079 28036
rect 31021 28027 31079 28033
rect 31386 28024 31392 28036
rect 31444 28024 31450 28076
rect 36354 28064 36360 28076
rect 36315 28036 36360 28064
rect 36354 28024 36360 28036
rect 36412 28024 36418 28076
rect 36446 28024 36452 28076
rect 36504 28064 36510 28076
rect 36541 28067 36599 28073
rect 36541 28064 36553 28067
rect 36504 28036 36553 28064
rect 36504 28024 36510 28036
rect 36541 28033 36553 28036
rect 36587 28033 36599 28067
rect 39114 28064 39120 28076
rect 39075 28036 39120 28064
rect 36541 28027 36599 28033
rect 39114 28024 39120 28036
rect 39172 28024 39178 28076
rect 39298 28064 39304 28076
rect 39259 28036 39304 28064
rect 39298 28024 39304 28036
rect 39356 28024 39362 28076
rect 41046 28064 41052 28076
rect 41007 28036 41052 28064
rect 41046 28024 41052 28036
rect 41104 28024 41110 28076
rect 41138 28024 41144 28076
rect 41196 28064 41202 28076
rect 41322 28064 41328 28076
rect 41196 28036 41241 28064
rect 41283 28036 41328 28064
rect 41196 28024 41202 28036
rect 41322 28024 41328 28036
rect 41380 28024 41386 28076
rect 41417 28067 41475 28073
rect 41417 28033 41429 28067
rect 41463 28033 41475 28067
rect 41417 28027 41475 28033
rect 25961 27999 26019 28005
rect 25961 27996 25973 27999
rect 24268 27968 25973 27996
rect 24268 27956 24274 27968
rect 25961 27965 25973 27968
rect 26007 27965 26019 27999
rect 25961 27959 26019 27965
rect 30374 27956 30380 28008
rect 30432 27996 30438 28008
rect 30929 27999 30987 28005
rect 30929 27996 30941 27999
rect 30432 27968 30941 27996
rect 30432 27956 30438 27968
rect 30929 27965 30941 27968
rect 30975 27965 30987 27999
rect 30929 27959 30987 27965
rect 39209 27999 39267 28005
rect 39209 27965 39221 27999
rect 39255 27996 39267 27999
rect 41230 27996 41236 28008
rect 39255 27968 41236 27996
rect 39255 27965 39267 27968
rect 39209 27959 39267 27965
rect 41230 27956 41236 27968
rect 41288 27996 41294 28008
rect 41432 27996 41460 28027
rect 41874 28024 41880 28076
rect 41932 28064 41938 28076
rect 42720 28073 42748 28104
rect 51445 28101 51457 28104
rect 51491 28101 51503 28135
rect 51445 28095 51503 28101
rect 57133 28135 57191 28141
rect 57133 28101 57145 28135
rect 57179 28132 57191 28135
rect 57238 28132 57244 28144
rect 57179 28104 57244 28132
rect 57179 28101 57191 28104
rect 57133 28095 57191 28101
rect 57238 28092 57244 28104
rect 57296 28092 57302 28144
rect 57333 28135 57391 28141
rect 57333 28101 57345 28135
rect 57379 28132 57391 28135
rect 57422 28132 57428 28144
rect 57379 28104 57428 28132
rect 57379 28101 57391 28104
rect 57333 28095 57391 28101
rect 57422 28092 57428 28104
rect 57480 28092 57486 28144
rect 42521 28067 42579 28073
rect 42521 28064 42533 28067
rect 41932 28036 42533 28064
rect 41932 28024 41938 28036
rect 42521 28033 42533 28036
rect 42567 28033 42579 28067
rect 42521 28027 42579 28033
rect 42613 28067 42671 28073
rect 42613 28033 42625 28067
rect 42659 28033 42671 28067
rect 42613 28027 42671 28033
rect 42705 28067 42763 28073
rect 42705 28033 42717 28067
rect 42751 28064 42763 28067
rect 42886 28064 42892 28076
rect 42751 28036 42892 28064
rect 42751 28033 42763 28036
rect 42705 28027 42763 28033
rect 41288 27968 41460 27996
rect 41288 27956 41294 27968
rect 42334 27956 42340 28008
rect 42392 27996 42398 28008
rect 42628 27996 42656 28027
rect 42886 28024 42892 28036
rect 42944 28024 42950 28076
rect 44729 28067 44787 28073
rect 44729 28033 44741 28067
rect 44775 28064 44787 28067
rect 44910 28064 44916 28076
rect 44775 28036 44916 28064
rect 44775 28033 44787 28036
rect 44729 28027 44787 28033
rect 44910 28024 44916 28036
rect 44968 28024 44974 28076
rect 51074 28024 51080 28076
rect 51132 28064 51138 28076
rect 51225 28067 51283 28073
rect 51132 28036 51177 28064
rect 51132 28024 51138 28036
rect 51225 28033 51237 28067
rect 51271 28064 51283 28067
rect 51271 28033 51304 28064
rect 51225 28027 51304 28033
rect 45002 27996 45008 28008
rect 42392 27968 42656 27996
rect 44963 27968 45008 27996
rect 42392 27956 42398 27968
rect 45002 27956 45008 27968
rect 45060 27956 45066 28008
rect 17126 27888 17132 27940
rect 17184 27928 17190 27940
rect 37642 27928 37648 27940
rect 17184 27900 37648 27928
rect 17184 27888 17190 27900
rect 37642 27888 37648 27900
rect 37700 27888 37706 27940
rect 44821 27931 44879 27937
rect 44821 27897 44833 27931
rect 44867 27928 44879 27931
rect 45094 27928 45100 27940
rect 44867 27900 45100 27928
rect 44867 27897 44879 27900
rect 44821 27891 44879 27897
rect 45094 27888 45100 27900
rect 45152 27888 45158 27940
rect 15565 27863 15623 27869
rect 15565 27829 15577 27863
rect 15611 27860 15623 27863
rect 18046 27860 18052 27872
rect 15611 27832 18052 27860
rect 15611 27829 15623 27832
rect 15565 27823 15623 27829
rect 18046 27820 18052 27832
rect 18104 27860 18110 27872
rect 18233 27863 18291 27869
rect 18233 27860 18245 27863
rect 18104 27832 18245 27860
rect 18104 27820 18110 27832
rect 18233 27829 18245 27832
rect 18279 27829 18291 27863
rect 24210 27860 24216 27872
rect 24171 27832 24216 27860
rect 18233 27823 18291 27829
rect 24210 27820 24216 27832
rect 24268 27820 24274 27872
rect 24765 27863 24823 27869
rect 24765 27829 24777 27863
rect 24811 27860 24823 27863
rect 25038 27860 25044 27872
rect 24811 27832 25044 27860
rect 24811 27829 24823 27832
rect 24765 27823 24823 27829
rect 25038 27820 25044 27832
rect 25096 27820 25102 27872
rect 29638 27860 29644 27872
rect 29599 27832 29644 27860
rect 29638 27820 29644 27832
rect 29696 27820 29702 27872
rect 30374 27860 30380 27872
rect 30335 27832 30380 27860
rect 30374 27820 30380 27832
rect 30432 27820 30438 27872
rect 44913 27863 44971 27869
rect 44913 27829 44925 27863
rect 44959 27860 44971 27863
rect 46842 27860 46848 27872
rect 44959 27832 46848 27860
rect 44959 27829 44971 27832
rect 44913 27823 44971 27829
rect 46842 27820 46848 27832
rect 46900 27820 46906 27872
rect 51276 27860 51304 28027
rect 51350 28024 51356 28076
rect 51408 28064 51414 28076
rect 51626 28073 51632 28076
rect 51583 28067 51632 28073
rect 51408 28036 51453 28064
rect 51408 28024 51414 28036
rect 51583 28033 51595 28067
rect 51629 28033 51632 28067
rect 51583 28027 51632 28033
rect 51626 28024 51632 28027
rect 51684 28024 51690 28076
rect 55306 28024 55312 28076
rect 55364 28064 55370 28076
rect 55493 28067 55551 28073
rect 55493 28064 55505 28067
rect 55364 28036 55505 28064
rect 55364 28024 55370 28036
rect 55493 28033 55505 28036
rect 55539 28033 55551 28067
rect 55493 28027 55551 28033
rect 55582 28024 55588 28076
rect 55640 28064 55646 28076
rect 55640 28036 55685 28064
rect 55640 28024 55646 28036
rect 55858 28024 55864 28076
rect 55916 28064 55922 28076
rect 55953 28067 56011 28073
rect 55953 28064 55965 28067
rect 55916 28036 55965 28064
rect 55916 28024 55922 28036
rect 55953 28033 55965 28036
rect 55999 28033 56011 28067
rect 55953 28027 56011 28033
rect 55677 27999 55735 28005
rect 55677 27965 55689 27999
rect 55723 27965 55735 27999
rect 55677 27959 55735 27965
rect 55692 27928 55720 27959
rect 55766 27956 55772 28008
rect 55824 27996 55830 28008
rect 55824 27968 55869 27996
rect 55824 27956 55830 27968
rect 56962 27928 56968 27940
rect 55692 27900 56968 27928
rect 56962 27888 56968 27900
rect 57020 27888 57026 27940
rect 51442 27860 51448 27872
rect 51276 27832 51448 27860
rect 51442 27820 51448 27832
rect 51500 27820 51506 27872
rect 51718 27860 51724 27872
rect 51679 27832 51724 27860
rect 51718 27820 51724 27832
rect 51776 27820 51782 27872
rect 57149 27863 57207 27869
rect 57149 27829 57161 27863
rect 57195 27860 57207 27863
rect 57974 27860 57980 27872
rect 57195 27832 57980 27860
rect 57195 27829 57207 27832
rect 57149 27823 57207 27829
rect 57974 27820 57980 27832
rect 58032 27820 58038 27872
rect 1104 27770 58880 27792
rect 1104 27718 4214 27770
rect 4266 27718 4278 27770
rect 4330 27718 4342 27770
rect 4394 27718 4406 27770
rect 4458 27718 4470 27770
rect 4522 27718 34934 27770
rect 34986 27718 34998 27770
rect 35050 27718 35062 27770
rect 35114 27718 35126 27770
rect 35178 27718 35190 27770
rect 35242 27718 58880 27770
rect 1104 27696 58880 27718
rect 3050 27616 3056 27668
rect 3108 27656 3114 27668
rect 3237 27659 3295 27665
rect 3237 27656 3249 27659
rect 3108 27628 3249 27656
rect 3108 27616 3114 27628
rect 3237 27625 3249 27628
rect 3283 27656 3295 27659
rect 27246 27656 27252 27668
rect 3283 27628 27252 27656
rect 3283 27625 3295 27628
rect 3237 27619 3295 27625
rect 27246 27616 27252 27628
rect 27304 27616 27310 27668
rect 41046 27616 41052 27668
rect 41104 27656 41110 27668
rect 45462 27656 45468 27668
rect 41104 27628 41552 27656
rect 45423 27628 45468 27656
rect 41104 27616 41110 27628
rect 2038 27588 2044 27600
rect 1999 27560 2044 27588
rect 2038 27548 2044 27560
rect 2096 27548 2102 27600
rect 5629 27591 5687 27597
rect 5629 27557 5641 27591
rect 5675 27588 5687 27591
rect 7466 27588 7472 27600
rect 5675 27560 5856 27588
rect 5675 27557 5687 27560
rect 5629 27551 5687 27557
rect 2501 27523 2559 27529
rect 2501 27489 2513 27523
rect 2547 27520 2559 27523
rect 2774 27520 2780 27532
rect 2547 27492 2780 27520
rect 2547 27489 2559 27492
rect 2501 27483 2559 27489
rect 2774 27480 2780 27492
rect 2832 27480 2838 27532
rect 2409 27455 2467 27461
rect 2409 27421 2421 27455
rect 2455 27452 2467 27455
rect 3970 27452 3976 27464
rect 2455 27424 3976 27452
rect 2455 27421 2467 27424
rect 2409 27415 2467 27421
rect 3970 27412 3976 27424
rect 4028 27452 4034 27464
rect 5534 27452 5540 27464
rect 4028 27424 5540 27452
rect 4028 27412 4034 27424
rect 5534 27412 5540 27424
rect 5592 27412 5598 27464
rect 5626 27384 5632 27396
rect 5587 27356 5632 27384
rect 5626 27344 5632 27356
rect 5684 27344 5690 27396
rect 5828 27384 5856 27560
rect 5920 27560 7472 27588
rect 5920 27461 5948 27560
rect 7466 27548 7472 27560
rect 7524 27588 7530 27600
rect 13262 27588 13268 27600
rect 7524 27560 13268 27588
rect 7524 27548 7530 27560
rect 13262 27548 13268 27560
rect 13320 27548 13326 27600
rect 14366 27548 14372 27600
rect 14424 27588 14430 27600
rect 14737 27591 14795 27597
rect 14737 27588 14749 27591
rect 14424 27560 14749 27588
rect 14424 27548 14430 27560
rect 14737 27557 14749 27560
rect 14783 27557 14795 27591
rect 15286 27588 15292 27600
rect 15247 27560 15292 27588
rect 14737 27551 14795 27557
rect 15286 27548 15292 27560
rect 15344 27548 15350 27600
rect 16853 27591 16911 27597
rect 16853 27557 16865 27591
rect 16899 27557 16911 27591
rect 17034 27588 17040 27600
rect 16995 27560 17040 27588
rect 16853 27551 16911 27557
rect 6917 27523 6975 27529
rect 6917 27489 6929 27523
rect 6963 27520 6975 27523
rect 11238 27520 11244 27532
rect 6963 27492 11244 27520
rect 6963 27489 6975 27492
rect 6917 27483 6975 27489
rect 11238 27480 11244 27492
rect 11296 27480 11302 27532
rect 13173 27523 13231 27529
rect 13173 27489 13185 27523
rect 13219 27520 13231 27523
rect 15304 27520 15332 27548
rect 13219 27492 14136 27520
rect 13219 27489 13231 27492
rect 13173 27483 13231 27489
rect 5905 27455 5963 27461
rect 5905 27421 5917 27455
rect 5951 27421 5963 27455
rect 5905 27415 5963 27421
rect 6365 27455 6423 27461
rect 6365 27421 6377 27455
rect 6411 27421 6423 27455
rect 6365 27415 6423 27421
rect 6380 27384 6408 27415
rect 6454 27412 6460 27464
rect 6512 27452 6518 27464
rect 6641 27455 6699 27461
rect 6512 27424 6557 27452
rect 6512 27412 6518 27424
rect 6641 27421 6653 27455
rect 6687 27421 6699 27455
rect 6641 27415 6699 27421
rect 6733 27455 6791 27461
rect 6733 27421 6745 27455
rect 6779 27452 6791 27455
rect 8018 27452 8024 27464
rect 6779 27424 8024 27452
rect 6779 27421 6791 27424
rect 6733 27415 6791 27421
rect 5828 27356 6408 27384
rect 6656 27384 6684 27415
rect 8018 27412 8024 27424
rect 8076 27412 8082 27464
rect 8389 27455 8447 27461
rect 8389 27421 8401 27455
rect 8435 27452 8447 27455
rect 8478 27452 8484 27464
rect 8435 27424 8484 27452
rect 8435 27421 8447 27424
rect 8389 27415 8447 27421
rect 8478 27412 8484 27424
rect 8536 27452 8542 27464
rect 8938 27452 8944 27464
rect 8536 27424 8944 27452
rect 8536 27412 8542 27424
rect 8938 27412 8944 27424
rect 8996 27412 9002 27464
rect 11790 27452 11796 27464
rect 10520 27424 11796 27452
rect 10520 27393 10548 27424
rect 11790 27412 11796 27424
rect 11848 27452 11854 27464
rect 13078 27452 13084 27464
rect 11848 27424 12434 27452
rect 13039 27424 13084 27452
rect 11848 27412 11854 27424
rect 7653 27387 7711 27393
rect 7653 27384 7665 27387
rect 6656 27356 7665 27384
rect 7653 27353 7665 27356
rect 7699 27384 7711 27387
rect 8297 27387 8355 27393
rect 8297 27384 8309 27387
rect 7699 27356 8309 27384
rect 7699 27353 7711 27356
rect 7653 27347 7711 27353
rect 8297 27353 8309 27356
rect 8343 27353 8355 27387
rect 10505 27387 10563 27393
rect 10505 27384 10517 27387
rect 8297 27347 8355 27353
rect 8864 27356 10517 27384
rect 5813 27319 5871 27325
rect 5813 27285 5825 27319
rect 5859 27316 5871 27319
rect 6270 27316 6276 27328
rect 5859 27288 6276 27316
rect 5859 27285 5871 27288
rect 5813 27279 5871 27285
rect 6270 27276 6276 27288
rect 6328 27276 6334 27328
rect 7190 27276 7196 27328
rect 7248 27316 7254 27328
rect 7561 27319 7619 27325
rect 7561 27316 7573 27319
rect 7248 27288 7573 27316
rect 7248 27276 7254 27288
rect 7561 27285 7573 27288
rect 7607 27285 7619 27319
rect 7561 27279 7619 27285
rect 8110 27276 8116 27328
rect 8168 27316 8174 27328
rect 8864 27316 8892 27356
rect 10505 27353 10517 27356
rect 10551 27353 10563 27387
rect 10686 27384 10692 27396
rect 10647 27356 10692 27384
rect 10505 27347 10563 27353
rect 10686 27344 10692 27356
rect 10744 27344 10750 27396
rect 12406 27384 12434 27424
rect 13078 27412 13084 27424
rect 13136 27412 13142 27464
rect 14108 27461 14136 27492
rect 14384 27492 15332 27520
rect 16577 27523 16635 27529
rect 13265 27455 13323 27461
rect 13265 27421 13277 27455
rect 13311 27421 13323 27455
rect 13265 27415 13323 27421
rect 14093 27455 14151 27461
rect 14093 27421 14105 27455
rect 14139 27421 14151 27455
rect 14274 27452 14280 27464
rect 14235 27424 14280 27452
rect 14093 27415 14151 27421
rect 13280 27384 13308 27415
rect 14274 27412 14280 27424
rect 14332 27412 14338 27464
rect 14384 27461 14412 27492
rect 16577 27489 16589 27523
rect 16623 27520 16635 27523
rect 16758 27520 16764 27532
rect 16623 27492 16764 27520
rect 16623 27489 16635 27492
rect 16577 27483 16635 27489
rect 16758 27480 16764 27492
rect 16816 27480 16822 27532
rect 14369 27455 14427 27461
rect 14369 27421 14381 27455
rect 14415 27421 14427 27455
rect 14369 27415 14427 27421
rect 14458 27412 14464 27464
rect 14516 27452 14522 27464
rect 14516 27424 14561 27452
rect 14516 27412 14522 27424
rect 12406 27356 13308 27384
rect 16868 27384 16896 27551
rect 17034 27548 17040 27560
rect 17092 27548 17098 27600
rect 17586 27588 17592 27600
rect 17547 27560 17592 27588
rect 17586 27548 17592 27560
rect 17644 27548 17650 27600
rect 22741 27591 22799 27597
rect 22741 27557 22753 27591
rect 22787 27588 22799 27591
rect 22830 27588 22836 27600
rect 22787 27560 22836 27588
rect 22787 27557 22799 27560
rect 22741 27551 22799 27557
rect 22830 27548 22836 27560
rect 22888 27548 22894 27600
rect 30926 27588 30932 27600
rect 25424 27560 28672 27588
rect 30887 27560 30932 27588
rect 16942 27480 16948 27532
rect 17000 27520 17006 27532
rect 17604 27520 17632 27548
rect 17000 27492 17632 27520
rect 17000 27480 17006 27492
rect 20346 27480 20352 27532
rect 20404 27520 20410 27532
rect 20993 27523 21051 27529
rect 20993 27520 21005 27523
rect 20404 27492 21005 27520
rect 20404 27480 20410 27492
rect 20993 27489 21005 27492
rect 21039 27520 21051 27523
rect 22002 27520 22008 27532
rect 21039 27492 22008 27520
rect 21039 27489 21051 27492
rect 20993 27483 21051 27489
rect 22002 27480 22008 27492
rect 22060 27480 22066 27532
rect 22278 27480 22284 27532
rect 22336 27520 22342 27532
rect 22373 27523 22431 27529
rect 22373 27520 22385 27523
rect 22336 27492 22385 27520
rect 22336 27480 22342 27492
rect 22373 27489 22385 27492
rect 22419 27489 22431 27523
rect 22373 27483 22431 27489
rect 20162 27412 20168 27464
rect 20220 27452 20226 27464
rect 20806 27452 20812 27464
rect 20220 27424 20812 27452
rect 20220 27412 20226 27424
rect 20806 27412 20812 27424
rect 20864 27452 20870 27464
rect 22848 27452 22876 27548
rect 25038 27520 25044 27532
rect 24999 27492 25044 27520
rect 25038 27480 25044 27492
rect 25096 27480 25102 27532
rect 23385 27455 23443 27461
rect 23385 27452 23397 27455
rect 20864 27424 22094 27452
rect 22848 27424 23397 27452
rect 20864 27412 20870 27424
rect 17954 27384 17960 27396
rect 16868 27356 17960 27384
rect 8168 27288 8892 27316
rect 8168 27276 8174 27288
rect 8938 27276 8944 27328
rect 8996 27316 9002 27328
rect 13280 27316 13308 27356
rect 17954 27344 17960 27356
rect 18012 27384 18018 27396
rect 22066 27384 22094 27424
rect 23385 27421 23397 27424
rect 23431 27421 23443 27455
rect 23658 27452 23664 27464
rect 23619 27424 23664 27452
rect 23385 27415 23443 27421
rect 23658 27412 23664 27424
rect 23716 27412 23722 27464
rect 25130 27452 25136 27464
rect 25091 27424 25136 27452
rect 25130 27412 25136 27424
rect 25188 27412 25194 27464
rect 25424 27384 25452 27560
rect 25501 27523 25559 27529
rect 25501 27489 25513 27523
rect 25547 27520 25559 27523
rect 25547 27492 27016 27520
rect 25547 27489 25559 27492
rect 25501 27483 25559 27489
rect 26142 27452 26148 27464
rect 26103 27424 26148 27452
rect 26142 27412 26148 27424
rect 26200 27412 26206 27464
rect 26344 27461 26372 27492
rect 26988 27461 27016 27492
rect 26329 27455 26387 27461
rect 26329 27421 26341 27455
rect 26375 27421 26387 27455
rect 26329 27415 26387 27421
rect 26789 27455 26847 27461
rect 26789 27421 26801 27455
rect 26835 27421 26847 27455
rect 26789 27415 26847 27421
rect 26973 27455 27031 27461
rect 26973 27421 26985 27455
rect 27019 27421 27031 27455
rect 26973 27415 27031 27421
rect 27157 27455 27215 27461
rect 27157 27421 27169 27455
rect 27203 27452 27215 27455
rect 27430 27452 27436 27464
rect 27203 27424 27436 27452
rect 27203 27421 27215 27424
rect 27157 27415 27215 27421
rect 18012 27356 18184 27384
rect 22066 27356 25452 27384
rect 26160 27384 26188 27412
rect 26804 27384 26832 27415
rect 27430 27412 27436 27424
rect 27488 27452 27494 27464
rect 27893 27455 27951 27461
rect 27893 27452 27905 27455
rect 27488 27424 27905 27452
rect 27488 27412 27494 27424
rect 27893 27421 27905 27424
rect 27939 27421 27951 27455
rect 28074 27452 28080 27464
rect 28035 27424 28080 27452
rect 27893 27415 27951 27421
rect 28074 27412 28080 27424
rect 28132 27412 28138 27464
rect 28353 27455 28411 27461
rect 28353 27421 28365 27455
rect 28399 27452 28411 27455
rect 28534 27452 28540 27464
rect 28399 27424 28540 27452
rect 28399 27421 28411 27424
rect 28353 27415 28411 27421
rect 28534 27412 28540 27424
rect 28592 27412 28598 27464
rect 28644 27452 28672 27560
rect 30926 27548 30932 27560
rect 30984 27588 30990 27600
rect 32858 27588 32864 27600
rect 30984 27560 32864 27588
rect 30984 27548 30990 27560
rect 32858 27548 32864 27560
rect 32916 27548 32922 27600
rect 33045 27591 33103 27597
rect 33045 27557 33057 27591
rect 33091 27588 33103 27591
rect 36354 27588 36360 27600
rect 33091 27560 36360 27588
rect 33091 27557 33103 27560
rect 33045 27551 33103 27557
rect 32585 27523 32643 27529
rect 32585 27520 32597 27523
rect 31726 27492 32597 27520
rect 29638 27452 29644 27464
rect 28644 27424 29644 27452
rect 29638 27412 29644 27424
rect 29696 27452 29702 27464
rect 29825 27455 29883 27461
rect 29825 27452 29837 27455
rect 29696 27424 29837 27452
rect 29696 27412 29702 27424
rect 29825 27421 29837 27424
rect 29871 27421 29883 27455
rect 29825 27415 29883 27421
rect 30101 27455 30159 27461
rect 30101 27421 30113 27455
rect 30147 27452 30159 27455
rect 30742 27452 30748 27464
rect 30147 27424 30748 27452
rect 30147 27421 30159 27424
rect 30101 27415 30159 27421
rect 30742 27412 30748 27424
rect 30800 27412 30806 27464
rect 26160 27356 26832 27384
rect 18012 27344 18018 27356
rect 17310 27316 17316 27328
rect 8996 27288 9041 27316
rect 13280 27288 17316 27316
rect 8996 27276 9002 27288
rect 17310 27276 17316 27288
rect 17368 27276 17374 27328
rect 18156 27325 18184 27356
rect 26878 27344 26884 27396
rect 26936 27384 26942 27396
rect 31726 27384 31754 27492
rect 32585 27489 32597 27492
rect 32631 27489 32643 27523
rect 33597 27523 33655 27529
rect 33597 27520 33609 27523
rect 32585 27483 32643 27489
rect 32692 27492 33609 27520
rect 32692 27461 32720 27492
rect 33597 27489 33609 27492
rect 33643 27520 33655 27523
rect 34514 27520 34520 27532
rect 33643 27492 34520 27520
rect 33643 27489 33655 27492
rect 33597 27483 33655 27489
rect 34514 27480 34520 27492
rect 34572 27520 34578 27532
rect 34698 27520 34704 27532
rect 34572 27492 34704 27520
rect 34572 27480 34578 27492
rect 34698 27480 34704 27492
rect 34756 27480 34762 27532
rect 36280 27461 36308 27560
rect 36354 27548 36360 27560
rect 36412 27548 36418 27600
rect 38565 27591 38623 27597
rect 38565 27557 38577 27591
rect 38611 27588 38623 27591
rect 39298 27588 39304 27600
rect 38611 27560 39304 27588
rect 38611 27557 38623 27560
rect 38565 27551 38623 27557
rect 39298 27548 39304 27560
rect 39356 27548 39362 27600
rect 41524 27597 41552 27628
rect 45462 27616 45468 27628
rect 45520 27616 45526 27668
rect 48314 27616 48320 27668
rect 48372 27656 48378 27668
rect 48685 27659 48743 27665
rect 48685 27656 48697 27659
rect 48372 27628 48697 27656
rect 48372 27616 48378 27628
rect 48685 27625 48697 27628
rect 48731 27656 48743 27659
rect 49142 27656 49148 27668
rect 48731 27628 49148 27656
rect 48731 27625 48743 27628
rect 48685 27619 48743 27625
rect 49142 27616 49148 27628
rect 49200 27616 49206 27668
rect 51258 27616 51264 27668
rect 51316 27656 51322 27668
rect 51445 27659 51503 27665
rect 51445 27656 51457 27659
rect 51316 27628 51457 27656
rect 51316 27616 51322 27628
rect 51445 27625 51457 27628
rect 51491 27625 51503 27659
rect 51445 27619 51503 27625
rect 41509 27591 41567 27597
rect 39408 27560 41414 27588
rect 38102 27520 38108 27532
rect 38063 27492 38108 27520
rect 38102 27480 38108 27492
rect 38160 27480 38166 27532
rect 32677 27455 32735 27461
rect 32677 27421 32689 27455
rect 32723 27421 32735 27455
rect 32677 27415 32735 27421
rect 36265 27455 36323 27461
rect 36265 27421 36277 27455
rect 36311 27421 36323 27455
rect 36265 27415 36323 27421
rect 36446 27412 36452 27464
rect 36504 27452 36510 27464
rect 38194 27452 38200 27464
rect 36504 27424 36549 27452
rect 38155 27424 38200 27452
rect 36504 27412 36510 27424
rect 38194 27412 38200 27424
rect 38252 27412 38258 27464
rect 39408 27384 39436 27560
rect 41230 27520 41236 27532
rect 41191 27492 41236 27520
rect 41230 27480 41236 27492
rect 41288 27480 41294 27532
rect 41386 27520 41414 27560
rect 41509 27557 41521 27591
rect 41555 27557 41567 27591
rect 41509 27551 41567 27557
rect 47765 27591 47823 27597
rect 47765 27557 47777 27591
rect 47811 27588 47823 27591
rect 48038 27588 48044 27600
rect 47811 27560 48044 27588
rect 47811 27557 47823 27560
rect 47765 27551 47823 27557
rect 48038 27548 48044 27560
rect 48096 27548 48102 27600
rect 48501 27591 48559 27597
rect 48501 27557 48513 27591
rect 48547 27557 48559 27591
rect 48501 27551 48559 27557
rect 45094 27520 45100 27532
rect 41386 27492 41828 27520
rect 45055 27492 45100 27520
rect 40862 27412 40868 27464
rect 40920 27452 40926 27464
rect 41322 27452 41328 27464
rect 40920 27424 41328 27452
rect 40920 27412 40926 27424
rect 41322 27412 41328 27424
rect 41380 27412 41386 27464
rect 41601 27455 41659 27461
rect 41601 27421 41613 27455
rect 41647 27421 41659 27455
rect 41601 27415 41659 27421
rect 26936 27356 31754 27384
rect 33152 27356 39436 27384
rect 26936 27344 26942 27356
rect 18141 27319 18199 27325
rect 18141 27285 18153 27319
rect 18187 27316 18199 27319
rect 18874 27316 18880 27328
rect 18187 27288 18880 27316
rect 18187 27285 18199 27288
rect 18141 27279 18199 27285
rect 18874 27276 18880 27288
rect 18932 27276 18938 27328
rect 19242 27276 19248 27328
rect 19300 27316 19306 27328
rect 22738 27316 22744 27328
rect 19300 27288 22744 27316
rect 19300 27276 19306 27288
rect 22738 27276 22744 27288
rect 22796 27276 22802 27328
rect 22833 27319 22891 27325
rect 22833 27285 22845 27319
rect 22879 27316 22891 27319
rect 22922 27316 22928 27328
rect 22879 27288 22928 27316
rect 22879 27285 22891 27288
rect 22833 27279 22891 27285
rect 22922 27276 22928 27288
rect 22980 27276 22986 27328
rect 23382 27316 23388 27328
rect 23343 27288 23388 27316
rect 23382 27276 23388 27288
rect 23440 27276 23446 27328
rect 26234 27316 26240 27328
rect 26195 27288 26240 27316
rect 26234 27276 26240 27288
rect 26292 27276 26298 27328
rect 28537 27319 28595 27325
rect 28537 27285 28549 27319
rect 28583 27316 28595 27319
rect 28626 27316 28632 27328
rect 28583 27288 28632 27316
rect 28583 27285 28595 27288
rect 28537 27279 28595 27285
rect 28626 27276 28632 27288
rect 28684 27276 28690 27328
rect 28718 27276 28724 27328
rect 28776 27316 28782 27328
rect 33152 27316 33180 27356
rect 41138 27344 41144 27396
rect 41196 27384 41202 27396
rect 41616 27384 41644 27415
rect 41196 27356 41644 27384
rect 41800 27384 41828 27492
rect 45094 27480 45100 27492
rect 45152 27480 45158 27532
rect 46842 27480 46848 27532
rect 46900 27520 46906 27532
rect 47305 27523 47363 27529
rect 47305 27520 47317 27523
rect 46900 27492 47317 27520
rect 46900 27480 46906 27492
rect 47305 27489 47317 27492
rect 47351 27520 47363 27523
rect 48516 27520 48544 27551
rect 51902 27548 51908 27600
rect 51960 27588 51966 27600
rect 52362 27588 52368 27600
rect 51960 27560 52368 27588
rect 51960 27548 51966 27560
rect 52362 27548 52368 27560
rect 52420 27548 52426 27600
rect 56962 27588 56968 27600
rect 52472 27560 56640 27588
rect 56923 27560 56968 27588
rect 52472 27520 52500 27560
rect 47351 27492 48544 27520
rect 48608 27492 52500 27520
rect 54588 27492 55536 27520
rect 47351 27489 47363 27492
rect 47305 27483 47363 27489
rect 44910 27412 44916 27464
rect 44968 27452 44974 27464
rect 45189 27455 45247 27461
rect 45189 27452 45201 27455
rect 44968 27424 45201 27452
rect 44968 27412 44974 27424
rect 45189 27421 45201 27424
rect 45235 27421 45247 27455
rect 47394 27452 47400 27464
rect 47355 27424 47400 27452
rect 45189 27415 45247 27421
rect 47394 27412 47400 27424
rect 47452 27412 47458 27464
rect 48608 27452 48636 27492
rect 49142 27452 49148 27464
rect 47504 27424 48636 27452
rect 49103 27424 49148 27452
rect 47504 27384 47532 27424
rect 49142 27412 49148 27424
rect 49200 27412 49206 27464
rect 49326 27452 49332 27464
rect 49287 27424 49332 27452
rect 49326 27412 49332 27424
rect 49384 27412 49390 27464
rect 50706 27412 50712 27464
rect 50764 27452 50770 27464
rect 50985 27455 51043 27461
rect 50985 27452 50997 27455
rect 50764 27424 50997 27452
rect 50764 27412 50770 27424
rect 50985 27421 50997 27424
rect 51031 27421 51043 27455
rect 51258 27452 51264 27464
rect 51219 27424 51264 27452
rect 50985 27415 51043 27421
rect 47946 27384 47952 27396
rect 41800 27356 47532 27384
rect 47596 27356 47952 27384
rect 41196 27344 41202 27356
rect 28776 27288 33180 27316
rect 36449 27319 36507 27325
rect 28776 27276 28782 27288
rect 36449 27285 36461 27319
rect 36495 27316 36507 27319
rect 37550 27316 37556 27328
rect 36495 27288 37556 27316
rect 36495 27285 36507 27288
rect 36449 27279 36507 27285
rect 37550 27276 37556 27288
rect 37608 27276 37614 27328
rect 41233 27319 41291 27325
rect 41233 27285 41245 27319
rect 41279 27316 41291 27319
rect 42334 27316 42340 27328
rect 41279 27288 42340 27316
rect 41279 27285 41291 27288
rect 41233 27279 41291 27285
rect 42334 27276 42340 27288
rect 42392 27276 42398 27328
rect 47394 27276 47400 27328
rect 47452 27316 47458 27328
rect 47596 27316 47624 27356
rect 47946 27344 47952 27356
rect 48004 27384 48010 27396
rect 48225 27387 48283 27393
rect 48225 27384 48237 27387
rect 48004 27356 48237 27384
rect 48004 27344 48010 27356
rect 48225 27353 48237 27356
rect 48271 27353 48283 27387
rect 51000 27384 51028 27415
rect 51258 27412 51264 27424
rect 51316 27412 51322 27464
rect 51718 27412 51724 27464
rect 51776 27452 51782 27464
rect 52181 27455 52239 27461
rect 52181 27452 52193 27455
rect 51776 27424 52193 27452
rect 51776 27412 51782 27424
rect 52181 27421 52193 27424
rect 52227 27452 52239 27455
rect 53926 27452 53932 27464
rect 52227 27424 53932 27452
rect 52227 27421 52239 27424
rect 52181 27415 52239 27421
rect 53926 27412 53932 27424
rect 53984 27412 53990 27464
rect 54113 27455 54171 27461
rect 54113 27421 54125 27455
rect 54159 27452 54171 27455
rect 54588 27452 54616 27492
rect 54159 27424 54616 27452
rect 54665 27455 54723 27461
rect 54159 27421 54171 27424
rect 54113 27415 54171 27421
rect 54665 27421 54677 27455
rect 54711 27452 54723 27455
rect 55306 27452 55312 27464
rect 54711 27424 55312 27452
rect 54711 27421 54723 27424
rect 54665 27415 54723 27421
rect 55306 27412 55312 27424
rect 55364 27412 55370 27464
rect 55508 27461 55536 27492
rect 55950 27480 55956 27532
rect 56008 27520 56014 27532
rect 56505 27523 56563 27529
rect 56505 27520 56517 27523
rect 56008 27492 56517 27520
rect 56008 27480 56014 27492
rect 56505 27489 56517 27492
rect 56551 27489 56563 27523
rect 56612 27520 56640 27560
rect 56962 27548 56968 27560
rect 57020 27548 57026 27600
rect 57977 27591 58035 27597
rect 57977 27557 57989 27591
rect 58023 27557 58035 27591
rect 57977 27551 58035 27557
rect 57992 27520 58020 27551
rect 56612 27492 58020 27520
rect 56505 27483 56563 27489
rect 55493 27455 55551 27461
rect 55493 27421 55505 27455
rect 55539 27452 55551 27455
rect 55582 27452 55588 27464
rect 55539 27424 55588 27452
rect 55539 27421 55551 27424
rect 55493 27415 55551 27421
rect 55582 27412 55588 27424
rect 55640 27412 55646 27464
rect 55769 27455 55827 27461
rect 55769 27421 55781 27455
rect 55815 27421 55827 27455
rect 56594 27452 56600 27464
rect 56555 27424 56600 27452
rect 55769 27415 55827 27421
rect 51350 27384 51356 27396
rect 51000 27356 51356 27384
rect 48225 27347 48283 27353
rect 51350 27344 51356 27356
rect 51408 27344 51414 27396
rect 52638 27344 52644 27396
rect 52696 27384 52702 27396
rect 52696 27356 53222 27384
rect 52696 27344 52702 27356
rect 55122 27344 55128 27396
rect 55180 27384 55186 27396
rect 55784 27384 55812 27415
rect 56594 27412 56600 27424
rect 56652 27412 56658 27464
rect 58158 27452 58164 27464
rect 58119 27424 58164 27452
rect 58158 27412 58164 27424
rect 58216 27412 58222 27464
rect 55180 27356 55812 27384
rect 55180 27344 55186 27356
rect 47452 27288 47624 27316
rect 49237 27319 49295 27325
rect 47452 27276 47458 27288
rect 49237 27285 49249 27319
rect 49283 27316 49295 27319
rect 51077 27319 51135 27325
rect 51077 27316 51089 27319
rect 49283 27288 51089 27316
rect 49283 27285 49295 27288
rect 49237 27279 49295 27285
rect 51077 27285 51089 27288
rect 51123 27316 51135 27319
rect 51166 27316 51172 27328
rect 51123 27288 51172 27316
rect 51123 27285 51135 27288
rect 51077 27279 51135 27285
rect 51166 27276 51172 27288
rect 51224 27276 51230 27328
rect 55953 27319 56011 27325
rect 55953 27285 55965 27319
rect 55999 27316 56011 27319
rect 56870 27316 56876 27328
rect 55999 27288 56876 27316
rect 55999 27285 56011 27288
rect 55953 27279 56011 27285
rect 56870 27276 56876 27288
rect 56928 27276 56934 27328
rect 1104 27226 58880 27248
rect 1104 27174 19574 27226
rect 19626 27174 19638 27226
rect 19690 27174 19702 27226
rect 19754 27174 19766 27226
rect 19818 27174 19830 27226
rect 19882 27174 50294 27226
rect 50346 27174 50358 27226
rect 50410 27174 50422 27226
rect 50474 27174 50486 27226
rect 50538 27174 50550 27226
rect 50602 27174 58880 27226
rect 1104 27152 58880 27174
rect 5626 27072 5632 27124
rect 5684 27112 5690 27124
rect 5813 27115 5871 27121
rect 5813 27112 5825 27115
rect 5684 27084 5825 27112
rect 5684 27072 5690 27084
rect 5813 27081 5825 27084
rect 5859 27112 5871 27115
rect 6638 27112 6644 27124
rect 5859 27084 6644 27112
rect 5859 27081 5871 27084
rect 5813 27075 5871 27081
rect 6638 27072 6644 27084
rect 6696 27072 6702 27124
rect 7282 27072 7288 27124
rect 7340 27112 7346 27124
rect 7377 27115 7435 27121
rect 7377 27112 7389 27115
rect 7340 27084 7389 27112
rect 7340 27072 7346 27084
rect 7377 27081 7389 27084
rect 7423 27081 7435 27115
rect 7377 27075 7435 27081
rect 7837 27115 7895 27121
rect 7837 27081 7849 27115
rect 7883 27081 7895 27115
rect 7837 27075 7895 27081
rect 1854 27044 1860 27056
rect 1815 27016 1860 27044
rect 1854 27004 1860 27016
rect 1912 27004 1918 27056
rect 5169 27047 5227 27053
rect 5169 27013 5181 27047
rect 5215 27044 5227 27047
rect 6730 27044 6736 27056
rect 5215 27016 6736 27044
rect 5215 27013 5227 27016
rect 5169 27007 5227 27013
rect 5644 26985 5672 27016
rect 6730 27004 6736 27016
rect 6788 27004 6794 27056
rect 7852 27044 7880 27075
rect 10134 27072 10140 27124
rect 10192 27112 10198 27124
rect 13081 27115 13139 27121
rect 13081 27112 13093 27115
rect 10192 27084 13093 27112
rect 10192 27072 10198 27084
rect 13081 27081 13093 27084
rect 13127 27112 13139 27115
rect 14642 27112 14648 27124
rect 13127 27084 14648 27112
rect 13127 27081 13139 27084
rect 13081 27075 13139 27081
rect 14642 27072 14648 27084
rect 14700 27072 14706 27124
rect 15102 27112 15108 27124
rect 15063 27084 15108 27112
rect 15102 27072 15108 27084
rect 15160 27072 15166 27124
rect 15470 27072 15476 27124
rect 15528 27112 15534 27124
rect 17957 27115 18015 27121
rect 17957 27112 17969 27115
rect 15528 27084 17969 27112
rect 15528 27072 15534 27084
rect 17957 27081 17969 27084
rect 18003 27112 18015 27115
rect 18414 27112 18420 27124
rect 18003 27084 18420 27112
rect 18003 27081 18015 27084
rect 17957 27075 18015 27081
rect 18414 27072 18420 27084
rect 18472 27072 18478 27124
rect 19058 27112 19064 27124
rect 19019 27084 19064 27112
rect 19058 27072 19064 27084
rect 19116 27072 19122 27124
rect 19978 27072 19984 27124
rect 20036 27112 20042 27124
rect 30558 27112 30564 27124
rect 20036 27084 30564 27112
rect 20036 27072 20042 27084
rect 30558 27072 30564 27084
rect 30616 27072 30622 27124
rect 35345 27115 35403 27121
rect 35345 27081 35357 27115
rect 35391 27112 35403 27115
rect 36446 27112 36452 27124
rect 35391 27084 36452 27112
rect 35391 27081 35403 27084
rect 35345 27075 35403 27081
rect 36446 27072 36452 27084
rect 36504 27072 36510 27124
rect 38933 27115 38991 27121
rect 38933 27081 38945 27115
rect 38979 27112 38991 27115
rect 40862 27112 40868 27124
rect 38979 27084 40868 27112
rect 38979 27081 38991 27084
rect 38933 27075 38991 27081
rect 40862 27072 40868 27084
rect 40920 27072 40926 27124
rect 41322 27112 41328 27124
rect 41283 27084 41328 27112
rect 41322 27072 41328 27084
rect 41380 27072 41386 27124
rect 44637 27115 44695 27121
rect 44637 27081 44649 27115
rect 44683 27112 44695 27115
rect 44910 27112 44916 27124
rect 44683 27084 44916 27112
rect 44683 27081 44695 27084
rect 44637 27075 44695 27081
rect 44910 27072 44916 27084
rect 44968 27072 44974 27124
rect 45002 27072 45008 27124
rect 45060 27112 45066 27124
rect 45097 27115 45155 27121
rect 45097 27112 45109 27115
rect 45060 27084 45109 27112
rect 45060 27072 45066 27084
rect 45097 27081 45109 27084
rect 45143 27081 45155 27115
rect 45097 27075 45155 27081
rect 50801 27115 50859 27121
rect 50801 27081 50813 27115
rect 50847 27112 50859 27115
rect 51258 27112 51264 27124
rect 50847 27084 51264 27112
rect 50847 27081 50859 27084
rect 50801 27075 50859 27081
rect 51258 27072 51264 27084
rect 51316 27072 51322 27124
rect 55861 27115 55919 27121
rect 55861 27081 55873 27115
rect 55907 27112 55919 27115
rect 56594 27112 56600 27124
rect 55907 27084 56600 27112
rect 55907 27081 55919 27084
rect 55861 27075 55919 27081
rect 56594 27072 56600 27084
rect 56652 27072 56658 27124
rect 58158 27112 58164 27124
rect 58119 27084 58164 27112
rect 58158 27072 58164 27084
rect 58216 27072 58222 27124
rect 8018 27053 8024 27056
rect 6932 27016 7880 27044
rect 8005 27047 8024 27053
rect 5629 26979 5687 26985
rect 5629 26945 5641 26979
rect 5675 26945 5687 26979
rect 6822 26976 6828 26988
rect 6783 26948 6828 26976
rect 5629 26939 5687 26945
rect 6822 26936 6828 26948
rect 6880 26936 6886 26988
rect 6932 26985 6960 27016
rect 8005 27013 8017 27047
rect 8005 27007 8024 27013
rect 8018 27004 8024 27007
rect 8076 27004 8082 27056
rect 8205 27047 8263 27053
rect 8205 27013 8217 27047
rect 8251 27013 8263 27047
rect 10042 27044 10048 27056
rect 10003 27016 10048 27044
rect 8205 27007 8263 27013
rect 6917 26979 6975 26985
rect 6917 26945 6929 26979
rect 6963 26945 6975 26979
rect 7098 26976 7104 26988
rect 7059 26948 7104 26976
rect 6917 26939 6975 26945
rect 7098 26936 7104 26948
rect 7156 26936 7162 26988
rect 7193 26979 7251 26985
rect 7193 26945 7205 26979
rect 7239 26976 7251 26979
rect 8110 26976 8116 26988
rect 7239 26948 8116 26976
rect 7239 26945 7251 26948
rect 7193 26939 7251 26945
rect 8110 26936 8116 26948
rect 8168 26936 8174 26988
rect 6270 26868 6276 26920
rect 6328 26908 6334 26920
rect 8220 26908 8248 27007
rect 10042 27004 10048 27016
rect 10100 27004 10106 27056
rect 10245 27047 10303 27053
rect 10245 27044 10257 27047
rect 10244 27013 10257 27044
rect 10291 27013 10303 27047
rect 10244 27007 10303 27013
rect 12069 27047 12127 27053
rect 12069 27013 12081 27047
rect 12115 27044 12127 27047
rect 12250 27044 12256 27056
rect 12115 27016 12256 27044
rect 12115 27013 12127 27016
rect 12069 27007 12127 27013
rect 9766 26936 9772 26988
rect 9824 26976 9830 26988
rect 10244 26976 10272 27007
rect 12250 27004 12256 27016
rect 12308 27004 12314 27056
rect 13262 27004 13268 27056
rect 13320 27044 13326 27056
rect 13725 27047 13783 27053
rect 13725 27044 13737 27047
rect 13320 27016 13737 27044
rect 13320 27004 13326 27016
rect 13725 27013 13737 27016
rect 13771 27013 13783 27047
rect 13725 27007 13783 27013
rect 14001 27047 14059 27053
rect 14001 27013 14013 27047
rect 14047 27044 14059 27047
rect 15841 27047 15899 27053
rect 14047 27016 14872 27044
rect 14047 27013 14059 27016
rect 14001 27007 14059 27013
rect 11422 26976 11428 26988
rect 9824 26948 11428 26976
rect 9824 26936 9830 26948
rect 11422 26936 11428 26948
rect 11480 26936 11486 26988
rect 13597 26979 13655 26985
rect 13597 26976 13609 26979
rect 13582 26945 13609 26976
rect 13643 26945 13655 26979
rect 13582 26939 13655 26945
rect 13582 26920 13610 26939
rect 13814 26936 13820 26988
rect 13872 26976 13878 26988
rect 14458 26976 14464 26988
rect 13872 26948 13917 26976
rect 14419 26948 14464 26976
rect 13872 26936 13878 26948
rect 14458 26936 14464 26948
rect 14516 26936 14522 26988
rect 14550 26936 14556 26988
rect 14608 26976 14614 26988
rect 14844 26985 14872 27016
rect 15841 27013 15853 27047
rect 15887 27044 15899 27047
rect 16022 27044 16028 27056
rect 15887 27016 16028 27044
rect 15887 27013 15899 27016
rect 15841 27007 15899 27013
rect 16022 27004 16028 27016
rect 16080 27004 16086 27056
rect 18690 27004 18696 27056
rect 18748 27044 18754 27056
rect 24762 27044 24768 27056
rect 18748 27016 24768 27044
rect 18748 27004 18754 27016
rect 24762 27004 24768 27016
rect 24820 27004 24826 27056
rect 26234 27004 26240 27056
rect 26292 27044 26298 27056
rect 27249 27047 27307 27053
rect 27249 27044 27261 27047
rect 26292 27016 27261 27044
rect 26292 27004 26298 27016
rect 27249 27013 27261 27016
rect 27295 27013 27307 27047
rect 27430 27044 27436 27056
rect 27391 27016 27436 27044
rect 27249 27007 27307 27013
rect 27430 27004 27436 27016
rect 27488 27004 27494 27056
rect 28626 27004 28632 27056
rect 28684 27044 28690 27056
rect 29089 27047 29147 27053
rect 29089 27044 29101 27047
rect 28684 27016 29101 27044
rect 28684 27004 28690 27016
rect 29089 27013 29101 27016
rect 29135 27013 29147 27047
rect 29089 27007 29147 27013
rect 38194 27004 38200 27056
rect 38252 27044 38258 27056
rect 38749 27047 38807 27053
rect 38749 27044 38761 27047
rect 38252 27016 38761 27044
rect 38252 27004 38258 27016
rect 38749 27013 38761 27016
rect 38795 27013 38807 27047
rect 38749 27007 38807 27013
rect 39942 27004 39948 27056
rect 40000 27044 40006 27056
rect 40313 27047 40371 27053
rect 40313 27044 40325 27047
rect 40000 27016 40325 27044
rect 40000 27004 40006 27016
rect 40313 27013 40325 27016
rect 40359 27044 40371 27047
rect 40957 27047 41015 27053
rect 40957 27044 40969 27047
rect 40359 27016 40969 27044
rect 40359 27013 40371 27016
rect 40313 27007 40371 27013
rect 40957 27013 40969 27016
rect 41003 27013 41015 27047
rect 41157 27047 41215 27053
rect 41157 27044 41169 27047
rect 40957 27007 41015 27013
rect 41064 27016 41169 27044
rect 14737 26979 14795 26985
rect 14608 26948 14653 26976
rect 14608 26936 14614 26948
rect 14737 26945 14749 26979
rect 14783 26945 14795 26979
rect 14737 26939 14795 26945
rect 14829 26979 14887 26985
rect 14829 26945 14841 26979
rect 14875 26945 14887 26979
rect 14829 26939 14887 26945
rect 6328 26880 8248 26908
rect 6328 26868 6334 26880
rect 13538 26868 13544 26920
rect 13596 26880 13610 26920
rect 13909 26911 13967 26917
rect 13596 26868 13602 26880
rect 13909 26877 13921 26911
rect 13955 26908 13967 26911
rect 14274 26908 14280 26920
rect 13955 26880 14280 26908
rect 13955 26877 13967 26880
rect 13909 26871 13967 26877
rect 14274 26868 14280 26880
rect 14332 26868 14338 26920
rect 14642 26868 14648 26920
rect 14700 26908 14706 26920
rect 14752 26908 14780 26939
rect 14700 26880 14780 26908
rect 14844 26908 14872 26939
rect 14918 26936 14924 26988
rect 14976 26985 14982 26988
rect 14976 26979 15025 26985
rect 14976 26945 14979 26979
rect 15013 26976 15025 26979
rect 15657 26979 15715 26985
rect 15657 26976 15669 26979
rect 15013 26948 15669 26976
rect 15013 26945 15025 26948
rect 14976 26939 15025 26945
rect 15657 26945 15669 26948
rect 15703 26945 15715 26979
rect 15657 26939 15715 26945
rect 14976 26936 14982 26939
rect 16482 26936 16488 26988
rect 16540 26976 16546 26988
rect 20257 26979 20315 26985
rect 20257 26976 20269 26979
rect 16540 26948 20269 26976
rect 16540 26936 16546 26948
rect 20257 26945 20269 26948
rect 20303 26976 20315 26979
rect 20530 26976 20536 26988
rect 20303 26948 20536 26976
rect 20303 26945 20315 26948
rect 20257 26939 20315 26945
rect 20530 26936 20536 26948
rect 20588 26936 20594 26988
rect 22186 26936 22192 26988
rect 22244 26976 22250 26988
rect 22741 26979 22799 26985
rect 22741 26976 22753 26979
rect 22244 26948 22753 26976
rect 22244 26936 22250 26948
rect 22741 26945 22753 26948
rect 22787 26945 22799 26979
rect 22741 26939 22799 26945
rect 22830 26936 22836 26988
rect 22888 26976 22894 26988
rect 22925 26979 22983 26985
rect 22925 26976 22937 26979
rect 22888 26948 22937 26976
rect 22888 26936 22894 26948
rect 22925 26945 22937 26948
rect 22971 26976 22983 26979
rect 23658 26976 23664 26988
rect 22971 26948 23664 26976
rect 22971 26945 22983 26948
rect 22925 26939 22983 26945
rect 23658 26936 23664 26948
rect 23716 26936 23722 26988
rect 14844 26880 15056 26908
rect 14700 26868 14706 26880
rect 15028 26852 15056 26880
rect 15286 26868 15292 26920
rect 15344 26908 15350 26920
rect 20162 26908 20168 26920
rect 15344 26880 20168 26908
rect 15344 26868 15350 26880
rect 20162 26868 20168 26880
rect 20220 26868 20226 26920
rect 20346 26908 20352 26920
rect 20307 26880 20352 26908
rect 20346 26868 20352 26880
rect 20404 26868 20410 26920
rect 21174 26908 21180 26920
rect 20456 26880 21180 26908
rect 2041 26843 2099 26849
rect 2041 26809 2053 26843
rect 2087 26840 2099 26843
rect 5442 26840 5448 26852
rect 2087 26812 5448 26840
rect 2087 26809 2099 26812
rect 2041 26803 2099 26809
rect 5442 26800 5448 26812
rect 5500 26800 5506 26852
rect 11882 26840 11888 26852
rect 11795 26812 11888 26840
rect 11882 26800 11888 26812
rect 11940 26840 11946 26852
rect 11940 26812 14504 26840
rect 11940 26800 11946 26812
rect 6638 26732 6644 26784
rect 6696 26772 6702 26784
rect 8021 26775 8079 26781
rect 8021 26772 8033 26775
rect 6696 26744 8033 26772
rect 6696 26732 6702 26744
rect 8021 26741 8033 26744
rect 8067 26741 8079 26775
rect 8021 26735 8079 26741
rect 9858 26732 9864 26784
rect 9916 26772 9922 26784
rect 10229 26775 10287 26781
rect 10229 26772 10241 26775
rect 9916 26744 10241 26772
rect 9916 26732 9922 26744
rect 10229 26741 10241 26744
rect 10275 26741 10287 26775
rect 10229 26735 10287 26741
rect 10318 26732 10324 26784
rect 10376 26772 10382 26784
rect 10413 26775 10471 26781
rect 10413 26772 10425 26775
rect 10376 26744 10425 26772
rect 10376 26732 10382 26744
rect 10413 26741 10425 26744
rect 10459 26741 10471 26775
rect 14476 26772 14504 26812
rect 15010 26800 15016 26852
rect 15068 26800 15074 26852
rect 19242 26840 19248 26852
rect 17972 26812 19248 26840
rect 17972 26784 18000 26812
rect 19242 26800 19248 26812
rect 19300 26800 19306 26852
rect 17954 26772 17960 26784
rect 14476 26744 17960 26772
rect 10413 26735 10471 26741
rect 17954 26732 17960 26744
rect 18012 26732 18018 26784
rect 18414 26732 18420 26784
rect 18472 26772 18478 26784
rect 20456 26772 20484 26880
rect 21174 26868 21180 26880
rect 21232 26868 21238 26920
rect 21634 26868 21640 26920
rect 21692 26908 21698 26920
rect 26878 26908 26884 26920
rect 21692 26880 26884 26908
rect 21692 26868 21698 26880
rect 26878 26868 26884 26880
rect 26936 26868 26942 26920
rect 27448 26908 27476 27004
rect 28077 26979 28135 26985
rect 28077 26945 28089 26979
rect 28123 26976 28135 26979
rect 28534 26976 28540 26988
rect 28123 26948 28540 26976
rect 28123 26945 28135 26948
rect 28077 26939 28135 26945
rect 28534 26936 28540 26948
rect 28592 26936 28598 26988
rect 32858 26936 32864 26988
rect 32916 26976 32922 26988
rect 34977 26979 35035 26985
rect 34977 26976 34989 26979
rect 32916 26948 34989 26976
rect 32916 26936 32922 26948
rect 34977 26945 34989 26948
rect 35023 26976 35035 26979
rect 35342 26976 35348 26988
rect 35023 26948 35348 26976
rect 35023 26945 35035 26948
rect 34977 26939 35035 26945
rect 35342 26936 35348 26948
rect 35400 26936 35406 26988
rect 37642 26936 37648 26988
rect 37700 26976 37706 26988
rect 38102 26976 38108 26988
rect 37700 26948 38108 26976
rect 37700 26936 37706 26948
rect 38102 26936 38108 26948
rect 38160 26976 38166 26988
rect 38565 26979 38623 26985
rect 38565 26976 38577 26979
rect 38160 26948 38577 26976
rect 38160 26936 38166 26948
rect 38565 26945 38577 26948
rect 38611 26945 38623 26979
rect 40218 26976 40224 26988
rect 40179 26948 40224 26976
rect 38565 26939 38623 26945
rect 40218 26936 40224 26948
rect 40276 26936 40282 26988
rect 40494 26976 40500 26988
rect 40455 26948 40500 26976
rect 40494 26936 40500 26948
rect 40552 26976 40558 26988
rect 41064 26976 41092 27016
rect 41157 27013 41169 27016
rect 41203 27013 41215 27047
rect 51166 27044 51172 27056
rect 41157 27007 41215 27013
rect 50724 27016 51172 27044
rect 44266 26976 44272 26988
rect 40552 26948 41092 26976
rect 44227 26948 44272 26976
rect 40552 26936 40558 26948
rect 44266 26936 44272 26948
rect 44324 26976 44330 26988
rect 50724 26985 50752 27016
rect 51166 27004 51172 27016
rect 51224 27044 51230 27056
rect 51350 27044 51356 27056
rect 51224 27016 51356 27044
rect 51224 27004 51230 27016
rect 51350 27004 51356 27016
rect 51408 27004 51414 27056
rect 53745 27047 53803 27053
rect 53745 27013 53757 27047
rect 53791 27044 53803 27047
rect 55306 27044 55312 27056
rect 53791 27016 55312 27044
rect 53791 27013 53803 27016
rect 53745 27007 53803 27013
rect 55306 27004 55312 27016
rect 55364 27004 55370 27056
rect 45097 26979 45155 26985
rect 45097 26976 45109 26979
rect 44324 26948 45109 26976
rect 44324 26936 44330 26948
rect 45097 26945 45109 26948
rect 45143 26945 45155 26979
rect 45097 26939 45155 26945
rect 45281 26979 45339 26985
rect 45281 26945 45293 26979
rect 45327 26945 45339 26979
rect 45281 26939 45339 26945
rect 50709 26979 50767 26985
rect 50709 26945 50721 26979
rect 50755 26945 50767 26979
rect 50890 26976 50896 26988
rect 50851 26948 50896 26976
rect 50709 26939 50767 26945
rect 28353 26911 28411 26917
rect 28353 26908 28365 26911
rect 27448 26880 28365 26908
rect 28353 26877 28365 26880
rect 28399 26877 28411 26911
rect 30466 26908 30472 26920
rect 28353 26871 28411 26877
rect 28460 26880 30472 26908
rect 20714 26800 20720 26852
rect 20772 26840 20778 26852
rect 28460 26840 28488 26880
rect 30466 26868 30472 26880
rect 30524 26868 30530 26920
rect 34514 26868 34520 26920
rect 34572 26908 34578 26920
rect 34885 26911 34943 26917
rect 34885 26908 34897 26911
rect 34572 26880 34897 26908
rect 34572 26868 34578 26880
rect 34885 26877 34897 26880
rect 34931 26877 34943 26911
rect 44174 26908 44180 26920
rect 44135 26880 44180 26908
rect 34885 26871 34943 26877
rect 44174 26868 44180 26880
rect 44232 26908 44238 26920
rect 45296 26908 45324 26939
rect 50890 26936 50896 26948
rect 50948 26936 50954 26988
rect 53374 26976 53380 26988
rect 53335 26948 53380 26976
rect 53374 26936 53380 26948
rect 53432 26936 53438 26988
rect 53561 26979 53619 26985
rect 53561 26945 53573 26979
rect 53607 26976 53619 26979
rect 54018 26976 54024 26988
rect 53607 26948 54024 26976
rect 53607 26945 53619 26948
rect 53561 26939 53619 26945
rect 54018 26936 54024 26948
rect 54076 26976 54082 26988
rect 55122 26976 55128 26988
rect 54076 26948 55128 26976
rect 54076 26936 54082 26948
rect 55122 26936 55128 26948
rect 55180 26976 55186 26988
rect 55677 26979 55735 26985
rect 55677 26976 55689 26979
rect 55180 26948 55689 26976
rect 55180 26936 55186 26948
rect 55677 26945 55689 26948
rect 55723 26945 55735 26979
rect 55677 26939 55735 26945
rect 55950 26936 55956 26988
rect 56008 26976 56014 26988
rect 56962 26976 56968 26988
rect 56008 26948 56053 26976
rect 56923 26948 56968 26976
rect 56008 26936 56014 26948
rect 56962 26936 56968 26948
rect 57020 26936 57026 26988
rect 56870 26908 56876 26920
rect 44232 26880 45324 26908
rect 56831 26880 56876 26908
rect 44232 26868 44238 26880
rect 56870 26868 56876 26880
rect 56928 26868 56934 26920
rect 20772 26812 28488 26840
rect 28629 26843 28687 26849
rect 20772 26800 20778 26812
rect 28629 26809 28641 26843
rect 28675 26840 28687 26843
rect 29365 26843 29423 26849
rect 29365 26840 29377 26843
rect 28675 26812 29377 26840
rect 28675 26809 28687 26812
rect 28629 26803 28687 26809
rect 29365 26809 29377 26812
rect 29411 26809 29423 26843
rect 29365 26803 29423 26809
rect 40497 26843 40555 26849
rect 40497 26809 40509 26843
rect 40543 26840 40555 26843
rect 41046 26840 41052 26852
rect 40543 26812 41052 26840
rect 40543 26809 40555 26812
rect 40497 26803 40555 26809
rect 41046 26800 41052 26812
rect 41104 26800 41110 26852
rect 55677 26843 55735 26849
rect 55677 26809 55689 26843
rect 55723 26840 55735 26843
rect 55858 26840 55864 26852
rect 55723 26812 55864 26840
rect 55723 26809 55735 26812
rect 55677 26803 55735 26809
rect 55858 26800 55864 26812
rect 55916 26800 55922 26852
rect 20622 26772 20628 26784
rect 18472 26744 20484 26772
rect 20583 26744 20628 26772
rect 18472 26732 18478 26744
rect 20622 26732 20628 26744
rect 20680 26732 20686 26784
rect 20806 26732 20812 26784
rect 20864 26772 20870 26784
rect 21085 26775 21143 26781
rect 21085 26772 21097 26775
rect 20864 26744 21097 26772
rect 20864 26732 20870 26744
rect 21085 26741 21097 26744
rect 21131 26741 21143 26775
rect 21085 26735 21143 26741
rect 22833 26775 22891 26781
rect 22833 26741 22845 26775
rect 22879 26772 22891 26775
rect 23566 26772 23572 26784
rect 22879 26744 23572 26772
rect 22879 26741 22891 26744
rect 22833 26735 22891 26741
rect 23566 26732 23572 26744
rect 23624 26732 23630 26784
rect 27617 26775 27675 26781
rect 27617 26741 27629 26775
rect 27663 26772 27675 26775
rect 27890 26772 27896 26784
rect 27663 26744 27896 26772
rect 27663 26741 27675 26744
rect 27617 26735 27675 26741
rect 27890 26732 27896 26744
rect 27948 26732 27954 26784
rect 28074 26732 28080 26784
rect 28132 26772 28138 26784
rect 28169 26775 28227 26781
rect 28169 26772 28181 26775
rect 28132 26744 28181 26772
rect 28132 26732 28138 26744
rect 28169 26741 28181 26744
rect 28215 26741 28227 26775
rect 29546 26772 29552 26784
rect 29507 26744 29552 26772
rect 28169 26735 28227 26741
rect 29546 26732 29552 26744
rect 29604 26732 29610 26784
rect 33594 26732 33600 26784
rect 33652 26772 33658 26784
rect 34790 26772 34796 26784
rect 33652 26744 34796 26772
rect 33652 26732 33658 26744
rect 34790 26732 34796 26744
rect 34848 26732 34854 26784
rect 41138 26772 41144 26784
rect 41099 26744 41144 26772
rect 41138 26732 41144 26744
rect 41196 26732 41202 26784
rect 57333 26775 57391 26781
rect 57333 26741 57345 26775
rect 57379 26772 57391 26775
rect 57882 26772 57888 26784
rect 57379 26744 57888 26772
rect 57379 26741 57391 26744
rect 57333 26735 57391 26741
rect 57882 26732 57888 26744
rect 57940 26732 57946 26784
rect 1104 26682 58880 26704
rect 1104 26630 4214 26682
rect 4266 26630 4278 26682
rect 4330 26630 4342 26682
rect 4394 26630 4406 26682
rect 4458 26630 4470 26682
rect 4522 26630 34934 26682
rect 34986 26630 34998 26682
rect 35050 26630 35062 26682
rect 35114 26630 35126 26682
rect 35178 26630 35190 26682
rect 35242 26630 58880 26682
rect 1104 26608 58880 26630
rect 1673 26571 1731 26577
rect 1673 26537 1685 26571
rect 1719 26568 1731 26571
rect 1854 26568 1860 26580
rect 1719 26540 1860 26568
rect 1719 26537 1731 26540
rect 1673 26531 1731 26537
rect 1854 26528 1860 26540
rect 1912 26528 1918 26580
rect 3142 26528 3148 26580
rect 3200 26568 3206 26580
rect 3881 26571 3939 26577
rect 3881 26568 3893 26571
rect 3200 26540 3893 26568
rect 3200 26528 3206 26540
rect 3881 26537 3893 26540
rect 3927 26568 3939 26571
rect 4062 26568 4068 26580
rect 3927 26540 4068 26568
rect 3927 26537 3939 26540
rect 3881 26531 3939 26537
rect 4062 26528 4068 26540
rect 4120 26528 4126 26580
rect 6457 26571 6515 26577
rect 6457 26537 6469 26571
rect 6503 26568 6515 26571
rect 6822 26568 6828 26580
rect 6503 26540 6828 26568
rect 6503 26537 6515 26540
rect 6457 26531 6515 26537
rect 6822 26528 6828 26540
rect 6880 26528 6886 26580
rect 10689 26571 10747 26577
rect 10689 26537 10701 26571
rect 10735 26568 10747 26571
rect 10962 26568 10968 26580
rect 10735 26540 10968 26568
rect 10735 26537 10747 26540
rect 10689 26531 10747 26537
rect 10962 26528 10968 26540
rect 11020 26528 11026 26580
rect 13538 26528 13544 26580
rect 13596 26568 13602 26580
rect 14090 26568 14096 26580
rect 13596 26540 14096 26568
rect 13596 26528 13602 26540
rect 14090 26528 14096 26540
rect 14148 26528 14154 26580
rect 18138 26568 18144 26580
rect 17052 26540 18144 26568
rect 8018 26500 8024 26512
rect 6196 26472 8024 26500
rect 6196 26373 6224 26472
rect 8018 26460 8024 26472
rect 8076 26500 8082 26512
rect 15194 26500 15200 26512
rect 8076 26472 15200 26500
rect 8076 26460 8082 26472
rect 15194 26460 15200 26472
rect 15252 26460 15258 26512
rect 6638 26392 6644 26444
rect 6696 26432 6702 26444
rect 6917 26435 6975 26441
rect 6917 26432 6929 26435
rect 6696 26404 6929 26432
rect 6696 26392 6702 26404
rect 6917 26401 6929 26404
rect 6963 26401 6975 26435
rect 11882 26432 11888 26444
rect 6917 26395 6975 26401
rect 10428 26404 11888 26432
rect 6181 26367 6239 26373
rect 6181 26333 6193 26367
rect 6227 26333 6239 26367
rect 6181 26327 6239 26333
rect 6270 26324 6276 26376
rect 6328 26364 6334 26376
rect 6457 26367 6515 26373
rect 6328 26336 6373 26364
rect 6328 26324 6334 26336
rect 6457 26333 6469 26367
rect 6503 26364 6515 26367
rect 7193 26367 7251 26373
rect 7193 26364 7205 26367
rect 6503 26336 7205 26364
rect 6503 26333 6515 26336
rect 6457 26327 6515 26333
rect 7193 26333 7205 26336
rect 7239 26364 7251 26367
rect 8018 26364 8024 26376
rect 7239 26336 8024 26364
rect 7239 26333 7251 26336
rect 7193 26327 7251 26333
rect 8018 26324 8024 26336
rect 8076 26364 8082 26376
rect 9858 26364 9864 26376
rect 8076 26336 9864 26364
rect 8076 26324 8082 26336
rect 9858 26324 9864 26336
rect 9916 26324 9922 26376
rect 10134 26364 10140 26376
rect 10095 26336 10140 26364
rect 10134 26324 10140 26336
rect 10192 26324 10198 26376
rect 10229 26367 10287 26373
rect 10229 26333 10241 26367
rect 10275 26364 10287 26367
rect 10318 26364 10324 26376
rect 10275 26336 10324 26364
rect 10275 26333 10287 26336
rect 10229 26327 10287 26333
rect 10318 26324 10324 26336
rect 10376 26324 10382 26376
rect 10428 26373 10456 26404
rect 11882 26392 11888 26404
rect 11940 26392 11946 26444
rect 15010 26432 15016 26444
rect 14971 26404 15016 26432
rect 15010 26392 15016 26404
rect 15068 26392 15074 26444
rect 10413 26367 10471 26373
rect 10413 26333 10425 26367
rect 10459 26333 10471 26367
rect 10413 26327 10471 26333
rect 10505 26367 10563 26373
rect 10505 26333 10517 26367
rect 10551 26333 10563 26367
rect 16758 26364 16764 26376
rect 10505 26327 10563 26333
rect 11256 26336 16764 26364
rect 10520 26296 10548 26327
rect 11256 26308 11284 26336
rect 16758 26324 16764 26336
rect 16816 26364 16822 26376
rect 17052 26373 17080 26540
rect 18138 26528 18144 26540
rect 18196 26528 18202 26580
rect 18690 26568 18696 26580
rect 18651 26540 18696 26568
rect 18690 26528 18696 26540
rect 18748 26528 18754 26580
rect 19058 26528 19064 26580
rect 19116 26568 19122 26580
rect 19610 26568 19616 26580
rect 19116 26540 19616 26568
rect 19116 26528 19122 26540
rect 19610 26528 19616 26540
rect 19668 26528 19674 26580
rect 19889 26571 19947 26577
rect 19889 26537 19901 26571
rect 19935 26568 19947 26571
rect 19978 26568 19984 26580
rect 19935 26540 19984 26568
rect 19935 26537 19947 26540
rect 19889 26531 19947 26537
rect 19978 26528 19984 26540
rect 20036 26528 20042 26580
rect 21450 26528 21456 26580
rect 21508 26568 21514 26580
rect 24489 26571 24547 26577
rect 21508 26540 24440 26568
rect 21508 26528 21514 26540
rect 17589 26503 17647 26509
rect 17589 26469 17601 26503
rect 17635 26469 17647 26503
rect 17589 26463 17647 26469
rect 17604 26432 17632 26463
rect 17678 26460 17684 26512
rect 17736 26500 17742 26512
rect 21082 26500 21088 26512
rect 17736 26472 21088 26500
rect 17736 26460 17742 26472
rect 21082 26460 21088 26472
rect 21140 26460 21146 26512
rect 21177 26503 21235 26509
rect 21177 26469 21189 26503
rect 21223 26500 21235 26503
rect 21223 26472 22416 26500
rect 21223 26469 21235 26472
rect 21177 26463 21235 26469
rect 17604 26404 18828 26432
rect 17037 26367 17095 26373
rect 17037 26364 17049 26367
rect 16816 26336 17049 26364
rect 16816 26324 16822 26336
rect 17037 26333 17049 26336
rect 17083 26333 17095 26367
rect 17310 26364 17316 26376
rect 17271 26336 17316 26364
rect 17037 26327 17095 26333
rect 17310 26324 17316 26336
rect 17368 26324 17374 26376
rect 17405 26367 17463 26373
rect 17405 26333 17417 26367
rect 17451 26364 17463 26367
rect 17678 26364 17684 26376
rect 17451 26336 17684 26364
rect 17451 26333 17463 26336
rect 17405 26327 17463 26333
rect 17678 26324 17684 26336
rect 17736 26324 17742 26376
rect 17770 26324 17776 26376
rect 17828 26364 17834 26376
rect 18049 26367 18107 26373
rect 18049 26364 18061 26367
rect 17828 26336 18061 26364
rect 17828 26324 17834 26336
rect 18049 26333 18061 26336
rect 18095 26333 18107 26367
rect 18049 26327 18107 26333
rect 18138 26324 18144 26376
rect 18196 26364 18202 26376
rect 18414 26364 18420 26376
rect 18196 26336 18241 26364
rect 18375 26336 18420 26364
rect 18196 26324 18202 26336
rect 18414 26324 18420 26336
rect 18472 26324 18478 26376
rect 18555 26367 18613 26373
rect 18555 26333 18567 26367
rect 18601 26364 18613 26367
rect 18690 26364 18696 26376
rect 18601 26336 18696 26364
rect 18601 26333 18613 26336
rect 18555 26327 18613 26333
rect 18690 26324 18696 26336
rect 18748 26324 18754 26376
rect 18800 26364 18828 26404
rect 20622 26392 20628 26444
rect 20680 26432 20686 26444
rect 22388 26441 22416 26472
rect 22738 26460 22744 26512
rect 22796 26500 22802 26512
rect 22796 26472 24072 26500
rect 22796 26460 22802 26472
rect 21453 26435 21511 26441
rect 21453 26432 21465 26435
rect 20680 26404 21465 26432
rect 20680 26392 20686 26404
rect 21453 26401 21465 26404
rect 21499 26432 21511 26435
rect 22373 26435 22431 26441
rect 21499 26404 22094 26432
rect 21499 26401 21511 26404
rect 21453 26395 21511 26401
rect 19245 26367 19303 26373
rect 19245 26364 19257 26367
rect 18800 26336 19257 26364
rect 19245 26333 19257 26336
rect 19291 26333 19303 26367
rect 19245 26327 19303 26333
rect 19334 26324 19340 26376
rect 19392 26364 19398 26376
rect 19702 26364 19708 26376
rect 19392 26336 19437 26364
rect 19661 26336 19708 26364
rect 19392 26324 19398 26336
rect 19702 26324 19708 26336
rect 19760 26373 19766 26376
rect 19760 26367 19809 26373
rect 19760 26333 19763 26367
rect 19797 26364 19809 26367
rect 22066 26364 22094 26404
rect 22373 26401 22385 26435
rect 22419 26432 22431 26435
rect 22830 26432 22836 26444
rect 22419 26404 22836 26432
rect 22419 26401 22431 26404
rect 22373 26395 22431 26401
rect 22830 26392 22836 26404
rect 22888 26392 22894 26444
rect 23201 26435 23259 26441
rect 23201 26401 23213 26435
rect 23247 26432 23259 26435
rect 23382 26432 23388 26444
rect 23247 26404 23388 26432
rect 23247 26401 23259 26404
rect 23201 26395 23259 26401
rect 23382 26392 23388 26404
rect 23440 26392 23446 26444
rect 22186 26364 22192 26376
rect 19797 26336 21956 26364
rect 22066 26336 22192 26364
rect 19797 26333 19809 26336
rect 19760 26327 19809 26333
rect 19760 26324 19766 26327
rect 11238 26296 11244 26308
rect 10244 26268 10548 26296
rect 11199 26268 11244 26296
rect 10244 26240 10272 26268
rect 11238 26256 11244 26268
rect 11296 26256 11302 26308
rect 11422 26296 11428 26308
rect 11383 26268 11428 26296
rect 11422 26256 11428 26268
rect 11480 26256 11486 26308
rect 14829 26299 14887 26305
rect 14829 26265 14841 26299
rect 14875 26296 14887 26299
rect 15194 26296 15200 26308
rect 14875 26268 15200 26296
rect 14875 26265 14887 26268
rect 14829 26259 14887 26265
rect 15194 26256 15200 26268
rect 15252 26256 15258 26308
rect 17221 26299 17279 26305
rect 17221 26265 17233 26299
rect 17267 26265 17279 26299
rect 17221 26259 17279 26265
rect 18325 26299 18383 26305
rect 18325 26265 18337 26299
rect 18371 26265 18383 26299
rect 19521 26299 19579 26305
rect 19521 26296 19533 26299
rect 18325 26259 18383 26265
rect 18524 26268 19533 26296
rect 10226 26188 10232 26240
rect 10284 26188 10290 26240
rect 17236 26228 17264 26259
rect 17402 26228 17408 26240
rect 17236 26200 17408 26228
rect 17402 26188 17408 26200
rect 17460 26188 17466 26240
rect 18340 26228 18368 26259
rect 18524 26228 18552 26268
rect 19521 26265 19533 26268
rect 19567 26265 19579 26299
rect 19521 26259 19579 26265
rect 18340 26200 18552 26228
rect 19536 26228 19564 26259
rect 19610 26256 19616 26308
rect 19668 26296 19674 26308
rect 19668 26268 19713 26296
rect 19668 26256 19674 26268
rect 21928 26240 21956 26336
rect 22186 26324 22192 26336
rect 22244 26324 22250 26376
rect 23290 26364 23296 26376
rect 23251 26336 23296 26364
rect 23290 26324 23296 26336
rect 23348 26324 23354 26376
rect 23566 26364 23572 26376
rect 23527 26336 23572 26364
rect 23566 26324 23572 26336
rect 23624 26324 23630 26376
rect 23661 26367 23719 26373
rect 23661 26333 23673 26367
rect 23707 26364 23719 26367
rect 23934 26364 23940 26376
rect 23707 26336 23940 26364
rect 23707 26333 23719 26336
rect 23661 26327 23719 26333
rect 23934 26324 23940 26336
rect 23992 26324 23998 26376
rect 24044 26364 24072 26472
rect 24412 26432 24440 26540
rect 24489 26537 24501 26571
rect 24535 26568 24547 26571
rect 25130 26568 25136 26580
rect 24535 26540 25136 26568
rect 24535 26537 24547 26540
rect 24489 26531 24547 26537
rect 25130 26528 25136 26540
rect 25188 26528 25194 26580
rect 34149 26571 34207 26577
rect 34149 26537 34161 26571
rect 34195 26568 34207 26571
rect 34422 26568 34428 26580
rect 34195 26540 34428 26568
rect 34195 26537 34207 26540
rect 34149 26531 34207 26537
rect 34422 26528 34428 26540
rect 34480 26528 34486 26580
rect 34790 26568 34796 26580
rect 34751 26540 34796 26568
rect 34790 26528 34796 26540
rect 34848 26528 34854 26580
rect 35161 26571 35219 26577
rect 35161 26537 35173 26571
rect 35207 26568 35219 26571
rect 38194 26568 38200 26580
rect 35207 26540 38200 26568
rect 35207 26537 35219 26540
rect 35161 26531 35219 26537
rect 38194 26528 38200 26540
rect 38252 26528 38258 26580
rect 41417 26571 41475 26577
rect 41417 26537 41429 26571
rect 41463 26568 41475 26571
rect 44266 26568 44272 26580
rect 41463 26540 44272 26568
rect 41463 26537 41475 26540
rect 41417 26531 41475 26537
rect 44266 26528 44272 26540
rect 44324 26528 44330 26580
rect 50706 26568 50712 26580
rect 50667 26540 50712 26568
rect 50706 26528 50712 26540
rect 50764 26528 50770 26580
rect 53101 26571 53159 26577
rect 53101 26537 53113 26571
rect 53147 26568 53159 26571
rect 53374 26568 53380 26580
rect 53147 26540 53380 26568
rect 53147 26537 53159 26540
rect 53101 26531 53159 26537
rect 53374 26528 53380 26540
rect 53432 26528 53438 26580
rect 55766 26528 55772 26580
rect 55824 26568 55830 26580
rect 55953 26571 56011 26577
rect 55953 26568 55965 26571
rect 55824 26540 55965 26568
rect 55824 26528 55830 26540
rect 55953 26537 55965 26540
rect 55999 26537 56011 26571
rect 55953 26531 56011 26537
rect 29546 26460 29552 26512
rect 29604 26500 29610 26512
rect 43162 26500 43168 26512
rect 29604 26472 34468 26500
rect 29604 26460 29610 26472
rect 33686 26432 33692 26444
rect 24412 26404 31754 26432
rect 33647 26404 33692 26432
rect 24394 26364 24400 26376
rect 24044 26336 24400 26364
rect 24394 26324 24400 26336
rect 24452 26324 24458 26376
rect 24581 26367 24639 26373
rect 24581 26333 24593 26367
rect 24627 26333 24639 26367
rect 27890 26364 27896 26376
rect 27851 26336 27896 26364
rect 24581 26327 24639 26333
rect 24118 26256 24124 26308
rect 24176 26296 24182 26308
rect 24596 26296 24624 26327
rect 27890 26324 27896 26336
rect 27948 26324 27954 26376
rect 30558 26364 30564 26376
rect 30519 26336 30564 26364
rect 30558 26324 30564 26336
rect 30616 26324 30622 26376
rect 30742 26364 30748 26376
rect 30703 26336 30748 26364
rect 30742 26324 30748 26336
rect 30800 26324 30806 26376
rect 31726 26364 31754 26404
rect 33686 26392 33692 26404
rect 33744 26432 33750 26444
rect 34440 26432 34468 26472
rect 34900 26472 43168 26500
rect 34900 26432 34928 26472
rect 43162 26460 43168 26472
rect 43220 26460 43226 26512
rect 33744 26404 33916 26432
rect 34440 26404 34928 26432
rect 38473 26435 38531 26441
rect 33744 26392 33750 26404
rect 33134 26364 33140 26376
rect 31726 26336 33140 26364
rect 33134 26324 33140 26336
rect 33192 26324 33198 26376
rect 33594 26324 33600 26376
rect 33652 26364 33658 26376
rect 33781 26367 33839 26373
rect 33781 26364 33793 26367
rect 33652 26336 33793 26364
rect 33652 26324 33658 26336
rect 33781 26333 33793 26336
rect 33827 26333 33839 26367
rect 33888 26364 33916 26404
rect 38473 26401 38485 26435
rect 38519 26432 38531 26435
rect 40494 26432 40500 26444
rect 38519 26404 40500 26432
rect 38519 26401 38531 26404
rect 38473 26395 38531 26401
rect 40494 26392 40500 26404
rect 40552 26432 40558 26444
rect 41233 26435 41291 26441
rect 41233 26432 41245 26435
rect 40552 26404 41245 26432
rect 40552 26392 40558 26404
rect 41233 26401 41245 26404
rect 41279 26401 41291 26435
rect 41233 26395 41291 26401
rect 49970 26392 49976 26444
rect 50028 26432 50034 26444
rect 50249 26435 50307 26441
rect 50249 26432 50261 26435
rect 50028 26404 50261 26432
rect 50028 26392 50034 26404
rect 50249 26401 50261 26404
rect 50295 26432 50307 26435
rect 50890 26432 50896 26444
rect 50295 26404 50896 26432
rect 50295 26401 50307 26404
rect 50249 26395 50307 26401
rect 50890 26392 50896 26404
rect 50948 26432 50954 26444
rect 50948 26404 51074 26432
rect 50948 26392 50954 26404
rect 34701 26367 34759 26373
rect 34701 26364 34713 26367
rect 33888 26336 34713 26364
rect 33781 26327 33839 26333
rect 34701 26333 34713 26336
rect 34747 26333 34759 26367
rect 34701 26327 34759 26333
rect 37185 26367 37243 26373
rect 37185 26333 37197 26367
rect 37231 26333 37243 26367
rect 37185 26327 37243 26333
rect 37369 26367 37427 26373
rect 37369 26333 37381 26367
rect 37415 26364 37427 26367
rect 37458 26364 37464 26376
rect 37415 26336 37464 26364
rect 37415 26333 37427 26336
rect 37369 26327 37427 26333
rect 25041 26299 25099 26305
rect 25041 26296 25053 26299
rect 24176 26268 25053 26296
rect 24176 26256 24182 26268
rect 25041 26265 25053 26268
rect 25087 26265 25099 26299
rect 25041 26259 25099 26265
rect 31573 26299 31631 26305
rect 31573 26265 31585 26299
rect 31619 26296 31631 26299
rect 37200 26296 37228 26327
rect 37458 26324 37464 26336
rect 37516 26324 37522 26376
rect 37737 26367 37795 26373
rect 37737 26333 37749 26367
rect 37783 26364 37795 26367
rect 38102 26364 38108 26376
rect 37783 26336 38108 26364
rect 37783 26333 37795 26336
rect 37737 26327 37795 26333
rect 38102 26324 38108 26336
rect 38160 26364 38166 26376
rect 38381 26367 38439 26373
rect 38381 26364 38393 26367
rect 38160 26336 38393 26364
rect 38160 26324 38166 26336
rect 38381 26333 38393 26336
rect 38427 26333 38439 26367
rect 38381 26327 38439 26333
rect 38565 26367 38623 26373
rect 38565 26333 38577 26367
rect 38611 26364 38623 26367
rect 38746 26364 38752 26376
rect 38611 26336 38752 26364
rect 38611 26333 38623 26336
rect 38565 26327 38623 26333
rect 38746 26324 38752 26336
rect 38804 26324 38810 26376
rect 40218 26324 40224 26376
rect 40276 26364 40282 26376
rect 41138 26364 41144 26376
rect 40276 26336 41144 26364
rect 40276 26324 40282 26336
rect 41138 26324 41144 26336
rect 41196 26324 41202 26376
rect 50062 26324 50068 26376
rect 50120 26364 50126 26376
rect 50341 26367 50399 26373
rect 50341 26364 50353 26367
rect 50120 26336 50353 26364
rect 50120 26324 50126 26336
rect 50341 26333 50353 26336
rect 50387 26333 50399 26367
rect 51046 26364 51074 26404
rect 51169 26367 51227 26373
rect 51169 26364 51181 26367
rect 51046 26336 51181 26364
rect 50341 26327 50399 26333
rect 51169 26333 51181 26336
rect 51215 26333 51227 26367
rect 51350 26364 51356 26376
rect 51311 26336 51356 26364
rect 51169 26327 51227 26333
rect 51350 26324 51356 26336
rect 51408 26324 51414 26376
rect 52822 26364 52828 26376
rect 52783 26336 52828 26364
rect 52822 26324 52828 26336
rect 52880 26324 52886 26376
rect 55950 26364 55956 26376
rect 55911 26336 55956 26364
rect 55950 26324 55956 26336
rect 56008 26324 56014 26376
rect 56137 26367 56195 26373
rect 56137 26333 56149 26367
rect 56183 26364 56195 26367
rect 56594 26364 56600 26376
rect 56183 26336 56600 26364
rect 56183 26333 56195 26336
rect 56137 26327 56195 26333
rect 56594 26324 56600 26336
rect 56652 26324 56658 26376
rect 37274 26296 37280 26308
rect 31619 26268 37280 26296
rect 31619 26265 31631 26268
rect 31573 26259 31631 26265
rect 37274 26256 37280 26268
rect 37332 26256 37338 26308
rect 37645 26299 37703 26305
rect 37645 26265 37657 26299
rect 37691 26296 37703 26299
rect 45094 26296 45100 26308
rect 37691 26268 45100 26296
rect 37691 26265 37703 26268
rect 37645 26259 37703 26265
rect 45094 26256 45100 26268
rect 45152 26256 45158 26308
rect 51537 26299 51595 26305
rect 51537 26265 51549 26299
rect 51583 26296 51595 26299
rect 52270 26296 52276 26308
rect 51583 26268 52276 26296
rect 51583 26265 51595 26268
rect 51537 26259 51595 26265
rect 52270 26256 52276 26268
rect 52328 26256 52334 26308
rect 52365 26299 52423 26305
rect 52365 26265 52377 26299
rect 52411 26296 52423 26299
rect 52454 26296 52460 26308
rect 52411 26268 52460 26296
rect 52411 26265 52423 26268
rect 52365 26259 52423 26265
rect 52454 26256 52460 26268
rect 52512 26296 52518 26308
rect 53101 26299 53159 26305
rect 53101 26296 53113 26299
rect 52512 26268 53113 26296
rect 52512 26256 52518 26268
rect 53101 26265 53113 26268
rect 53147 26296 53159 26299
rect 53561 26299 53619 26305
rect 53561 26296 53573 26299
rect 53147 26268 53573 26296
rect 53147 26265 53159 26268
rect 53101 26259 53159 26265
rect 53561 26265 53573 26268
rect 53607 26296 53619 26299
rect 53650 26296 53656 26308
rect 53607 26268 53656 26296
rect 53607 26265 53619 26268
rect 53561 26259 53619 26265
rect 53650 26256 53656 26268
rect 53708 26256 53714 26308
rect 20622 26228 20628 26240
rect 19536 26200 20628 26228
rect 20622 26188 20628 26200
rect 20680 26188 20686 26240
rect 20993 26231 21051 26237
rect 20993 26197 21005 26231
rect 21039 26228 21051 26231
rect 21082 26228 21088 26240
rect 21039 26200 21088 26228
rect 21039 26197 21051 26200
rect 20993 26191 21051 26197
rect 21082 26188 21088 26200
rect 21140 26188 21146 26240
rect 21910 26188 21916 26240
rect 21968 26228 21974 26240
rect 22005 26231 22063 26237
rect 22005 26228 22017 26231
rect 21968 26200 22017 26228
rect 21968 26188 21974 26200
rect 22005 26197 22017 26200
rect 22051 26197 22063 26231
rect 22005 26191 22063 26197
rect 23845 26231 23903 26237
rect 23845 26197 23857 26231
rect 23891 26228 23903 26231
rect 24026 26228 24032 26240
rect 23891 26200 24032 26228
rect 23891 26197 23903 26200
rect 23845 26191 23903 26197
rect 24026 26188 24032 26200
rect 24084 26188 24090 26240
rect 27985 26231 28043 26237
rect 27985 26197 27997 26231
rect 28031 26228 28043 26231
rect 28074 26228 28080 26240
rect 28031 26200 28080 26228
rect 28031 26197 28043 26200
rect 27985 26191 28043 26197
rect 28074 26188 28080 26200
rect 28132 26188 28138 26240
rect 39942 26188 39948 26240
rect 40000 26228 40006 26240
rect 40773 26231 40831 26237
rect 40773 26228 40785 26231
rect 40000 26200 40785 26228
rect 40000 26188 40006 26200
rect 40773 26197 40785 26200
rect 40819 26197 40831 26231
rect 40773 26191 40831 26197
rect 52917 26231 52975 26237
rect 52917 26197 52929 26231
rect 52963 26228 52975 26231
rect 53190 26228 53196 26240
rect 52963 26200 53196 26228
rect 52963 26197 52975 26200
rect 52917 26191 52975 26197
rect 53190 26188 53196 26200
rect 53248 26188 53254 26240
rect 1104 26138 58880 26160
rect 1104 26086 19574 26138
rect 19626 26086 19638 26138
rect 19690 26086 19702 26138
rect 19754 26086 19766 26138
rect 19818 26086 19830 26138
rect 19882 26086 50294 26138
rect 50346 26086 50358 26138
rect 50410 26086 50422 26138
rect 50474 26086 50486 26138
rect 50538 26086 50550 26138
rect 50602 26086 58880 26138
rect 1104 26064 58880 26086
rect 2774 25984 2780 26036
rect 2832 26024 2838 26036
rect 4062 26024 4068 26036
rect 2832 25996 4068 26024
rect 2832 25984 2838 25996
rect 4062 25984 4068 25996
rect 4120 26024 4126 26036
rect 4120 25996 4292 26024
rect 4120 25984 4126 25996
rect 4264 25965 4292 25996
rect 6270 25984 6276 26036
rect 6328 26024 6334 26036
rect 6457 26027 6515 26033
rect 6457 26024 6469 26027
rect 6328 25996 6469 26024
rect 6328 25984 6334 25996
rect 6457 25993 6469 25996
rect 6503 25993 6515 26027
rect 9950 26024 9956 26036
rect 9911 25996 9956 26024
rect 6457 25987 6515 25993
rect 9950 25984 9956 25996
rect 10008 25984 10014 26036
rect 10594 26024 10600 26036
rect 10060 25996 10600 26024
rect 4249 25959 4307 25965
rect 4249 25925 4261 25959
rect 4295 25925 4307 25959
rect 10060 25956 10088 25996
rect 10594 25984 10600 25996
rect 10652 25984 10658 26036
rect 10686 25984 10692 26036
rect 10744 26024 10750 26036
rect 13817 26027 13875 26033
rect 10744 25996 13768 26024
rect 10744 25984 10750 25996
rect 11238 25956 11244 25968
rect 4249 25919 4307 25925
rect 9232 25928 10088 25956
rect 10152 25928 11244 25956
rect 3142 25888 3148 25900
rect 3103 25860 3148 25888
rect 3142 25848 3148 25860
rect 3200 25848 3206 25900
rect 5813 25891 5871 25897
rect 5813 25857 5825 25891
rect 5859 25888 5871 25891
rect 6641 25891 6699 25897
rect 6641 25888 6653 25891
rect 5859 25860 6653 25888
rect 5859 25857 5871 25860
rect 5813 25851 5871 25857
rect 6641 25857 6653 25860
rect 6687 25888 6699 25891
rect 6914 25888 6920 25900
rect 6687 25860 6920 25888
rect 6687 25857 6699 25860
rect 6641 25851 6699 25857
rect 6914 25848 6920 25860
rect 6972 25848 6978 25900
rect 9232 25897 9260 25928
rect 8113 25891 8171 25897
rect 8113 25888 8125 25891
rect 7760 25860 8125 25888
rect 3053 25823 3111 25829
rect 3053 25789 3065 25823
rect 3099 25789 3111 25823
rect 3053 25783 3111 25789
rect 3068 25752 3096 25783
rect 3142 25752 3148 25764
rect 3068 25724 3148 25752
rect 3142 25712 3148 25724
rect 3200 25712 3206 25764
rect 3970 25752 3976 25764
rect 3931 25724 3976 25752
rect 3970 25712 3976 25724
rect 4028 25712 4034 25764
rect 6638 25712 6644 25764
rect 6696 25752 6702 25764
rect 7760 25752 7788 25860
rect 8113 25857 8125 25860
rect 8159 25857 8171 25891
rect 8113 25851 8171 25857
rect 9217 25891 9275 25897
rect 9217 25857 9229 25891
rect 9263 25857 9275 25891
rect 9398 25888 9404 25900
rect 9359 25860 9404 25888
rect 9217 25851 9275 25857
rect 7837 25823 7895 25829
rect 7837 25789 7849 25823
rect 7883 25820 7895 25823
rect 9232 25820 9260 25851
rect 9398 25848 9404 25860
rect 9456 25848 9462 25900
rect 9493 25891 9551 25897
rect 9493 25857 9505 25891
rect 9539 25888 9551 25891
rect 9766 25888 9772 25900
rect 9539 25860 9772 25888
rect 9539 25857 9551 25860
rect 9493 25851 9551 25857
rect 9766 25848 9772 25860
rect 9824 25848 9830 25900
rect 10152 25897 10180 25928
rect 11238 25916 11244 25928
rect 11296 25916 11302 25968
rect 12986 25916 12992 25968
rect 13044 25956 13050 25968
rect 13541 25959 13599 25965
rect 13541 25956 13553 25959
rect 13044 25928 13553 25956
rect 13044 25916 13050 25928
rect 13541 25925 13553 25928
rect 13587 25925 13599 25959
rect 13740 25956 13768 25996
rect 13817 25993 13829 26027
rect 13863 26024 13875 26027
rect 14458 26024 14464 26036
rect 13863 25996 14464 26024
rect 13863 25993 13875 25996
rect 13817 25987 13875 25993
rect 14458 25984 14464 25996
rect 14516 25984 14522 26036
rect 17770 26024 17776 26036
rect 17731 25996 17776 26024
rect 17770 25984 17776 25996
rect 17828 25984 17834 26036
rect 18230 25984 18236 26036
rect 18288 26024 18294 26036
rect 18325 26027 18383 26033
rect 18325 26024 18337 26027
rect 18288 25996 18337 26024
rect 18288 25984 18294 25996
rect 18325 25993 18337 25996
rect 18371 26024 18383 26027
rect 19058 26024 19064 26036
rect 18371 25996 19064 26024
rect 18371 25993 18383 25996
rect 18325 25987 18383 25993
rect 19058 25984 19064 25996
rect 19116 25984 19122 26036
rect 20622 25984 20628 26036
rect 20680 26024 20686 26036
rect 22005 26027 22063 26033
rect 22005 26024 22017 26027
rect 20680 25996 22017 26024
rect 20680 25984 20686 25996
rect 22005 25993 22017 25996
rect 22051 25993 22063 26027
rect 22005 25987 22063 25993
rect 27893 26027 27951 26033
rect 27893 25993 27905 26027
rect 27939 26024 27951 26027
rect 28166 26024 28172 26036
rect 27939 25996 28172 26024
rect 27939 25993 27951 25996
rect 27893 25987 27951 25993
rect 28166 25984 28172 25996
rect 28224 25984 28230 26036
rect 38746 26024 38752 26036
rect 38707 25996 38752 26024
rect 38746 25984 38752 25996
rect 38804 25984 38810 26036
rect 43993 26027 44051 26033
rect 43993 25993 44005 26027
rect 44039 26024 44051 26027
rect 44174 26024 44180 26036
rect 44039 25996 44180 26024
rect 44039 25993 44051 25996
rect 43993 25987 44051 25993
rect 44174 25984 44180 25996
rect 44232 25984 44238 26036
rect 47946 26024 47952 26036
rect 47907 25996 47952 26024
rect 47946 25984 47952 25996
rect 48004 25984 48010 26036
rect 49326 26024 49332 26036
rect 48700 25996 49332 26024
rect 13740 25928 14412 25956
rect 13541 25919 13599 25925
rect 10137 25891 10195 25897
rect 10137 25857 10149 25891
rect 10183 25857 10195 25891
rect 10137 25851 10195 25857
rect 10226 25848 10232 25900
rect 10284 25888 10290 25900
rect 10413 25891 10471 25897
rect 10284 25860 10377 25888
rect 10284 25848 10290 25860
rect 10413 25857 10425 25891
rect 10459 25857 10471 25891
rect 10413 25851 10471 25857
rect 10505 25891 10563 25897
rect 10505 25857 10517 25891
rect 10551 25857 10563 25891
rect 10505 25851 10563 25857
rect 7883 25792 9260 25820
rect 7883 25789 7895 25792
rect 7837 25783 7895 25789
rect 9674 25780 9680 25832
rect 9732 25820 9738 25832
rect 10244 25820 10272 25848
rect 9732 25792 10272 25820
rect 9732 25780 9738 25792
rect 10318 25780 10324 25832
rect 10376 25820 10382 25832
rect 10428 25820 10456 25851
rect 10376 25792 10456 25820
rect 10520 25820 10548 25851
rect 10594 25848 10600 25900
rect 10652 25888 10658 25900
rect 11517 25891 11575 25897
rect 11517 25888 11529 25891
rect 10652 25860 11529 25888
rect 10652 25848 10658 25860
rect 11517 25857 11529 25860
rect 11563 25857 11575 25891
rect 11517 25851 11575 25857
rect 11701 25891 11759 25897
rect 11701 25857 11713 25891
rect 11747 25857 11759 25891
rect 11701 25851 11759 25857
rect 10520 25792 11560 25820
rect 10376 25780 10382 25792
rect 6696 25724 7788 25752
rect 9217 25755 9275 25761
rect 6696 25712 6702 25724
rect 9217 25721 9229 25755
rect 9263 25752 9275 25755
rect 10134 25752 10140 25764
rect 9263 25724 10140 25752
rect 9263 25721 9275 25724
rect 9217 25715 9275 25721
rect 10134 25712 10140 25724
rect 10192 25712 10198 25764
rect 11532 25761 11560 25792
rect 11517 25755 11575 25761
rect 11517 25721 11529 25755
rect 11563 25721 11575 25755
rect 11517 25715 11575 25721
rect 3418 25644 3424 25696
rect 3476 25684 3482 25696
rect 3789 25687 3847 25693
rect 3789 25684 3801 25687
rect 3476 25656 3801 25684
rect 3476 25644 3482 25656
rect 3789 25653 3801 25656
rect 3835 25653 3847 25687
rect 3789 25647 3847 25653
rect 9398 25644 9404 25696
rect 9456 25684 9462 25696
rect 11054 25684 11060 25696
rect 9456 25656 11060 25684
rect 9456 25644 9462 25656
rect 11054 25644 11060 25656
rect 11112 25684 11118 25696
rect 11716 25684 11744 25851
rect 11790 25848 11796 25900
rect 11848 25888 11854 25900
rect 13262 25888 13268 25900
rect 11848 25860 11893 25888
rect 13223 25860 13268 25888
rect 11848 25848 11854 25860
rect 13262 25848 13268 25860
rect 13320 25848 13326 25900
rect 13449 25891 13507 25897
rect 13449 25857 13461 25891
rect 13495 25857 13507 25891
rect 13630 25888 13636 25900
rect 13591 25860 13636 25888
rect 13449 25851 13507 25857
rect 13170 25780 13176 25832
rect 13228 25820 13234 25832
rect 13464 25820 13492 25851
rect 13630 25848 13636 25860
rect 13688 25888 13694 25900
rect 14277 25891 14335 25897
rect 14277 25888 14289 25891
rect 13688 25860 14289 25888
rect 13688 25848 13694 25860
rect 14277 25857 14289 25860
rect 14323 25857 14335 25891
rect 14384 25888 14412 25928
rect 15194 25916 15200 25968
rect 15252 25956 15258 25968
rect 17497 25959 17555 25965
rect 17497 25956 17509 25959
rect 15252 25928 17509 25956
rect 15252 25916 15258 25928
rect 17497 25925 17509 25928
rect 17543 25925 17555 25959
rect 17497 25919 17555 25925
rect 18138 25916 18144 25968
rect 18196 25956 18202 25968
rect 18969 25959 19027 25965
rect 18969 25956 18981 25959
rect 18196 25928 18981 25956
rect 18196 25916 18202 25928
rect 18969 25925 18981 25928
rect 19015 25925 19027 25959
rect 21082 25956 21088 25968
rect 21043 25928 21088 25956
rect 18969 25919 19027 25925
rect 21082 25916 21088 25928
rect 21140 25916 21146 25968
rect 21726 25916 21732 25968
rect 21784 25956 21790 25968
rect 24305 25959 24363 25965
rect 24305 25956 24317 25959
rect 21784 25928 24317 25956
rect 21784 25916 21790 25928
rect 24305 25925 24317 25928
rect 24351 25925 24363 25959
rect 24305 25919 24363 25925
rect 24397 25959 24455 25965
rect 24397 25925 24409 25959
rect 24443 25956 24455 25959
rect 24443 25928 24717 25956
rect 24443 25925 24455 25928
rect 24397 25919 24455 25925
rect 14734 25888 14740 25900
rect 14384 25860 14740 25888
rect 14277 25851 14335 25857
rect 14734 25848 14740 25860
rect 14792 25888 14798 25900
rect 17218 25888 17224 25900
rect 14792 25860 17224 25888
rect 14792 25848 14798 25860
rect 17218 25848 17224 25860
rect 17276 25848 17282 25900
rect 17402 25888 17408 25900
rect 17363 25860 17408 25888
rect 17402 25848 17408 25860
rect 17460 25848 17466 25900
rect 17589 25891 17647 25897
rect 17589 25857 17601 25891
rect 17635 25888 17647 25891
rect 17678 25888 17684 25900
rect 17635 25860 17684 25888
rect 17635 25857 17647 25860
rect 17589 25851 17647 25857
rect 17678 25848 17684 25860
rect 17736 25848 17742 25900
rect 22189 25891 22247 25897
rect 22189 25857 22201 25891
rect 22235 25857 22247 25891
rect 22189 25851 22247 25857
rect 13722 25820 13728 25832
rect 13228 25792 13728 25820
rect 13228 25780 13234 25792
rect 13722 25780 13728 25792
rect 13780 25780 13786 25832
rect 22204 25820 22232 25851
rect 22278 25848 22284 25900
rect 22336 25888 22342 25900
rect 24026 25888 24032 25900
rect 22336 25860 22381 25888
rect 23987 25860 24032 25888
rect 22336 25848 22342 25860
rect 24026 25848 24032 25860
rect 24084 25848 24090 25900
rect 24177 25891 24235 25897
rect 24177 25857 24189 25891
rect 24223 25888 24235 25891
rect 24223 25857 24256 25888
rect 24177 25851 24256 25857
rect 22922 25820 22928 25832
rect 22204 25792 22928 25820
rect 22922 25780 22928 25792
rect 22980 25780 22986 25832
rect 24228 25820 24256 25851
rect 24486 25848 24492 25900
rect 24544 25897 24550 25900
rect 24544 25888 24552 25897
rect 24689 25888 24717 25928
rect 24762 25916 24768 25968
rect 24820 25956 24826 25968
rect 48700 25965 48728 25996
rect 49326 25984 49332 25996
rect 49384 25984 49390 26036
rect 50062 26024 50068 26036
rect 50023 25996 50068 26024
rect 50062 25984 50068 25996
rect 50120 25984 50126 26036
rect 52822 25984 52828 26036
rect 52880 25984 52886 26036
rect 53190 26024 53196 26036
rect 53151 25996 53196 26024
rect 53190 25984 53196 25996
rect 53248 25984 53254 26036
rect 53853 26027 53911 26033
rect 53853 26024 53865 26027
rect 53300 25996 53865 26024
rect 47765 25959 47823 25965
rect 47765 25956 47777 25959
rect 24820 25928 30420 25956
rect 24820 25916 24826 25928
rect 24946 25888 24952 25900
rect 24544 25860 24589 25888
rect 24689 25860 24952 25888
rect 24544 25851 24552 25860
rect 24544 25848 24550 25851
rect 24946 25848 24952 25860
rect 25004 25848 25010 25900
rect 28074 25888 28080 25900
rect 28035 25860 28080 25888
rect 28074 25848 28080 25860
rect 28132 25848 28138 25900
rect 24578 25820 24584 25832
rect 24228 25792 24584 25820
rect 24578 25780 24584 25792
rect 24636 25780 24642 25832
rect 28258 25820 28264 25832
rect 28219 25792 28264 25820
rect 28258 25780 28264 25792
rect 28316 25780 28322 25832
rect 30392 25829 30420 25928
rect 47044 25928 47777 25956
rect 47044 25900 47072 25928
rect 47765 25925 47777 25928
rect 47811 25925 47823 25959
rect 47765 25919 47823 25925
rect 48685 25959 48743 25965
rect 48685 25925 48697 25959
rect 48731 25925 48743 25959
rect 52840 25956 52868 25984
rect 53300 25956 53328 25996
rect 53853 25993 53865 25996
rect 53899 25993 53911 26027
rect 54018 26024 54024 26036
rect 53979 25996 54024 26024
rect 53853 25987 53911 25993
rect 54018 25984 54024 25996
rect 54076 25984 54082 26036
rect 55950 25984 55956 26036
rect 56008 26024 56014 26036
rect 56229 26027 56287 26033
rect 56229 26024 56241 26027
rect 56008 25996 56241 26024
rect 56008 25984 56014 25996
rect 56229 25993 56241 25996
rect 56275 25993 56287 26027
rect 56229 25987 56287 25993
rect 53650 25956 53656 25968
rect 48685 25919 48743 25925
rect 48792 25928 50200 25956
rect 52840 25928 53328 25956
rect 53611 25928 53656 25956
rect 30469 25891 30527 25897
rect 30469 25857 30481 25891
rect 30515 25888 30527 25891
rect 30742 25888 30748 25900
rect 30515 25860 30748 25888
rect 30515 25857 30527 25860
rect 30469 25851 30527 25857
rect 30742 25848 30748 25860
rect 30800 25848 30806 25900
rect 37458 25888 37464 25900
rect 37419 25860 37464 25888
rect 37458 25848 37464 25860
rect 37516 25848 37522 25900
rect 43625 25891 43683 25897
rect 43625 25857 43637 25891
rect 43671 25888 43683 25891
rect 43806 25888 43812 25900
rect 43671 25860 43812 25888
rect 43671 25857 43683 25860
rect 43625 25851 43683 25857
rect 43806 25848 43812 25860
rect 43864 25848 43870 25900
rect 46842 25888 46848 25900
rect 46803 25860 46848 25888
rect 46842 25848 46848 25860
rect 46900 25848 46906 25900
rect 47026 25888 47032 25900
rect 46987 25860 47032 25888
rect 47026 25848 47032 25860
rect 47084 25848 47090 25900
rect 47578 25888 47584 25900
rect 47539 25860 47584 25888
rect 47578 25848 47584 25860
rect 47636 25848 47642 25900
rect 48792 25888 48820 25928
rect 50172 25900 50200 25928
rect 53650 25916 53656 25928
rect 53708 25916 53714 25968
rect 48332 25874 48820 25888
rect 49973 25891 50031 25897
rect 48332 25860 48806 25874
rect 30377 25823 30435 25829
rect 30377 25789 30389 25823
rect 30423 25789 30435 25823
rect 30377 25783 30435 25789
rect 37274 25780 37280 25832
rect 37332 25820 37338 25832
rect 37369 25823 37427 25829
rect 37369 25820 37381 25823
rect 37332 25792 37381 25820
rect 37332 25780 37338 25792
rect 37369 25789 37381 25792
rect 37415 25789 37427 25823
rect 37369 25783 37427 25789
rect 37829 25823 37887 25829
rect 37829 25789 37841 25823
rect 37875 25820 37887 25823
rect 38010 25820 38016 25832
rect 37875 25792 38016 25820
rect 37875 25789 37887 25792
rect 37829 25783 37887 25789
rect 38010 25780 38016 25792
rect 38068 25820 38074 25832
rect 38289 25823 38347 25829
rect 38289 25820 38301 25823
rect 38068 25792 38301 25820
rect 38068 25780 38074 25792
rect 38289 25789 38301 25792
rect 38335 25789 38347 25823
rect 43714 25820 43720 25832
rect 43675 25792 43720 25820
rect 38289 25783 38347 25789
rect 43714 25780 43720 25792
rect 43772 25780 43778 25832
rect 46937 25823 46995 25829
rect 46937 25789 46949 25823
rect 46983 25820 46995 25823
rect 48332 25820 48360 25860
rect 49973 25857 49985 25891
rect 50019 25857 50031 25891
rect 49973 25851 50031 25857
rect 49234 25820 49240 25832
rect 46983 25792 48360 25820
rect 49195 25792 49240 25820
rect 46983 25789 46995 25792
rect 46937 25783 46995 25789
rect 49234 25780 49240 25792
rect 49292 25820 49298 25832
rect 49988 25820 50016 25851
rect 50154 25848 50160 25900
rect 50212 25888 50218 25900
rect 50212 25860 50305 25888
rect 50212 25848 50218 25860
rect 52362 25848 52368 25900
rect 52420 25888 52426 25900
rect 52733 25891 52791 25897
rect 52733 25888 52745 25891
rect 52420 25860 52745 25888
rect 52420 25848 52426 25860
rect 52733 25857 52745 25860
rect 52779 25857 52791 25891
rect 52733 25851 52791 25857
rect 52825 25891 52883 25897
rect 52825 25857 52837 25891
rect 52871 25857 52883 25891
rect 52825 25851 52883 25857
rect 53009 25891 53067 25897
rect 53009 25857 53021 25891
rect 53055 25888 53067 25891
rect 53098 25888 53104 25900
rect 53055 25860 53104 25888
rect 53055 25857 53067 25860
rect 53009 25851 53067 25857
rect 49292 25792 50016 25820
rect 49292 25780 49298 25792
rect 52270 25780 52276 25832
rect 52328 25820 52334 25832
rect 52840 25820 52868 25851
rect 53098 25848 53104 25860
rect 53156 25848 53162 25900
rect 55861 25891 55919 25897
rect 55861 25857 55873 25891
rect 55907 25888 55919 25891
rect 55950 25888 55956 25900
rect 55907 25860 55956 25888
rect 55907 25857 55919 25860
rect 55861 25851 55919 25857
rect 55950 25848 55956 25860
rect 56008 25848 56014 25900
rect 52914 25820 52920 25832
rect 52328 25792 52920 25820
rect 52328 25780 52334 25792
rect 52914 25780 52920 25792
rect 52972 25780 52978 25832
rect 55766 25820 55772 25832
rect 55727 25792 55772 25820
rect 55766 25780 55772 25792
rect 55824 25780 55830 25832
rect 13078 25712 13084 25764
rect 13136 25752 13142 25764
rect 14090 25752 14096 25764
rect 13136 25724 14096 25752
rect 13136 25712 13142 25724
rect 14090 25712 14096 25724
rect 14148 25752 14154 25764
rect 14461 25755 14519 25761
rect 14461 25752 14473 25755
rect 14148 25724 14473 25752
rect 14148 25712 14154 25724
rect 14461 25721 14473 25724
rect 14507 25721 14519 25755
rect 14461 25715 14519 25721
rect 19153 25755 19211 25761
rect 19153 25721 19165 25755
rect 19199 25752 19211 25755
rect 20898 25752 20904 25764
rect 19199 25724 20904 25752
rect 19199 25721 19211 25724
rect 19153 25715 19211 25721
rect 20898 25712 20904 25724
rect 20956 25712 20962 25764
rect 21269 25755 21327 25761
rect 21269 25721 21281 25755
rect 21315 25752 21327 25755
rect 21542 25752 21548 25764
rect 21315 25724 21548 25752
rect 21315 25721 21327 25724
rect 21269 25715 21327 25721
rect 21542 25712 21548 25724
rect 21600 25712 21606 25764
rect 24673 25755 24731 25761
rect 24673 25721 24685 25755
rect 24719 25752 24731 25755
rect 34514 25752 34520 25764
rect 24719 25724 34520 25752
rect 24719 25721 24731 25724
rect 24673 25715 24731 25721
rect 34514 25712 34520 25724
rect 34572 25712 34578 25764
rect 37182 25712 37188 25764
rect 37240 25752 37246 25764
rect 38565 25755 38623 25761
rect 38565 25752 38577 25755
rect 37240 25724 38577 25752
rect 37240 25712 37246 25724
rect 38565 25721 38577 25724
rect 38611 25721 38623 25755
rect 38565 25715 38623 25721
rect 11112 25656 11744 25684
rect 11112 25644 11118 25656
rect 18046 25644 18052 25696
rect 18104 25684 18110 25696
rect 23109 25687 23167 25693
rect 23109 25684 23121 25687
rect 18104 25656 23121 25684
rect 18104 25644 18110 25656
rect 23109 25653 23121 25656
rect 23155 25684 23167 25687
rect 23934 25684 23940 25696
rect 23155 25656 23940 25684
rect 23155 25653 23167 25656
rect 23109 25647 23167 25653
rect 23934 25644 23940 25656
rect 23992 25644 23998 25696
rect 30745 25687 30803 25693
rect 30745 25653 30757 25687
rect 30791 25684 30803 25687
rect 40126 25684 40132 25696
rect 30791 25656 40132 25684
rect 30791 25653 30803 25656
rect 30745 25647 30803 25653
rect 40126 25644 40132 25656
rect 40184 25644 40190 25696
rect 53190 25644 53196 25696
rect 53248 25684 53254 25696
rect 53837 25687 53895 25693
rect 53837 25684 53849 25687
rect 53248 25656 53849 25684
rect 53248 25644 53254 25656
rect 53837 25653 53849 25656
rect 53883 25653 53895 25687
rect 53837 25647 53895 25653
rect 1104 25594 58880 25616
rect 1104 25542 4214 25594
rect 4266 25542 4278 25594
rect 4330 25542 4342 25594
rect 4394 25542 4406 25594
rect 4458 25542 4470 25594
rect 4522 25542 34934 25594
rect 34986 25542 34998 25594
rect 35050 25542 35062 25594
rect 35114 25542 35126 25594
rect 35178 25542 35190 25594
rect 35242 25542 58880 25594
rect 1104 25520 58880 25542
rect 6549 25483 6607 25489
rect 6549 25449 6561 25483
rect 6595 25480 6607 25483
rect 6638 25480 6644 25492
rect 6595 25452 6644 25480
rect 6595 25449 6607 25452
rect 6549 25443 6607 25449
rect 6638 25440 6644 25452
rect 6696 25440 6702 25492
rect 9858 25440 9864 25492
rect 9916 25480 9922 25492
rect 10137 25483 10195 25489
rect 10137 25480 10149 25483
rect 9916 25452 10149 25480
rect 9916 25440 9922 25452
rect 10137 25449 10149 25452
rect 10183 25449 10195 25483
rect 10318 25480 10324 25492
rect 10279 25452 10324 25480
rect 10137 25443 10195 25449
rect 10318 25440 10324 25452
rect 10376 25440 10382 25492
rect 18509 25483 18567 25489
rect 18509 25449 18521 25483
rect 18555 25480 18567 25483
rect 20714 25480 20720 25492
rect 18555 25452 20720 25480
rect 18555 25449 18567 25452
rect 18509 25443 18567 25449
rect 20714 25440 20720 25452
rect 20772 25440 20778 25492
rect 21726 25480 21732 25492
rect 21687 25452 21732 25480
rect 21726 25440 21732 25452
rect 21784 25480 21790 25492
rect 22186 25480 22192 25492
rect 21784 25452 22192 25480
rect 21784 25440 21790 25452
rect 22186 25440 22192 25452
rect 22244 25440 22250 25492
rect 43806 25480 43812 25492
rect 28920 25452 41414 25480
rect 43767 25452 43812 25480
rect 3050 25372 3056 25424
rect 3108 25372 3114 25424
rect 3510 25372 3516 25424
rect 3568 25412 3574 25424
rect 4341 25415 4399 25421
rect 4341 25412 4353 25415
rect 3568 25384 4353 25412
rect 3568 25372 3574 25384
rect 4341 25381 4353 25384
rect 4387 25381 4399 25415
rect 4341 25375 4399 25381
rect 14550 25372 14556 25424
rect 14608 25372 14614 25424
rect 17221 25415 17279 25421
rect 17221 25381 17233 25415
rect 17267 25381 17279 25415
rect 17221 25375 17279 25381
rect 3068 25344 3096 25372
rect 2976 25316 3096 25344
rect 2041 25279 2099 25285
rect 2041 25245 2053 25279
rect 2087 25276 2099 25279
rect 2498 25276 2504 25288
rect 2087 25248 2504 25276
rect 2087 25245 2099 25248
rect 2041 25239 2099 25245
rect 2498 25236 2504 25248
rect 2556 25276 2562 25288
rect 2976 25285 3004 25316
rect 3970 25304 3976 25356
rect 4028 25304 4034 25356
rect 4062 25304 4068 25356
rect 4120 25344 4126 25356
rect 7745 25347 7803 25353
rect 4120 25316 5028 25344
rect 4120 25304 4126 25316
rect 2685 25279 2743 25285
rect 2685 25276 2697 25279
rect 2556 25248 2697 25276
rect 2556 25236 2562 25248
rect 2685 25245 2697 25248
rect 2731 25245 2743 25279
rect 2685 25239 2743 25245
rect 2961 25279 3019 25285
rect 2961 25245 2973 25279
rect 3007 25245 3019 25279
rect 2961 25239 3019 25245
rect 3053 25279 3111 25285
rect 3053 25245 3065 25279
rect 3099 25276 3111 25279
rect 3142 25276 3148 25288
rect 3099 25248 3148 25276
rect 3099 25245 3111 25248
rect 3053 25239 3111 25245
rect 3142 25236 3148 25248
rect 3200 25236 3206 25288
rect 3786 25276 3792 25288
rect 3747 25248 3792 25276
rect 3786 25236 3792 25248
rect 3844 25236 3850 25288
rect 3988 25276 4016 25304
rect 4157 25279 4215 25285
rect 3988 25248 4108 25276
rect 1854 25208 1860 25220
rect 1815 25180 1860 25208
rect 1854 25168 1860 25180
rect 1912 25168 1918 25220
rect 2590 25168 2596 25220
rect 2648 25208 2654 25220
rect 4080 25217 4108 25248
rect 4157 25245 4169 25279
rect 4203 25245 4215 25279
rect 4157 25239 4215 25245
rect 2869 25211 2927 25217
rect 2869 25208 2881 25211
rect 2648 25180 2881 25208
rect 2648 25168 2654 25180
rect 2869 25177 2881 25180
rect 2915 25177 2927 25211
rect 2869 25171 2927 25177
rect 3973 25211 4031 25217
rect 3973 25177 3985 25211
rect 4019 25177 4031 25211
rect 3973 25171 4031 25177
rect 4065 25211 4123 25217
rect 4065 25177 4077 25211
rect 4111 25177 4123 25211
rect 4172 25208 4200 25239
rect 4246 25236 4252 25288
rect 4304 25276 4310 25288
rect 5000 25285 5028 25316
rect 7745 25313 7757 25347
rect 7791 25344 7803 25347
rect 9398 25344 9404 25356
rect 7791 25316 9404 25344
rect 7791 25313 7803 25316
rect 7745 25307 7803 25313
rect 9398 25304 9404 25316
rect 9456 25304 9462 25356
rect 13630 25344 13636 25356
rect 13372 25316 13636 25344
rect 4801 25279 4859 25285
rect 4801 25276 4813 25279
rect 4304 25248 4813 25276
rect 4304 25236 4310 25248
rect 4801 25245 4813 25248
rect 4847 25245 4859 25279
rect 4801 25239 4859 25245
rect 4985 25279 5043 25285
rect 4985 25245 4997 25279
rect 5031 25245 5043 25279
rect 8021 25279 8079 25285
rect 8021 25276 8033 25279
rect 4985 25239 5043 25245
rect 6380 25248 8033 25276
rect 4893 25211 4951 25217
rect 4893 25208 4905 25211
rect 4172 25180 4905 25208
rect 4065 25171 4123 25177
rect 4893 25177 4905 25180
rect 4939 25177 4951 25211
rect 4893 25171 4951 25177
rect 3237 25143 3295 25149
rect 3237 25109 3249 25143
rect 3283 25140 3295 25143
rect 3988 25140 4016 25171
rect 6270 25168 6276 25220
rect 6328 25208 6334 25220
rect 6380 25217 6408 25248
rect 8021 25245 8033 25248
rect 8067 25245 8079 25279
rect 8021 25239 8079 25245
rect 12434 25236 12440 25288
rect 12492 25276 12498 25288
rect 12986 25276 12992 25288
rect 12492 25248 12992 25276
rect 12492 25236 12498 25248
rect 12986 25236 12992 25248
rect 13044 25236 13050 25288
rect 13372 25285 13400 25316
rect 13630 25304 13636 25316
rect 13688 25304 13694 25356
rect 13998 25304 14004 25356
rect 14056 25344 14062 25356
rect 14568 25344 14596 25372
rect 14056 25316 14596 25344
rect 14056 25304 14062 25316
rect 14292 25285 14320 25316
rect 13357 25279 13415 25285
rect 13357 25245 13369 25279
rect 13403 25245 13415 25279
rect 14093 25279 14151 25285
rect 14093 25276 14105 25279
rect 13357 25239 13415 25245
rect 13556 25248 14105 25276
rect 6365 25211 6423 25217
rect 6365 25208 6377 25211
rect 6328 25180 6377 25208
rect 6328 25168 6334 25180
rect 6365 25177 6377 25180
rect 6411 25177 6423 25211
rect 6365 25171 6423 25177
rect 6565 25211 6623 25217
rect 6565 25177 6577 25211
rect 6611 25208 6623 25211
rect 6822 25208 6828 25220
rect 6611 25180 6828 25208
rect 6611 25177 6623 25180
rect 6565 25171 6623 25177
rect 6822 25168 6828 25180
rect 6880 25168 6886 25220
rect 9953 25211 10011 25217
rect 9953 25177 9965 25211
rect 9999 25208 10011 25211
rect 10042 25208 10048 25220
rect 9999 25180 10048 25208
rect 9999 25177 10011 25180
rect 9953 25171 10011 25177
rect 10042 25168 10048 25180
rect 10100 25168 10106 25220
rect 10169 25211 10227 25217
rect 10169 25177 10181 25211
rect 10215 25208 10227 25211
rect 10686 25208 10692 25220
rect 10215 25180 10692 25208
rect 10215 25177 10227 25180
rect 10169 25171 10227 25177
rect 10686 25168 10692 25180
rect 10744 25168 10750 25220
rect 13170 25208 13176 25220
rect 13131 25180 13176 25208
rect 13170 25168 13176 25180
rect 13228 25168 13234 25220
rect 13265 25211 13323 25217
rect 13265 25177 13277 25211
rect 13311 25177 13323 25211
rect 13265 25171 13323 25177
rect 3283 25112 4016 25140
rect 6733 25143 6791 25149
rect 3283 25109 3295 25112
rect 3237 25103 3295 25109
rect 6733 25109 6745 25143
rect 6779 25140 6791 25143
rect 7006 25140 7012 25152
rect 6779 25112 7012 25140
rect 6779 25109 6791 25112
rect 6733 25103 6791 25109
rect 7006 25100 7012 25112
rect 7064 25100 7070 25152
rect 12710 25100 12716 25152
rect 12768 25140 12774 25152
rect 13280 25140 13308 25171
rect 13556 25149 13584 25248
rect 14093 25245 14105 25248
rect 14139 25245 14151 25279
rect 14093 25239 14151 25245
rect 14241 25279 14320 25285
rect 14241 25245 14253 25279
rect 14287 25248 14320 25279
rect 14599 25279 14657 25285
rect 14287 25245 14299 25248
rect 14241 25239 14299 25245
rect 14599 25245 14611 25279
rect 14645 25276 14657 25279
rect 14918 25276 14924 25288
rect 14645 25248 14924 25276
rect 14645 25245 14657 25248
rect 14599 25239 14657 25245
rect 14918 25236 14924 25248
rect 14976 25236 14982 25288
rect 16669 25279 16727 25285
rect 16669 25245 16681 25279
rect 16715 25276 16727 25279
rect 16758 25276 16764 25288
rect 16715 25248 16764 25276
rect 16715 25245 16727 25248
rect 16669 25239 16727 25245
rect 16758 25236 16764 25248
rect 16816 25236 16822 25288
rect 17037 25279 17095 25285
rect 17037 25245 17049 25279
rect 17083 25276 17095 25279
rect 17126 25276 17132 25288
rect 17083 25248 17132 25276
rect 17083 25245 17095 25248
rect 17037 25239 17095 25245
rect 17126 25236 17132 25248
rect 17184 25236 17190 25288
rect 17236 25276 17264 25375
rect 20162 25372 20168 25424
rect 20220 25412 20226 25424
rect 20533 25415 20591 25421
rect 20533 25412 20545 25415
rect 20220 25384 20545 25412
rect 20220 25372 20226 25384
rect 20533 25381 20545 25384
rect 20579 25381 20591 25415
rect 20533 25375 20591 25381
rect 21542 25372 21548 25424
rect 21600 25412 21606 25424
rect 24486 25412 24492 25424
rect 21600 25384 24492 25412
rect 21600 25372 21606 25384
rect 24486 25372 24492 25384
rect 24544 25412 24550 25424
rect 24544 25384 24900 25412
rect 24544 25372 24550 25384
rect 17402 25304 17408 25356
rect 17460 25344 17466 25356
rect 23661 25347 23719 25353
rect 17460 25316 22094 25344
rect 17460 25304 17466 25316
rect 17865 25279 17923 25285
rect 17865 25276 17877 25279
rect 17236 25248 17877 25276
rect 17865 25245 17877 25248
rect 17911 25245 17923 25279
rect 17865 25239 17923 25245
rect 17954 25236 17960 25288
rect 18012 25276 18018 25288
rect 18230 25276 18236 25288
rect 18012 25248 18057 25276
rect 18191 25248 18236 25276
rect 18012 25236 18018 25248
rect 18230 25236 18236 25248
rect 18288 25236 18294 25288
rect 18322 25236 18328 25288
rect 18380 25285 18386 25288
rect 18380 25276 18388 25285
rect 18380 25248 18425 25276
rect 18380 25239 18388 25248
rect 18380 25236 18386 25239
rect 20622 25236 20628 25288
rect 20680 25276 20686 25288
rect 21637 25279 21695 25285
rect 21637 25276 21649 25279
rect 20680 25248 21649 25276
rect 20680 25236 20686 25248
rect 21637 25245 21649 25248
rect 21683 25245 21695 25279
rect 22066 25276 22094 25316
rect 23661 25313 23673 25347
rect 23707 25344 23719 25347
rect 23707 25316 24440 25344
rect 23707 25313 23719 25316
rect 23661 25307 23719 25313
rect 22925 25279 22983 25285
rect 22925 25276 22937 25279
rect 22066 25248 22937 25276
rect 21637 25239 21695 25245
rect 22925 25245 22937 25248
rect 22971 25276 22983 25279
rect 23382 25276 23388 25288
rect 22971 25248 23388 25276
rect 22971 25245 22983 25248
rect 22925 25239 22983 25245
rect 23382 25236 23388 25248
rect 23440 25236 23446 25288
rect 23566 25276 23572 25288
rect 23527 25248 23572 25276
rect 23566 25236 23572 25248
rect 23624 25236 23630 25288
rect 23750 25276 23756 25288
rect 23711 25248 23756 25276
rect 23750 25236 23756 25248
rect 23808 25236 23814 25288
rect 24412 25285 24440 25316
rect 24578 25285 24584 25288
rect 24397 25279 24455 25285
rect 24397 25245 24409 25279
rect 24443 25245 24455 25279
rect 24397 25239 24455 25245
rect 24545 25279 24584 25285
rect 24545 25245 24557 25279
rect 24545 25239 24584 25245
rect 24578 25236 24584 25239
rect 24636 25236 24642 25288
rect 24872 25285 24900 25384
rect 27706 25304 27712 25356
rect 27764 25344 27770 25356
rect 28258 25344 28264 25356
rect 27764 25316 28264 25344
rect 27764 25304 27770 25316
rect 28258 25304 28264 25316
rect 28316 25344 28322 25356
rect 28920 25353 28948 25452
rect 30650 25412 30656 25424
rect 30611 25384 30656 25412
rect 30650 25372 30656 25384
rect 30708 25412 30714 25424
rect 31757 25415 31815 25421
rect 30708 25384 31432 25412
rect 30708 25372 30714 25384
rect 28905 25347 28963 25353
rect 28316 25316 28396 25344
rect 28316 25304 28322 25316
rect 24862 25279 24920 25285
rect 24862 25245 24874 25279
rect 24908 25245 24920 25279
rect 27614 25276 27620 25288
rect 27575 25248 27620 25276
rect 24862 25239 24920 25245
rect 27614 25236 27620 25248
rect 27672 25236 27678 25288
rect 27801 25279 27859 25285
rect 27801 25245 27813 25279
rect 27847 25276 27859 25279
rect 28166 25276 28172 25288
rect 27847 25248 28172 25276
rect 27847 25245 27859 25248
rect 27801 25239 27859 25245
rect 28166 25236 28172 25248
rect 28224 25236 28230 25288
rect 28368 25285 28396 25316
rect 28905 25313 28917 25347
rect 28951 25313 28963 25347
rect 31294 25344 31300 25356
rect 31255 25316 31300 25344
rect 28905 25307 28963 25313
rect 31294 25304 31300 25316
rect 31352 25304 31358 25356
rect 31404 25288 31432 25384
rect 31757 25381 31769 25415
rect 31803 25412 31815 25415
rect 33686 25412 33692 25424
rect 31803 25384 33692 25412
rect 31803 25381 31815 25384
rect 31757 25375 31815 25381
rect 33686 25372 33692 25384
rect 33744 25372 33750 25424
rect 34606 25412 34612 25424
rect 33796 25384 34612 25412
rect 28353 25279 28411 25285
rect 28353 25245 28365 25279
rect 28399 25245 28411 25279
rect 28718 25276 28724 25288
rect 28679 25248 28724 25276
rect 28353 25239 28411 25245
rect 28718 25236 28724 25248
rect 28776 25236 28782 25288
rect 31386 25276 31392 25288
rect 31299 25248 31392 25276
rect 31386 25236 31392 25248
rect 31444 25236 31450 25288
rect 14369 25211 14427 25217
rect 14369 25177 14381 25211
rect 14415 25177 14427 25211
rect 14369 25171 14427 25177
rect 12768 25112 13308 25140
rect 13541 25143 13599 25149
rect 12768 25100 12774 25112
rect 13541 25109 13553 25143
rect 13587 25109 13599 25143
rect 13541 25103 13599 25109
rect 14090 25100 14096 25152
rect 14148 25140 14154 25152
rect 14384 25140 14412 25171
rect 14458 25168 14464 25220
rect 14516 25208 14522 25220
rect 16850 25208 16856 25220
rect 14516 25180 14561 25208
rect 16811 25180 16856 25208
rect 14516 25168 14522 25180
rect 16850 25168 16856 25180
rect 16908 25168 16914 25220
rect 16945 25211 17003 25217
rect 16945 25177 16957 25211
rect 16991 25208 17003 25211
rect 17310 25208 17316 25220
rect 16991 25180 17316 25208
rect 16991 25177 17003 25180
rect 16945 25171 17003 25177
rect 17310 25168 17316 25180
rect 17368 25168 17374 25220
rect 18138 25208 18144 25220
rect 18099 25180 18144 25208
rect 18138 25168 18144 25180
rect 18196 25168 18202 25220
rect 18248 25208 18276 25236
rect 18690 25208 18696 25220
rect 18248 25180 18696 25208
rect 18690 25168 18696 25180
rect 18748 25168 18754 25220
rect 21726 25168 21732 25220
rect 21784 25208 21790 25220
rect 22741 25211 22799 25217
rect 22741 25208 22753 25211
rect 21784 25180 22753 25208
rect 21784 25168 21790 25180
rect 22741 25177 22753 25180
rect 22787 25208 22799 25211
rect 24673 25211 24731 25217
rect 24673 25208 24685 25211
rect 22787 25180 24685 25208
rect 22787 25177 22799 25180
rect 22741 25171 22799 25177
rect 24673 25177 24685 25180
rect 24719 25177 24731 25211
rect 24673 25171 24731 25177
rect 24762 25168 24768 25220
rect 24820 25208 24826 25220
rect 33796 25208 33824 25384
rect 34606 25372 34612 25384
rect 34664 25372 34670 25424
rect 35253 25415 35311 25421
rect 35253 25381 35265 25415
rect 35299 25412 35311 25415
rect 37458 25412 37464 25424
rect 35299 25384 37464 25412
rect 35299 25381 35311 25384
rect 35253 25375 35311 25381
rect 37458 25372 37464 25384
rect 37516 25372 37522 25424
rect 38010 25412 38016 25424
rect 37971 25384 38016 25412
rect 38010 25372 38016 25384
rect 38068 25372 38074 25424
rect 38102 25372 38108 25424
rect 38160 25412 38166 25424
rect 41386 25412 41414 25452
rect 43806 25440 43812 25452
rect 43864 25440 43870 25492
rect 46477 25483 46535 25489
rect 46477 25449 46489 25483
rect 46523 25480 46535 25483
rect 47578 25480 47584 25492
rect 46523 25452 47584 25480
rect 46523 25449 46535 25452
rect 46477 25443 46535 25449
rect 47578 25440 47584 25452
rect 47636 25440 47642 25492
rect 50154 25480 50160 25492
rect 50115 25452 50160 25480
rect 50154 25440 50160 25452
rect 50212 25440 50218 25492
rect 52822 25480 52828 25492
rect 52783 25452 52828 25480
rect 52822 25440 52828 25452
rect 52880 25440 52886 25492
rect 54665 25483 54723 25489
rect 54665 25449 54677 25483
rect 54711 25480 54723 25483
rect 55950 25480 55956 25492
rect 54711 25452 55812 25480
rect 55911 25452 55956 25480
rect 54711 25449 54723 25452
rect 54665 25443 54723 25449
rect 52546 25412 52552 25424
rect 38160 25384 38205 25412
rect 41386 25384 52552 25412
rect 38160 25372 38166 25384
rect 52546 25372 52552 25384
rect 52604 25372 52610 25424
rect 34793 25347 34851 25353
rect 34793 25344 34805 25347
rect 24820 25180 24865 25208
rect 25056 25180 33824 25208
rect 34072 25316 34805 25344
rect 24820 25168 24826 25180
rect 14734 25140 14740 25152
rect 14148 25112 14412 25140
rect 14695 25112 14740 25140
rect 14148 25100 14154 25112
rect 14734 25100 14740 25112
rect 14792 25100 14798 25152
rect 18230 25100 18236 25152
rect 18288 25140 18294 25152
rect 18506 25140 18512 25152
rect 18288 25112 18512 25140
rect 18288 25100 18294 25112
rect 18506 25100 18512 25112
rect 18564 25140 18570 25152
rect 21358 25140 21364 25152
rect 18564 25112 21364 25140
rect 18564 25100 18570 25112
rect 21358 25100 21364 25112
rect 21416 25100 21422 25152
rect 25056 25149 25084 25180
rect 34072 25152 34100 25316
rect 34793 25313 34805 25316
rect 34839 25313 34851 25347
rect 34793 25307 34851 25313
rect 40497 25347 40555 25353
rect 40497 25313 40509 25347
rect 40543 25344 40555 25347
rect 40543 25316 41184 25344
rect 40543 25313 40555 25316
rect 40497 25307 40555 25313
rect 34698 25236 34704 25288
rect 34756 25276 34762 25288
rect 34885 25279 34943 25285
rect 34885 25276 34897 25279
rect 34756 25248 34897 25276
rect 34756 25236 34762 25248
rect 34885 25245 34897 25248
rect 34931 25276 34943 25279
rect 35713 25279 35771 25285
rect 35713 25276 35725 25279
rect 34931 25248 35725 25276
rect 34931 25245 34943 25248
rect 34885 25239 34943 25245
rect 35713 25245 35725 25248
rect 35759 25245 35771 25279
rect 40126 25276 40132 25288
rect 40087 25248 40132 25276
rect 35713 25239 35771 25245
rect 40126 25236 40132 25248
rect 40184 25236 40190 25288
rect 40954 25276 40960 25288
rect 40915 25248 40960 25276
rect 40954 25236 40960 25248
rect 41012 25236 41018 25288
rect 41156 25285 41184 25316
rect 49234 25304 49240 25356
rect 49292 25344 49298 25356
rect 50249 25347 50307 25353
rect 50249 25344 50261 25347
rect 49292 25316 50261 25344
rect 49292 25304 49298 25316
rect 50249 25313 50261 25316
rect 50295 25313 50307 25347
rect 50249 25307 50307 25313
rect 52362 25304 52368 25356
rect 52420 25344 52426 25356
rect 52825 25347 52883 25353
rect 52825 25344 52837 25347
rect 52420 25316 52837 25344
rect 52420 25304 52426 25316
rect 52825 25313 52837 25316
rect 52871 25313 52883 25347
rect 52825 25307 52883 25313
rect 52914 25304 52920 25356
rect 52972 25344 52978 25356
rect 53101 25347 53159 25353
rect 52972 25316 53017 25344
rect 52972 25304 52978 25316
rect 53101 25313 53113 25347
rect 53147 25344 53159 25347
rect 53147 25316 53696 25344
rect 53147 25313 53159 25316
rect 53101 25307 53159 25313
rect 53668 25288 53696 25316
rect 55582 25304 55588 25356
rect 55640 25344 55646 25356
rect 55784 25353 55812 25452
rect 55950 25440 55956 25452
rect 56008 25440 56014 25492
rect 55769 25347 55827 25353
rect 55640 25316 55685 25344
rect 55640 25304 55646 25316
rect 55769 25313 55781 25347
rect 55815 25344 55827 25347
rect 55858 25344 55864 25356
rect 55815 25316 55864 25344
rect 55815 25313 55827 25316
rect 55769 25307 55827 25313
rect 55858 25304 55864 25316
rect 55916 25304 55922 25356
rect 41141 25279 41199 25285
rect 41141 25245 41153 25279
rect 41187 25245 41199 25279
rect 41141 25239 41199 25245
rect 41325 25279 41383 25285
rect 41325 25245 41337 25279
rect 41371 25276 41383 25279
rect 41874 25276 41880 25288
rect 41371 25248 41880 25276
rect 41371 25245 41383 25248
rect 41325 25239 41383 25245
rect 41874 25236 41880 25248
rect 41932 25276 41938 25288
rect 41969 25279 42027 25285
rect 41969 25276 41981 25279
rect 41932 25248 41981 25276
rect 41932 25236 41938 25248
rect 41969 25245 41981 25248
rect 42015 25245 42027 25279
rect 41969 25239 42027 25245
rect 42153 25279 42211 25285
rect 42153 25245 42165 25279
rect 42199 25276 42211 25279
rect 42613 25279 42671 25285
rect 42613 25276 42625 25279
rect 42199 25248 42625 25276
rect 42199 25245 42211 25248
rect 42153 25239 42211 25245
rect 42613 25245 42625 25248
rect 42659 25245 42671 25279
rect 42794 25276 42800 25288
rect 42755 25248 42800 25276
rect 42613 25239 42671 25245
rect 42794 25236 42800 25248
rect 42852 25236 42858 25288
rect 42981 25279 43039 25285
rect 42981 25245 42993 25279
rect 43027 25276 43039 25279
rect 43714 25276 43720 25288
rect 43027 25248 43720 25276
rect 43027 25245 43039 25248
rect 42981 25239 43039 25245
rect 43714 25236 43720 25248
rect 43772 25236 43778 25288
rect 45738 25236 45744 25288
rect 45796 25276 45802 25288
rect 45833 25279 45891 25285
rect 45833 25276 45845 25279
rect 45796 25248 45845 25276
rect 45796 25236 45802 25248
rect 45833 25245 45845 25248
rect 45879 25245 45891 25279
rect 45833 25239 45891 25245
rect 45922 25236 45928 25288
rect 45980 25276 45986 25288
rect 46017 25279 46075 25285
rect 46017 25276 46029 25279
rect 45980 25248 46029 25276
rect 45980 25236 45986 25248
rect 46017 25245 46029 25248
rect 46063 25245 46075 25279
rect 46017 25239 46075 25245
rect 46106 25236 46112 25288
rect 46164 25276 46170 25288
rect 46290 25285 46296 25288
rect 46247 25279 46296 25285
rect 46164 25248 46209 25276
rect 46164 25236 46170 25248
rect 46247 25245 46259 25279
rect 46293 25245 46296 25279
rect 46247 25239 46296 25245
rect 46290 25236 46296 25239
rect 46348 25276 46354 25288
rect 46842 25276 46848 25288
rect 46348 25248 46848 25276
rect 46348 25236 46354 25248
rect 46842 25236 46848 25248
rect 46900 25236 46906 25288
rect 50154 25276 50160 25288
rect 50115 25248 50160 25276
rect 50154 25236 50160 25248
rect 50212 25236 50218 25288
rect 53190 25276 53196 25288
rect 53151 25248 53196 25276
rect 53190 25236 53196 25248
rect 53248 25236 53254 25288
rect 53650 25236 53656 25288
rect 53708 25276 53714 25288
rect 54573 25279 54631 25285
rect 54573 25276 54585 25279
rect 53708 25248 54585 25276
rect 53708 25236 53714 25248
rect 54573 25245 54585 25248
rect 54619 25245 54631 25279
rect 54573 25239 54631 25245
rect 55398 25236 55404 25288
rect 55456 25276 55462 25288
rect 55493 25279 55551 25285
rect 55493 25276 55505 25279
rect 55456 25248 55505 25276
rect 55456 25236 55462 25248
rect 55493 25245 55505 25248
rect 55539 25245 55551 25279
rect 55493 25239 55551 25245
rect 55677 25279 55735 25285
rect 55677 25245 55689 25279
rect 55723 25276 55735 25279
rect 57882 25276 57888 25288
rect 55723 25248 55812 25276
rect 57843 25248 57888 25276
rect 55723 25245 55735 25248
rect 55677 25239 55735 25245
rect 37182 25168 37188 25220
rect 37240 25208 37246 25220
rect 37645 25211 37703 25217
rect 37645 25208 37657 25211
rect 37240 25180 37657 25208
rect 37240 25168 37246 25180
rect 37645 25177 37657 25180
rect 37691 25177 37703 25211
rect 40310 25208 40316 25220
rect 40271 25180 40316 25208
rect 37645 25171 37703 25177
rect 40310 25168 40316 25180
rect 40368 25168 40374 25220
rect 41598 25168 41604 25220
rect 41656 25208 41662 25220
rect 41785 25211 41843 25217
rect 41785 25208 41797 25211
rect 41656 25180 41797 25208
rect 41656 25168 41662 25180
rect 41785 25177 41797 25180
rect 41831 25177 41843 25211
rect 55784 25208 55812 25248
rect 57882 25236 57888 25248
rect 57940 25236 57946 25288
rect 41785 25171 41843 25177
rect 55692 25180 55812 25208
rect 55692 25152 55720 25180
rect 25041 25143 25099 25149
rect 25041 25109 25053 25143
rect 25087 25109 25099 25143
rect 25041 25103 25099 25109
rect 26602 25100 26608 25152
rect 26660 25140 26666 25152
rect 27525 25143 27583 25149
rect 27525 25140 27537 25143
rect 26660 25112 27537 25140
rect 26660 25100 26666 25112
rect 27525 25109 27537 25112
rect 27571 25109 27583 25143
rect 34054 25140 34060 25152
rect 34015 25112 34060 25140
rect 27525 25103 27583 25109
rect 34054 25100 34060 25112
rect 34112 25100 34118 25152
rect 44174 25140 44180 25152
rect 44135 25112 44180 25140
rect 44174 25100 44180 25112
rect 44232 25100 44238 25152
rect 50525 25143 50583 25149
rect 50525 25109 50537 25143
rect 50571 25140 50583 25143
rect 52270 25140 52276 25152
rect 50571 25112 52276 25140
rect 50571 25109 50583 25112
rect 50525 25103 50583 25109
rect 52270 25100 52276 25112
rect 52328 25100 52334 25152
rect 55674 25100 55680 25152
rect 55732 25100 55738 25152
rect 58066 25140 58072 25152
rect 58027 25112 58072 25140
rect 58066 25100 58072 25112
rect 58124 25100 58130 25152
rect 1104 25050 58880 25072
rect 1104 24998 19574 25050
rect 19626 24998 19638 25050
rect 19690 24998 19702 25050
rect 19754 24998 19766 25050
rect 19818 24998 19830 25050
rect 19882 24998 50294 25050
rect 50346 24998 50358 25050
rect 50410 24998 50422 25050
rect 50474 24998 50486 25050
rect 50538 24998 50550 25050
rect 50602 24998 58880 25050
rect 1104 24976 58880 24998
rect 1673 24939 1731 24945
rect 1673 24905 1685 24939
rect 1719 24936 1731 24939
rect 1854 24936 1860 24948
rect 1719 24908 1860 24936
rect 1719 24905 1731 24908
rect 1673 24899 1731 24905
rect 1854 24896 1860 24908
rect 1912 24896 1918 24948
rect 3050 24896 3056 24948
rect 3108 24936 3114 24948
rect 3237 24939 3295 24945
rect 3237 24936 3249 24939
rect 3108 24908 3249 24936
rect 3108 24896 3114 24908
rect 3237 24905 3249 24908
rect 3283 24936 3295 24939
rect 3878 24936 3884 24948
rect 3283 24908 3884 24936
rect 3283 24905 3295 24908
rect 3237 24899 3295 24905
rect 3878 24896 3884 24908
rect 3936 24936 3942 24948
rect 4065 24939 4123 24945
rect 4065 24936 4077 24939
rect 3936 24908 4077 24936
rect 3936 24896 3942 24908
rect 4065 24905 4077 24908
rect 4111 24905 4123 24939
rect 4065 24899 4123 24905
rect 8294 24896 8300 24948
rect 8352 24896 8358 24948
rect 8478 24896 8484 24948
rect 8536 24936 8542 24948
rect 15654 24936 15660 24948
rect 8536 24908 15660 24936
rect 8536 24896 8542 24908
rect 15654 24896 15660 24908
rect 15712 24896 15718 24948
rect 17954 24896 17960 24948
rect 18012 24936 18018 24948
rect 18012 24908 22416 24936
rect 18012 24896 18018 24908
rect 8202 24868 8208 24880
rect 8163 24840 8208 24868
rect 8202 24828 8208 24840
rect 8260 24828 8266 24880
rect 8312 24831 8340 24896
rect 8306 24825 8364 24831
rect 11974 24828 11980 24880
rect 12032 24868 12038 24880
rect 16482 24868 16488 24880
rect 12032 24840 16488 24868
rect 12032 24828 12038 24840
rect 16482 24828 16488 24840
rect 16540 24828 16546 24880
rect 17218 24828 17224 24880
rect 17276 24868 17282 24880
rect 17865 24871 17923 24877
rect 17865 24868 17877 24871
rect 17276 24840 17877 24868
rect 17276 24828 17282 24840
rect 17865 24837 17877 24840
rect 17911 24837 17923 24871
rect 17865 24831 17923 24837
rect 20162 24828 20168 24880
rect 20220 24868 20226 24880
rect 21266 24868 21272 24880
rect 20220 24840 21272 24868
rect 20220 24828 20226 24840
rect 2498 24800 2504 24812
rect 2459 24772 2504 24800
rect 2498 24760 2504 24772
rect 2556 24760 2562 24812
rect 2590 24760 2596 24812
rect 2648 24800 2654 24812
rect 2685 24803 2743 24809
rect 2685 24800 2697 24803
rect 2648 24772 2697 24800
rect 2648 24760 2654 24772
rect 2685 24769 2697 24772
rect 2731 24769 2743 24803
rect 3142 24800 3148 24812
rect 3103 24772 3148 24800
rect 2685 24763 2743 24769
rect 3142 24760 3148 24772
rect 3200 24760 3206 24812
rect 3418 24800 3424 24812
rect 3379 24772 3424 24800
rect 3418 24760 3424 24772
rect 3476 24760 3482 24812
rect 6917 24803 6975 24809
rect 6917 24769 6929 24803
rect 6963 24769 6975 24803
rect 6917 24763 6975 24769
rect 2317 24735 2375 24741
rect 2317 24701 2329 24735
rect 2363 24732 2375 24735
rect 3786 24732 3792 24744
rect 2363 24704 3792 24732
rect 2363 24701 2375 24704
rect 2317 24695 2375 24701
rect 3786 24692 3792 24704
rect 3844 24692 3850 24744
rect 6932 24732 6960 24763
rect 7006 24760 7012 24812
rect 7064 24800 7070 24812
rect 7190 24800 7196 24812
rect 7064 24772 7109 24800
rect 7151 24772 7196 24800
rect 7064 24760 7070 24772
rect 7190 24760 7196 24772
rect 7248 24760 7254 24812
rect 7282 24760 7288 24812
rect 7340 24800 7346 24812
rect 7466 24800 7472 24812
rect 7340 24772 7385 24800
rect 7427 24772 7472 24800
rect 7340 24760 7346 24772
rect 7466 24760 7472 24772
rect 7524 24760 7530 24812
rect 8018 24800 8024 24812
rect 7979 24772 8024 24800
rect 8018 24760 8024 24772
rect 8076 24760 8082 24812
rect 8306 24791 8318 24825
rect 8352 24791 8364 24825
rect 8306 24785 8364 24791
rect 8662 24760 8668 24812
rect 8720 24800 8726 24812
rect 9674 24800 9680 24812
rect 8720 24772 9680 24800
rect 8720 24760 8726 24772
rect 9674 24760 9680 24772
rect 9732 24760 9738 24812
rect 10042 24760 10048 24812
rect 10100 24800 10106 24812
rect 10229 24803 10287 24809
rect 10229 24800 10241 24803
rect 10100 24772 10241 24800
rect 10100 24760 10106 24772
rect 10229 24769 10241 24772
rect 10275 24769 10287 24803
rect 10229 24763 10287 24769
rect 13449 24803 13507 24809
rect 13449 24769 13461 24803
rect 13495 24800 13507 24803
rect 13538 24800 13544 24812
rect 13495 24772 13544 24800
rect 13495 24769 13507 24772
rect 13449 24763 13507 24769
rect 13538 24760 13544 24772
rect 13596 24760 13602 24812
rect 15194 24800 15200 24812
rect 14936 24772 15200 24800
rect 6932 24704 8064 24732
rect 8036 24673 8064 24704
rect 8386 24692 8392 24744
rect 8444 24732 8450 24744
rect 10060 24732 10088 24760
rect 8444 24704 10088 24732
rect 13265 24735 13323 24741
rect 8444 24692 8450 24704
rect 13265 24701 13277 24735
rect 13311 24732 13323 24735
rect 13354 24732 13360 24744
rect 13311 24704 13360 24732
rect 13311 24701 13323 24704
rect 13265 24695 13323 24701
rect 13354 24692 13360 24704
rect 13412 24732 13418 24744
rect 14936 24732 14964 24772
rect 15194 24760 15200 24772
rect 15252 24760 15258 24812
rect 17034 24760 17040 24812
rect 17092 24800 17098 24812
rect 17129 24803 17187 24809
rect 17129 24800 17141 24803
rect 17092 24772 17141 24800
rect 17092 24760 17098 24772
rect 17129 24769 17141 24772
rect 17175 24769 17187 24803
rect 20070 24800 20076 24812
rect 20031 24772 20076 24800
rect 17129 24763 17187 24769
rect 20070 24760 20076 24772
rect 20128 24760 20134 24812
rect 20732 24809 20760 24840
rect 21266 24828 21272 24840
rect 21324 24828 21330 24880
rect 21358 24828 21364 24880
rect 21416 24868 21422 24880
rect 22388 24868 22416 24908
rect 27614 24896 27620 24948
rect 27672 24936 27678 24948
rect 27985 24939 28043 24945
rect 27985 24936 27997 24939
rect 27672 24908 27997 24936
rect 27672 24896 27678 24908
rect 27985 24905 27997 24908
rect 28031 24905 28043 24939
rect 27985 24899 28043 24905
rect 31386 24896 31392 24948
rect 31444 24936 31450 24948
rect 34514 24936 34520 24948
rect 31444 24908 34520 24936
rect 31444 24896 31450 24908
rect 34514 24896 34520 24908
rect 34572 24896 34578 24948
rect 34698 24896 34704 24948
rect 34756 24936 34762 24948
rect 34977 24939 35035 24945
rect 34977 24936 34989 24939
rect 34756 24908 34989 24936
rect 34756 24896 34762 24908
rect 34977 24905 34989 24908
rect 35023 24905 35035 24939
rect 34977 24899 35035 24905
rect 40221 24939 40279 24945
rect 40221 24905 40233 24939
rect 40267 24936 40279 24939
rect 40954 24936 40960 24948
rect 40267 24908 40960 24936
rect 40267 24905 40279 24908
rect 40221 24899 40279 24905
rect 40954 24896 40960 24908
rect 41012 24896 41018 24948
rect 50065 24939 50123 24945
rect 50065 24905 50077 24939
rect 50111 24936 50123 24939
rect 50154 24936 50160 24948
rect 50111 24908 50160 24936
rect 50111 24905 50123 24908
rect 50065 24899 50123 24905
rect 50154 24896 50160 24908
rect 50212 24896 50218 24948
rect 53926 24896 53932 24948
rect 53984 24936 53990 24948
rect 57974 24936 57980 24948
rect 53984 24908 55812 24936
rect 57935 24908 57980 24936
rect 53984 24896 53990 24908
rect 34054 24868 34060 24880
rect 21416 24840 22324 24868
rect 22388 24840 34060 24868
rect 21416 24828 21422 24840
rect 20717 24803 20775 24809
rect 20717 24769 20729 24803
rect 20763 24769 20775 24803
rect 20717 24763 20775 24769
rect 20901 24803 20959 24809
rect 20901 24769 20913 24803
rect 20947 24769 20959 24803
rect 22296 24800 22324 24840
rect 34054 24828 34060 24840
rect 34112 24828 34118 24880
rect 45005 24871 45063 24877
rect 45005 24837 45017 24871
rect 45051 24868 45063 24871
rect 46201 24871 46259 24877
rect 45051 24840 46060 24868
rect 45051 24837 45063 24840
rect 45005 24831 45063 24837
rect 23474 24800 23480 24812
rect 22296 24772 23480 24800
rect 20901 24763 20959 24769
rect 13412 24704 14964 24732
rect 13412 24692 13418 24704
rect 17402 24692 17408 24744
rect 17460 24732 17466 24744
rect 18322 24732 18328 24744
rect 17460 24704 18328 24732
rect 17460 24692 17466 24704
rect 18322 24692 18328 24704
rect 18380 24692 18386 24744
rect 19334 24692 19340 24744
rect 19392 24732 19398 24744
rect 20806 24732 20812 24744
rect 19392 24704 20812 24732
rect 19392 24692 19398 24704
rect 20806 24692 20812 24704
rect 20864 24732 20870 24744
rect 20916 24732 20944 24763
rect 23474 24760 23480 24772
rect 23532 24800 23538 24812
rect 23750 24800 23756 24812
rect 23532 24772 23756 24800
rect 23532 24760 23538 24772
rect 23750 24760 23756 24772
rect 23808 24760 23814 24812
rect 24394 24800 24400 24812
rect 24355 24772 24400 24800
rect 24394 24760 24400 24772
rect 24452 24760 24458 24812
rect 25130 24760 25136 24812
rect 25188 24800 25194 24812
rect 25685 24803 25743 24809
rect 25685 24800 25697 24803
rect 25188 24772 25697 24800
rect 25188 24760 25194 24772
rect 25685 24769 25697 24772
rect 25731 24769 25743 24803
rect 25685 24763 25743 24769
rect 26145 24803 26203 24809
rect 26145 24769 26157 24803
rect 26191 24800 26203 24803
rect 26234 24800 26240 24812
rect 26191 24772 26240 24800
rect 26191 24769 26203 24772
rect 26145 24763 26203 24769
rect 26234 24760 26240 24772
rect 26292 24760 26298 24812
rect 27706 24760 27712 24812
rect 27764 24800 27770 24812
rect 27893 24803 27951 24809
rect 27893 24800 27905 24803
rect 27764 24772 27905 24800
rect 27764 24760 27770 24772
rect 27893 24769 27905 24772
rect 27939 24769 27951 24803
rect 28074 24800 28080 24812
rect 28035 24772 28080 24800
rect 27893 24763 27951 24769
rect 28074 24760 28080 24772
rect 28132 24760 28138 24812
rect 30561 24803 30619 24809
rect 30561 24769 30573 24803
rect 30607 24800 30619 24803
rect 33778 24800 33784 24812
rect 30607 24772 33784 24800
rect 30607 24769 30619 24772
rect 30561 24763 30619 24769
rect 25314 24732 25320 24744
rect 20864 24704 20944 24732
rect 25275 24704 25320 24732
rect 20864 24692 20870 24704
rect 25314 24692 25320 24704
rect 25372 24692 25378 24744
rect 25406 24692 25412 24744
rect 25464 24732 25470 24744
rect 30285 24735 30343 24741
rect 30285 24732 30297 24735
rect 25464 24704 30297 24732
rect 25464 24692 25470 24704
rect 30285 24701 30297 24704
rect 30331 24701 30343 24735
rect 30285 24695 30343 24701
rect 8021 24667 8079 24673
rect 8021 24633 8033 24667
rect 8067 24633 8079 24667
rect 8021 24627 8079 24633
rect 9493 24667 9551 24673
rect 9493 24633 9505 24667
rect 9539 24664 9551 24667
rect 10778 24664 10784 24676
rect 9539 24636 10784 24664
rect 9539 24633 9551 24636
rect 9493 24627 9551 24633
rect 10778 24624 10784 24636
rect 10836 24624 10842 24676
rect 13633 24667 13691 24673
rect 13633 24633 13645 24667
rect 13679 24664 13691 24667
rect 14182 24664 14188 24676
rect 13679 24636 14188 24664
rect 13679 24633 13691 24636
rect 13633 24627 13691 24633
rect 14182 24624 14188 24636
rect 14240 24624 14246 24676
rect 16758 24624 16764 24676
rect 16816 24664 16822 24676
rect 17126 24664 17132 24676
rect 16816 24636 17132 24664
rect 16816 24624 16822 24636
rect 17126 24624 17132 24636
rect 17184 24664 17190 24676
rect 17313 24667 17371 24673
rect 17313 24664 17325 24667
rect 17184 24636 17325 24664
rect 17184 24624 17190 24636
rect 17313 24633 17325 24636
rect 17359 24664 17371 24667
rect 17678 24664 17684 24676
rect 17359 24636 17684 24664
rect 17359 24633 17371 24636
rect 17313 24627 17371 24633
rect 17678 24624 17684 24636
rect 17736 24624 17742 24676
rect 18049 24667 18107 24673
rect 18049 24633 18061 24667
rect 18095 24664 18107 24667
rect 18506 24664 18512 24676
rect 18095 24636 18512 24664
rect 18095 24633 18107 24636
rect 18049 24627 18107 24633
rect 18506 24624 18512 24636
rect 18564 24624 18570 24676
rect 20254 24664 20260 24676
rect 20215 24636 20260 24664
rect 20254 24624 20260 24636
rect 20312 24624 20318 24676
rect 23658 24624 23664 24676
rect 23716 24664 23722 24676
rect 24213 24667 24271 24673
rect 24213 24664 24225 24667
rect 23716 24636 24225 24664
rect 23716 24624 23722 24636
rect 24213 24633 24225 24636
rect 24259 24633 24271 24667
rect 24213 24627 24271 24633
rect 26234 24624 26240 24676
rect 26292 24664 26298 24676
rect 26786 24664 26792 24676
rect 26292 24636 26792 24664
rect 26292 24624 26298 24636
rect 26786 24624 26792 24636
rect 26844 24664 26850 24676
rect 30576 24664 30604 24763
rect 33778 24760 33784 24772
rect 33836 24760 33842 24812
rect 33962 24800 33968 24812
rect 33875 24772 33968 24800
rect 33962 24760 33968 24772
rect 34020 24800 34026 24812
rect 34885 24803 34943 24809
rect 34885 24800 34897 24803
rect 34020 24772 34897 24800
rect 34020 24760 34026 24772
rect 34885 24769 34897 24772
rect 34931 24769 34943 24803
rect 34885 24763 34943 24769
rect 36538 24760 36544 24812
rect 36596 24800 36602 24812
rect 37737 24803 37795 24809
rect 37737 24800 37749 24803
rect 36596 24772 37749 24800
rect 36596 24760 36602 24772
rect 37737 24769 37749 24772
rect 37783 24800 37795 24803
rect 39114 24800 39120 24812
rect 37783 24772 39120 24800
rect 37783 24769 37795 24772
rect 37737 24763 37795 24769
rect 39114 24760 39120 24772
rect 39172 24760 39178 24812
rect 40037 24803 40095 24809
rect 40037 24769 40049 24803
rect 40083 24800 40095 24803
rect 40126 24800 40132 24812
rect 40083 24772 40132 24800
rect 40083 24769 40095 24772
rect 40037 24763 40095 24769
rect 40126 24760 40132 24772
rect 40184 24760 40190 24812
rect 40221 24803 40279 24809
rect 40221 24769 40233 24803
rect 40267 24800 40279 24803
rect 40310 24800 40316 24812
rect 40267 24772 40316 24800
rect 40267 24769 40279 24772
rect 40221 24763 40279 24769
rect 31110 24732 31116 24744
rect 31071 24704 31116 24732
rect 31110 24692 31116 24704
rect 31168 24692 31174 24744
rect 33873 24735 33931 24741
rect 33873 24732 33885 24735
rect 33244 24704 33885 24732
rect 26844 24636 30604 24664
rect 26844 24624 26850 24636
rect 33244 24608 33272 24704
rect 33873 24701 33885 24704
rect 33919 24701 33931 24735
rect 33873 24695 33931 24701
rect 37829 24735 37887 24741
rect 37829 24701 37841 24735
rect 37875 24732 37887 24735
rect 38562 24732 38568 24744
rect 37875 24704 38568 24732
rect 37875 24701 37887 24704
rect 37829 24695 37887 24701
rect 38562 24692 38568 24704
rect 38620 24692 38626 24744
rect 34333 24667 34391 24673
rect 34333 24633 34345 24667
rect 34379 24664 34391 24667
rect 40236 24664 40264 24763
rect 40310 24760 40316 24772
rect 40368 24760 40374 24812
rect 41598 24800 41604 24812
rect 41559 24772 41604 24800
rect 41598 24760 41604 24772
rect 41656 24760 41662 24812
rect 41785 24803 41843 24809
rect 41785 24769 41797 24803
rect 41831 24800 41843 24803
rect 41874 24800 41880 24812
rect 41831 24772 41880 24800
rect 41831 24769 41843 24772
rect 41785 24763 41843 24769
rect 41874 24760 41880 24772
rect 41932 24760 41938 24812
rect 44174 24760 44180 24812
rect 44232 24800 44238 24812
rect 44269 24803 44327 24809
rect 44269 24800 44281 24803
rect 44232 24772 44281 24800
rect 44232 24760 44238 24772
rect 44269 24769 44281 24772
rect 44315 24769 44327 24803
rect 44542 24800 44548 24812
rect 44503 24772 44548 24800
rect 44269 24763 44327 24769
rect 44542 24760 44548 24772
rect 44600 24760 44606 24812
rect 44913 24803 44971 24809
rect 44913 24769 44925 24803
rect 44959 24800 44971 24803
rect 45370 24800 45376 24812
rect 44959 24772 45376 24800
rect 44959 24769 44971 24772
rect 44913 24763 44971 24769
rect 45370 24760 45376 24772
rect 45428 24760 45434 24812
rect 45738 24800 45744 24812
rect 45480 24772 45744 24800
rect 41693 24735 41751 24741
rect 41693 24701 41705 24735
rect 41739 24732 41751 24735
rect 42794 24732 42800 24744
rect 41739 24704 42800 24732
rect 41739 24701 41751 24704
rect 41693 24695 41751 24701
rect 42794 24692 42800 24704
rect 42852 24692 42858 24744
rect 45094 24732 45100 24744
rect 45055 24704 45100 24732
rect 45094 24692 45100 24704
rect 45152 24692 45158 24744
rect 34379 24636 40264 24664
rect 42812 24664 42840 24692
rect 45480 24664 45508 24772
rect 45738 24760 45744 24772
rect 45796 24760 45802 24812
rect 45830 24760 45836 24812
rect 45888 24800 45894 24812
rect 46032 24809 46060 24840
rect 46201 24837 46213 24871
rect 46247 24868 46259 24871
rect 47026 24868 47032 24880
rect 46247 24840 47032 24868
rect 46247 24837 46259 24840
rect 46201 24831 46259 24837
rect 47026 24828 47032 24840
rect 47084 24828 47090 24880
rect 52914 24828 52920 24880
rect 52972 24868 52978 24880
rect 55582 24868 55588 24880
rect 52972 24840 55588 24868
rect 52972 24828 52978 24840
rect 55582 24828 55588 24840
rect 55640 24868 55646 24880
rect 55784 24877 55812 24908
rect 57974 24896 57980 24908
rect 58032 24896 58038 24948
rect 55677 24871 55735 24877
rect 55677 24868 55689 24871
rect 55640 24840 55689 24868
rect 55640 24828 55646 24840
rect 55677 24837 55689 24840
rect 55723 24837 55735 24871
rect 55677 24831 55735 24837
rect 55769 24871 55827 24877
rect 55769 24837 55781 24871
rect 55815 24837 55827 24871
rect 55769 24831 55827 24837
rect 46017 24803 46075 24809
rect 45888 24772 45933 24800
rect 45888 24760 45894 24772
rect 46017 24769 46029 24803
rect 46063 24800 46075 24803
rect 46290 24800 46296 24812
rect 46063 24772 46296 24800
rect 46063 24769 46075 24772
rect 46017 24763 46075 24769
rect 46290 24760 46296 24772
rect 46348 24760 46354 24812
rect 50709 24803 50767 24809
rect 50709 24800 50721 24803
rect 49528 24772 50721 24800
rect 45646 24692 45652 24744
rect 45704 24732 45710 24744
rect 46106 24732 46112 24744
rect 45704 24704 46112 24732
rect 45704 24692 45710 24704
rect 46106 24692 46112 24704
rect 46164 24692 46170 24744
rect 42812 24636 45508 24664
rect 34379 24633 34391 24636
rect 34333 24627 34391 24633
rect 49528 24608 49556 24772
rect 50709 24769 50721 24772
rect 50755 24769 50767 24803
rect 50709 24763 50767 24769
rect 51074 24760 51080 24812
rect 51132 24800 51138 24812
rect 51132 24772 51177 24800
rect 51132 24760 51138 24772
rect 53190 24760 53196 24812
rect 53248 24800 53254 24812
rect 55398 24800 55404 24812
rect 53248 24772 55404 24800
rect 53248 24760 53254 24772
rect 55398 24760 55404 24772
rect 55456 24760 55462 24812
rect 55490 24760 55496 24812
rect 55548 24800 55554 24812
rect 55548 24772 55593 24800
rect 55548 24760 55554 24772
rect 55674 24692 55680 24744
rect 55732 24732 55738 24744
rect 55784 24732 55812 24831
rect 55858 24760 55864 24812
rect 55916 24800 55922 24812
rect 56873 24803 56931 24809
rect 55916 24772 55961 24800
rect 55916 24760 55922 24772
rect 56873 24769 56885 24803
rect 56919 24769 56931 24803
rect 56873 24763 56931 24769
rect 56888 24732 56916 24763
rect 56962 24760 56968 24812
rect 57020 24800 57026 24812
rect 57149 24803 57207 24809
rect 57020 24772 57065 24800
rect 57020 24760 57026 24772
rect 57149 24769 57161 24803
rect 57195 24769 57207 24803
rect 57149 24763 57207 24769
rect 57054 24732 57060 24744
rect 55732 24704 55812 24732
rect 56060 24704 57060 24732
rect 55732 24692 55738 24704
rect 56060 24673 56088 24704
rect 57054 24692 57060 24704
rect 57112 24692 57118 24744
rect 57164 24732 57192 24763
rect 57238 24760 57244 24812
rect 57296 24800 57302 24812
rect 57333 24803 57391 24809
rect 57333 24800 57345 24803
rect 57296 24772 57345 24800
rect 57296 24760 57302 24772
rect 57333 24769 57345 24772
rect 57379 24769 57391 24803
rect 57882 24800 57888 24812
rect 57843 24772 57888 24800
rect 57333 24763 57391 24769
rect 57882 24760 57888 24772
rect 57940 24760 57946 24812
rect 57977 24803 58035 24809
rect 57977 24769 57989 24803
rect 58023 24769 58035 24803
rect 57977 24763 58035 24769
rect 58161 24803 58219 24809
rect 58161 24769 58173 24803
rect 58207 24769 58219 24803
rect 58161 24763 58219 24769
rect 57900 24732 57928 24760
rect 57164 24704 57928 24732
rect 56045 24667 56103 24673
rect 56045 24633 56057 24667
rect 56091 24633 56103 24667
rect 56045 24627 56103 24633
rect 56962 24624 56968 24676
rect 57020 24664 57026 24676
rect 57992 24664 58020 24763
rect 57020 24636 58020 24664
rect 57020 24624 57026 24636
rect 3602 24596 3608 24608
rect 3563 24568 3608 24596
rect 3602 24556 3608 24568
rect 3660 24556 3666 24608
rect 7190 24556 7196 24608
rect 7248 24596 7254 24608
rect 8662 24596 8668 24608
rect 7248 24568 8668 24596
rect 7248 24556 7254 24568
rect 8662 24556 8668 24568
rect 8720 24556 8726 24608
rect 9674 24556 9680 24608
rect 9732 24596 9738 24608
rect 10413 24599 10471 24605
rect 10413 24596 10425 24599
rect 9732 24568 10425 24596
rect 9732 24556 9738 24568
rect 10413 24565 10425 24568
rect 10459 24565 10471 24599
rect 14090 24596 14096 24608
rect 14051 24568 14096 24596
rect 10413 24559 10471 24565
rect 14090 24556 14096 24568
rect 14148 24556 14154 24608
rect 15010 24556 15016 24608
rect 15068 24596 15074 24608
rect 16482 24596 16488 24608
rect 15068 24568 16488 24596
rect 15068 24556 15074 24568
rect 16482 24556 16488 24568
rect 16540 24596 16546 24608
rect 20070 24596 20076 24608
rect 16540 24568 20076 24596
rect 16540 24556 16546 24568
rect 20070 24556 20076 24568
rect 20128 24556 20134 24608
rect 20530 24556 20536 24608
rect 20588 24596 20594 24608
rect 20717 24599 20775 24605
rect 20717 24596 20729 24599
rect 20588 24568 20729 24596
rect 20588 24556 20594 24568
rect 20717 24565 20729 24568
rect 20763 24565 20775 24599
rect 28534 24596 28540 24608
rect 28495 24568 28540 24596
rect 20717 24559 20775 24565
rect 28534 24556 28540 24568
rect 28592 24556 28598 24608
rect 33226 24596 33232 24608
rect 33187 24568 33232 24596
rect 33226 24556 33232 24568
rect 33284 24556 33290 24608
rect 33870 24556 33876 24608
rect 33928 24596 33934 24608
rect 37366 24596 37372 24608
rect 33928 24568 37372 24596
rect 33928 24556 33934 24568
rect 37366 24556 37372 24568
rect 37424 24556 37430 24608
rect 37734 24596 37740 24608
rect 37695 24568 37740 24596
rect 37734 24556 37740 24568
rect 37792 24556 37798 24608
rect 38105 24599 38163 24605
rect 38105 24565 38117 24599
rect 38151 24596 38163 24599
rect 39942 24596 39948 24608
rect 38151 24568 39948 24596
rect 38151 24565 38163 24568
rect 38105 24559 38163 24565
rect 39942 24556 39948 24568
rect 40000 24556 40006 24608
rect 40954 24556 40960 24608
rect 41012 24596 41018 24608
rect 45830 24596 45836 24608
rect 41012 24568 45836 24596
rect 41012 24556 41018 24568
rect 45830 24556 45836 24568
rect 45888 24556 45894 24608
rect 49510 24596 49516 24608
rect 49471 24568 49516 24596
rect 49510 24556 49516 24568
rect 49568 24556 49574 24608
rect 57146 24556 57152 24608
rect 57204 24596 57210 24608
rect 58176 24596 58204 24763
rect 57204 24568 58204 24596
rect 57204 24556 57210 24568
rect 1104 24506 58880 24528
rect 1104 24454 4214 24506
rect 4266 24454 4278 24506
rect 4330 24454 4342 24506
rect 4394 24454 4406 24506
rect 4458 24454 4470 24506
rect 4522 24454 34934 24506
rect 34986 24454 34998 24506
rect 35050 24454 35062 24506
rect 35114 24454 35126 24506
rect 35178 24454 35190 24506
rect 35242 24454 58880 24506
rect 1104 24432 58880 24454
rect 3878 24392 3884 24404
rect 3839 24364 3884 24392
rect 3878 24352 3884 24364
rect 3936 24352 3942 24404
rect 7745 24395 7803 24401
rect 7745 24361 7757 24395
rect 7791 24392 7803 24395
rect 8202 24392 8208 24404
rect 7791 24364 8208 24392
rect 7791 24361 7803 24364
rect 7745 24355 7803 24361
rect 8202 24352 8208 24364
rect 8260 24392 8266 24404
rect 8386 24392 8392 24404
rect 8260 24364 8392 24392
rect 8260 24352 8266 24364
rect 8386 24352 8392 24364
rect 8444 24352 8450 24404
rect 10689 24395 10747 24401
rect 10689 24361 10701 24395
rect 10735 24392 10747 24395
rect 10870 24392 10876 24404
rect 10735 24364 10876 24392
rect 10735 24361 10747 24364
rect 10689 24355 10747 24361
rect 10870 24352 10876 24364
rect 10928 24352 10934 24404
rect 12802 24352 12808 24404
rect 12860 24392 12866 24404
rect 13081 24395 13139 24401
rect 13081 24392 13093 24395
rect 12860 24364 13093 24392
rect 12860 24352 12866 24364
rect 13081 24361 13093 24364
rect 13127 24392 13139 24395
rect 17034 24392 17040 24404
rect 13127 24364 17040 24392
rect 13127 24361 13139 24364
rect 13081 24355 13139 24361
rect 17034 24352 17040 24364
rect 17092 24352 17098 24404
rect 17954 24392 17960 24404
rect 17915 24364 17960 24392
rect 17954 24352 17960 24364
rect 18012 24352 18018 24404
rect 20714 24392 20720 24404
rect 19812 24364 20720 24392
rect 7650 24284 7656 24336
rect 7708 24324 7714 24336
rect 13265 24327 13323 24333
rect 13265 24324 13277 24327
rect 7708 24296 13277 24324
rect 7708 24284 7714 24296
rect 13265 24293 13277 24296
rect 13311 24324 13323 24327
rect 13354 24324 13360 24336
rect 13311 24296 13360 24324
rect 13311 24293 13323 24296
rect 13265 24287 13323 24293
rect 13354 24284 13360 24296
rect 13412 24284 13418 24336
rect 14734 24324 14740 24336
rect 14695 24296 14740 24324
rect 14734 24284 14740 24296
rect 14792 24284 14798 24336
rect 14844 24296 17632 24324
rect 11532 24228 14366 24256
rect 6914 24148 6920 24200
rect 6972 24188 6978 24200
rect 7561 24191 7619 24197
rect 7561 24188 7573 24191
rect 6972 24160 7573 24188
rect 6972 24148 6978 24160
rect 7561 24157 7573 24160
rect 7607 24188 7619 24191
rect 8297 24191 8355 24197
rect 8297 24188 8309 24191
rect 7607 24160 8309 24188
rect 7607 24157 7619 24160
rect 7561 24151 7619 24157
rect 8297 24157 8309 24160
rect 8343 24188 8355 24191
rect 8386 24188 8392 24200
rect 8343 24160 8392 24188
rect 8343 24157 8355 24160
rect 8297 24151 8355 24157
rect 8386 24148 8392 24160
rect 8444 24148 8450 24200
rect 9214 24148 9220 24200
rect 9272 24188 9278 24200
rect 10137 24191 10195 24197
rect 10137 24188 10149 24191
rect 9272 24160 10149 24188
rect 9272 24148 9278 24160
rect 10137 24157 10149 24160
rect 10183 24157 10195 24191
rect 10137 24151 10195 24157
rect 10229 24191 10287 24197
rect 10229 24157 10241 24191
rect 10275 24188 10287 24191
rect 10318 24188 10324 24200
rect 10275 24160 10324 24188
rect 10275 24157 10287 24160
rect 10229 24151 10287 24157
rect 10318 24148 10324 24160
rect 10376 24148 10382 24200
rect 11532 24197 11560 24228
rect 10413 24191 10471 24197
rect 10413 24157 10425 24191
rect 10459 24157 10471 24191
rect 10413 24151 10471 24157
rect 10505 24191 10563 24197
rect 10505 24157 10517 24191
rect 10551 24188 10563 24191
rect 11517 24191 11575 24197
rect 11517 24188 11529 24191
rect 10551 24160 11529 24188
rect 10551 24157 10563 24160
rect 10505 24151 10563 24157
rect 11517 24157 11529 24160
rect 11563 24157 11575 24191
rect 11517 24151 11575 24157
rect 9306 24080 9312 24132
rect 9364 24120 9370 24132
rect 9401 24123 9459 24129
rect 9401 24120 9413 24123
rect 9364 24092 9413 24120
rect 9364 24080 9370 24092
rect 9401 24089 9413 24092
rect 9447 24089 9459 24123
rect 9401 24083 9459 24089
rect 9585 24123 9643 24129
rect 9585 24089 9597 24123
rect 9631 24120 9643 24123
rect 9766 24120 9772 24132
rect 9631 24092 9772 24120
rect 9631 24089 9643 24092
rect 9585 24083 9643 24089
rect 9766 24080 9772 24092
rect 9824 24080 9830 24132
rect 10428 24120 10456 24151
rect 12986 24148 12992 24200
rect 13044 24188 13050 24200
rect 14093 24191 14151 24197
rect 14093 24188 14105 24191
rect 13044 24160 14105 24188
rect 13044 24148 13050 24160
rect 14093 24157 14105 24160
rect 14139 24157 14151 24191
rect 14093 24151 14151 24157
rect 14182 24148 14188 24200
rect 14240 24188 14246 24200
rect 14338 24188 14366 24228
rect 14642 24216 14648 24268
rect 14700 24256 14706 24268
rect 14844 24256 14872 24296
rect 16482 24256 16488 24268
rect 14700 24228 14872 24256
rect 16316 24228 16488 24256
rect 14700 24216 14706 24228
rect 14458 24188 14464 24200
rect 14240 24160 14285 24188
rect 14338 24160 14464 24188
rect 14240 24148 14246 24160
rect 14458 24148 14464 24160
rect 14516 24148 14522 24200
rect 14550 24148 14556 24200
rect 14608 24197 14614 24200
rect 16316 24197 16344 24228
rect 16482 24216 16488 24228
rect 16540 24216 16546 24268
rect 17604 24256 17632 24296
rect 18601 24259 18659 24265
rect 18601 24256 18613 24259
rect 17604 24228 18613 24256
rect 14608 24188 14616 24197
rect 16301 24191 16359 24197
rect 14608 24160 14653 24188
rect 14608 24151 14616 24160
rect 16301 24157 16313 24191
rect 16347 24157 16359 24191
rect 16574 24188 16580 24200
rect 16301 24151 16359 24157
rect 16408 24160 16580 24188
rect 14608 24148 14614 24151
rect 10778 24120 10784 24132
rect 10428 24092 10784 24120
rect 10778 24080 10784 24092
rect 10836 24080 10842 24132
rect 11333 24123 11391 24129
rect 11333 24089 11345 24123
rect 11379 24120 11391 24123
rect 13538 24120 13544 24132
rect 11379 24092 12434 24120
rect 13499 24092 13544 24120
rect 11379 24089 11391 24092
rect 11333 24083 11391 24089
rect 12406 24052 12434 24092
rect 13538 24080 13544 24092
rect 13596 24080 13602 24132
rect 14369 24123 14427 24129
rect 14369 24120 14381 24123
rect 14108 24092 14381 24120
rect 14108 24064 14136 24092
rect 14369 24089 14381 24092
rect 14415 24089 14427 24123
rect 14476 24120 14504 24148
rect 16408 24120 16436 24160
rect 16574 24148 16580 24160
rect 16632 24148 16638 24200
rect 16669 24191 16727 24197
rect 16669 24157 16681 24191
rect 16715 24188 16727 24191
rect 16758 24188 16764 24200
rect 16715 24160 16764 24188
rect 16715 24157 16727 24160
rect 16669 24151 16727 24157
rect 16758 24148 16764 24160
rect 16816 24148 16822 24200
rect 17218 24148 17224 24200
rect 17276 24188 17282 24200
rect 17313 24191 17371 24197
rect 17313 24188 17325 24191
rect 17276 24160 17325 24188
rect 17276 24148 17282 24160
rect 17313 24157 17325 24160
rect 17359 24157 17371 24191
rect 17313 24151 17371 24157
rect 17402 24148 17408 24200
rect 17460 24188 17466 24200
rect 17460 24160 17553 24188
rect 17460 24148 17466 24160
rect 14476 24092 16436 24120
rect 14369 24083 14427 24089
rect 16482 24080 16488 24132
rect 16540 24120 16546 24132
rect 17420 24120 17448 24148
rect 17604 24129 17632 24228
rect 18601 24225 18613 24228
rect 18647 24256 18659 24259
rect 19058 24256 19064 24268
rect 18647 24228 19064 24256
rect 18647 24225 18659 24228
rect 18601 24219 18659 24225
rect 19058 24216 19064 24228
rect 19116 24216 19122 24268
rect 17770 24148 17776 24200
rect 17828 24197 17834 24200
rect 17828 24188 17836 24197
rect 17828 24160 17873 24188
rect 17828 24151 17836 24160
rect 17828 24148 17834 24151
rect 18506 24148 18512 24200
rect 18564 24188 18570 24200
rect 19812 24197 19840 24364
rect 20714 24352 20720 24364
rect 20772 24352 20778 24404
rect 21450 24392 21456 24404
rect 21411 24364 21456 24392
rect 21450 24352 21456 24364
rect 21508 24352 21514 24404
rect 24946 24392 24952 24404
rect 21560 24364 24952 24392
rect 20349 24327 20407 24333
rect 20349 24293 20361 24327
rect 20395 24293 20407 24327
rect 20349 24287 20407 24293
rect 19797 24191 19855 24197
rect 19797 24188 19809 24191
rect 18564 24160 19809 24188
rect 18564 24148 18570 24160
rect 19797 24157 19809 24160
rect 19843 24157 19855 24191
rect 20070 24188 20076 24200
rect 20031 24160 20076 24188
rect 19797 24151 19855 24157
rect 20070 24148 20076 24160
rect 20128 24148 20134 24200
rect 20162 24148 20168 24200
rect 20220 24188 20226 24200
rect 20364 24188 20392 24287
rect 21560 24256 21588 24364
rect 24946 24352 24952 24364
rect 25004 24352 25010 24404
rect 25130 24392 25136 24404
rect 25091 24364 25136 24392
rect 25130 24352 25136 24364
rect 25188 24352 25194 24404
rect 25590 24352 25596 24404
rect 25648 24392 25654 24404
rect 27706 24392 27712 24404
rect 25648 24364 27292 24392
rect 27667 24364 27712 24392
rect 25648 24352 25654 24364
rect 23382 24284 23388 24336
rect 23440 24324 23446 24336
rect 27157 24327 27215 24333
rect 27157 24324 27169 24327
rect 23440 24296 27169 24324
rect 23440 24284 23446 24296
rect 27157 24293 27169 24296
rect 27203 24293 27215 24327
rect 27264 24324 27292 24364
rect 27706 24352 27712 24364
rect 27764 24352 27770 24404
rect 27798 24352 27804 24404
rect 27856 24392 27862 24404
rect 27893 24395 27951 24401
rect 27893 24392 27905 24395
rect 27856 24364 27905 24392
rect 27856 24352 27862 24364
rect 27893 24361 27905 24364
rect 27939 24361 27951 24395
rect 27893 24355 27951 24361
rect 28537 24395 28595 24401
rect 28537 24361 28549 24395
rect 28583 24392 28595 24395
rect 28718 24392 28724 24404
rect 28583 24364 28724 24392
rect 28583 24361 28595 24364
rect 28537 24355 28595 24361
rect 28718 24352 28724 24364
rect 28776 24352 28782 24404
rect 31110 24392 31116 24404
rect 31071 24364 31116 24392
rect 31110 24352 31116 24364
rect 31168 24352 31174 24404
rect 33962 24392 33968 24404
rect 33923 24364 33968 24392
rect 33962 24352 33968 24364
rect 34020 24352 34026 24404
rect 38197 24395 38255 24401
rect 38197 24392 38209 24395
rect 37292 24364 38209 24392
rect 27264 24296 31754 24324
rect 27157 24287 27215 24293
rect 21192 24228 21588 24256
rect 20809 24191 20867 24197
rect 20809 24188 20821 24191
rect 20220 24160 20265 24188
rect 20364 24160 20821 24188
rect 20220 24148 20226 24160
rect 20809 24157 20821 24160
rect 20855 24157 20867 24191
rect 20809 24151 20867 24157
rect 20898 24148 20904 24200
rect 20956 24197 20962 24200
rect 20956 24191 21015 24197
rect 20956 24157 20969 24191
rect 21003 24188 21015 24191
rect 21192 24188 21220 24228
rect 23658 24216 23664 24268
rect 23716 24256 23722 24268
rect 24762 24256 24768 24268
rect 23716 24228 24768 24256
rect 23716 24216 23722 24228
rect 24762 24216 24768 24228
rect 24820 24256 24826 24268
rect 24820 24228 24900 24256
rect 24820 24216 24826 24228
rect 21003 24160 21220 24188
rect 21315 24191 21373 24197
rect 21003 24157 21015 24160
rect 20956 24151 21015 24157
rect 21315 24157 21327 24191
rect 21361 24188 21373 24191
rect 21450 24188 21456 24200
rect 21361 24160 21456 24188
rect 21361 24157 21373 24160
rect 21315 24151 21373 24157
rect 20956 24148 20962 24151
rect 21450 24148 21456 24160
rect 21508 24148 21514 24200
rect 23477 24191 23535 24197
rect 23477 24157 23489 24191
rect 23523 24188 23535 24191
rect 23566 24188 23572 24200
rect 23523 24160 23572 24188
rect 23523 24157 23535 24160
rect 23477 24151 23535 24157
rect 23566 24148 23572 24160
rect 23624 24148 23630 24200
rect 24486 24188 24492 24200
rect 24447 24160 24492 24188
rect 24486 24148 24492 24160
rect 24544 24148 24550 24200
rect 24578 24148 24584 24200
rect 24636 24188 24642 24200
rect 24872 24197 24900 24228
rect 25038 24197 25044 24200
rect 24857 24191 24915 24197
rect 24636 24160 24681 24188
rect 24636 24148 24642 24160
rect 24857 24157 24869 24191
rect 24903 24157 24915 24191
rect 24857 24151 24915 24157
rect 24995 24191 25044 24197
rect 24995 24157 25007 24191
rect 25041 24157 25044 24191
rect 24995 24151 25044 24157
rect 25038 24148 25044 24151
rect 25096 24148 25102 24200
rect 16540 24092 16585 24120
rect 16776 24092 17448 24120
rect 17589 24123 17647 24129
rect 16540 24080 16546 24092
rect 13262 24052 13268 24064
rect 12406 24024 13268 24052
rect 13262 24012 13268 24024
rect 13320 24052 13326 24064
rect 13814 24052 13820 24064
rect 13320 24024 13820 24052
rect 13320 24012 13326 24024
rect 13814 24012 13820 24024
rect 13872 24012 13878 24064
rect 14090 24012 14096 24064
rect 14148 24012 14154 24064
rect 14182 24012 14188 24064
rect 14240 24052 14246 24064
rect 16776 24052 16804 24092
rect 17589 24089 17601 24123
rect 17635 24089 17647 24123
rect 17589 24083 17647 24089
rect 17681 24123 17739 24129
rect 17681 24089 17693 24123
rect 17727 24120 17739 24123
rect 19978 24120 19984 24132
rect 17727 24092 19840 24120
rect 19939 24092 19984 24120
rect 17727 24089 17739 24092
rect 17681 24083 17739 24089
rect 14240 24024 16804 24052
rect 16853 24055 16911 24061
rect 14240 24012 14246 24024
rect 16853 24021 16865 24055
rect 16899 24052 16911 24055
rect 17862 24052 17868 24064
rect 16899 24024 17868 24052
rect 16899 24021 16911 24024
rect 16853 24015 16911 24021
rect 17862 24012 17868 24024
rect 17920 24012 17926 24064
rect 19812 24052 19840 24092
rect 19978 24080 19984 24092
rect 20036 24080 20042 24132
rect 20438 24080 20444 24132
rect 20496 24120 20502 24132
rect 20916 24120 20944 24148
rect 21085 24123 21143 24129
rect 21085 24120 21097 24123
rect 20496 24092 20944 24120
rect 21008 24092 21097 24120
rect 20496 24080 20502 24092
rect 21008 24064 21036 24092
rect 21085 24089 21097 24092
rect 21131 24089 21143 24123
rect 21085 24083 21143 24089
rect 21174 24080 21180 24132
rect 21232 24120 21238 24132
rect 21232 24092 21277 24120
rect 21232 24080 21238 24092
rect 23014 24080 23020 24132
rect 23072 24120 23078 24132
rect 23934 24120 23940 24132
rect 23072 24092 23940 24120
rect 23072 24080 23078 24092
rect 23934 24080 23940 24092
rect 23992 24080 23998 24132
rect 24765 24123 24823 24129
rect 24765 24089 24777 24123
rect 24811 24089 24823 24123
rect 27172 24120 27200 24287
rect 28534 24188 28540 24200
rect 27908 24160 28540 24188
rect 27908 24129 27936 24160
rect 28534 24148 28540 24160
rect 28592 24148 28598 24200
rect 28810 24188 28816 24200
rect 28771 24160 28816 24188
rect 28810 24148 28816 24160
rect 28868 24188 28874 24200
rect 30377 24191 30435 24197
rect 30377 24188 30389 24191
rect 28868 24160 30389 24188
rect 28868 24148 28874 24160
rect 30377 24157 30389 24160
rect 30423 24157 30435 24191
rect 30377 24151 30435 24157
rect 27861 24123 27936 24129
rect 27861 24120 27873 24123
rect 27172 24092 27873 24120
rect 24765 24083 24823 24089
rect 27861 24089 27873 24092
rect 27907 24092 27936 24123
rect 28077 24123 28135 24129
rect 27907 24089 27919 24092
rect 27861 24083 27919 24089
rect 28077 24089 28089 24123
rect 28123 24089 28135 24123
rect 30392 24120 30420 24151
rect 30929 24123 30987 24129
rect 30929 24120 30941 24123
rect 30392 24092 30941 24120
rect 28077 24083 28135 24089
rect 30929 24089 30941 24092
rect 30975 24089 30987 24123
rect 31726 24120 31754 24296
rect 33413 24191 33471 24197
rect 33413 24157 33425 24191
rect 33459 24188 33471 24191
rect 33870 24188 33876 24200
rect 33459 24160 33876 24188
rect 33459 24157 33471 24160
rect 33413 24151 33471 24157
rect 33870 24148 33876 24160
rect 33928 24148 33934 24200
rect 33980 24188 34008 24352
rect 37292 24197 37320 24364
rect 38197 24361 38209 24364
rect 38243 24361 38255 24395
rect 38562 24392 38568 24404
rect 38523 24364 38568 24392
rect 38197 24355 38255 24361
rect 38562 24352 38568 24364
rect 38620 24352 38626 24404
rect 39114 24392 39120 24404
rect 39075 24364 39120 24392
rect 39114 24352 39120 24364
rect 39172 24352 39178 24404
rect 39209 24395 39267 24401
rect 39209 24361 39221 24395
rect 39255 24392 39267 24395
rect 40218 24392 40224 24404
rect 39255 24364 40224 24392
rect 39255 24361 39267 24364
rect 39209 24355 39267 24361
rect 40218 24352 40224 24364
rect 40276 24352 40282 24404
rect 42245 24395 42303 24401
rect 42245 24361 42257 24395
rect 42291 24392 42303 24395
rect 44542 24392 44548 24404
rect 42291 24364 44548 24392
rect 42291 24361 42303 24364
rect 42245 24355 42303 24361
rect 44542 24352 44548 24364
rect 44600 24352 44606 24404
rect 45646 24392 45652 24404
rect 45607 24364 45652 24392
rect 45646 24352 45652 24364
rect 45704 24352 45710 24404
rect 55490 24352 55496 24404
rect 55548 24392 55554 24404
rect 56321 24395 56379 24401
rect 56321 24392 56333 24395
rect 55548 24364 56333 24392
rect 55548 24352 55554 24364
rect 56321 24361 56333 24364
rect 56367 24361 56379 24395
rect 56321 24355 56379 24361
rect 37642 24324 37648 24336
rect 37603 24296 37648 24324
rect 37642 24284 37648 24296
rect 37700 24284 37706 24336
rect 37369 24259 37427 24265
rect 37369 24225 37381 24259
rect 37415 24225 37427 24259
rect 38580 24256 38608 24352
rect 41417 24327 41475 24333
rect 41417 24293 41429 24327
rect 41463 24324 41475 24327
rect 43806 24324 43812 24336
rect 41463 24296 43812 24324
rect 41463 24293 41475 24296
rect 41417 24287 41475 24293
rect 43806 24284 43812 24296
rect 43864 24284 43870 24336
rect 43901 24327 43959 24333
rect 43901 24293 43913 24327
rect 43947 24293 43959 24327
rect 43901 24287 43959 24293
rect 39301 24259 39359 24265
rect 39301 24256 39313 24259
rect 38580 24228 39313 24256
rect 37369 24219 37427 24225
rect 39301 24225 39313 24228
rect 39347 24225 39359 24259
rect 39301 24219 39359 24225
rect 34701 24191 34759 24197
rect 34701 24188 34713 24191
rect 33980 24160 34713 24188
rect 34701 24157 34713 24160
rect 34747 24157 34759 24191
rect 37277 24191 37335 24197
rect 37277 24188 37289 24191
rect 34701 24151 34759 24157
rect 34900 24160 37289 24188
rect 34900 24120 34928 24160
rect 37277 24157 37289 24160
rect 37323 24157 37335 24191
rect 37384 24188 37412 24219
rect 40586 24216 40592 24268
rect 40644 24256 40650 24268
rect 40957 24259 41015 24265
rect 40957 24256 40969 24259
rect 40644 24228 40969 24256
rect 40644 24216 40650 24228
rect 40957 24225 40969 24228
rect 41003 24256 41015 24259
rect 43916 24256 43944 24287
rect 45094 24256 45100 24268
rect 41003 24228 42196 24256
rect 43916 24228 45100 24256
rect 41003 24225 41015 24228
rect 40957 24219 41015 24225
rect 38102 24188 38108 24200
rect 37384 24160 38108 24188
rect 37277 24151 37335 24157
rect 38102 24148 38108 24160
rect 38160 24148 38166 24200
rect 39025 24191 39083 24197
rect 39025 24157 39037 24191
rect 39071 24157 39083 24191
rect 41046 24188 41052 24200
rect 41007 24160 41052 24188
rect 39025 24151 39083 24157
rect 31726 24092 34928 24120
rect 34977 24123 35035 24129
rect 30929 24083 30987 24089
rect 34977 24089 34989 24123
rect 35023 24089 35035 24123
rect 34977 24083 35035 24089
rect 20254 24052 20260 24064
rect 19812 24024 20260 24052
rect 20254 24012 20260 24024
rect 20312 24012 20318 24064
rect 20990 24012 20996 24064
rect 21048 24012 21054 24064
rect 21358 24012 21364 24064
rect 21416 24052 21422 24064
rect 22005 24055 22063 24061
rect 22005 24052 22017 24055
rect 21416 24024 22017 24052
rect 21416 24012 21422 24024
rect 22005 24021 22017 24024
rect 22051 24021 22063 24055
rect 22005 24015 22063 24021
rect 22738 24012 22744 24064
rect 22796 24052 22802 24064
rect 23569 24055 23627 24061
rect 23569 24052 23581 24055
rect 22796 24024 23581 24052
rect 22796 24012 22802 24024
rect 23569 24021 23581 24024
rect 23615 24021 23627 24055
rect 23569 24015 23627 24021
rect 24578 24012 24584 24064
rect 24636 24052 24642 24064
rect 24780 24052 24808 24083
rect 25958 24052 25964 24064
rect 24636 24024 25964 24052
rect 24636 24012 24642 24024
rect 25958 24012 25964 24024
rect 26016 24012 26022 24064
rect 28092 24052 28120 24083
rect 28721 24055 28779 24061
rect 28721 24052 28733 24055
rect 28092 24024 28733 24052
rect 28721 24021 28733 24024
rect 28767 24052 28779 24055
rect 29454 24052 29460 24064
rect 28767 24024 29460 24052
rect 28767 24021 28779 24024
rect 28721 24015 28779 24021
rect 29454 24012 29460 24024
rect 29512 24012 29518 24064
rect 29638 24012 29644 24064
rect 29696 24052 29702 24064
rect 29825 24055 29883 24061
rect 29825 24052 29837 24055
rect 29696 24024 29837 24052
rect 29696 24012 29702 24024
rect 29825 24021 29837 24024
rect 29871 24052 29883 24055
rect 31113 24055 31171 24061
rect 31113 24052 31125 24055
rect 29871 24024 31125 24052
rect 29871 24021 29883 24024
rect 29825 24015 29883 24021
rect 31113 24021 31125 24024
rect 31159 24021 31171 24055
rect 31294 24052 31300 24064
rect 31255 24024 31300 24052
rect 31113 24015 31171 24021
rect 31294 24012 31300 24024
rect 31352 24012 31358 24064
rect 33778 24012 33784 24064
rect 33836 24052 33842 24064
rect 34330 24052 34336 24064
rect 33836 24024 34336 24052
rect 33836 24012 33842 24024
rect 34330 24012 34336 24024
rect 34388 24052 34394 24064
rect 34992 24052 35020 24083
rect 37734 24080 37740 24132
rect 37792 24120 37798 24132
rect 39040 24120 39068 24151
rect 41046 24148 41052 24160
rect 41104 24188 41110 24200
rect 42061 24191 42119 24197
rect 42061 24188 42073 24191
rect 41104 24160 42073 24188
rect 41104 24148 41110 24160
rect 42061 24157 42073 24160
rect 42107 24157 42119 24191
rect 42061 24151 42119 24157
rect 37792 24092 39068 24120
rect 41877 24123 41935 24129
rect 37792 24080 37798 24092
rect 41877 24089 41889 24123
rect 41923 24120 41935 24123
rect 42168 24120 42196 24228
rect 45094 24216 45100 24228
rect 45152 24256 45158 24268
rect 48869 24259 48927 24265
rect 45152 24228 45324 24256
rect 45152 24216 45158 24228
rect 43625 24191 43683 24197
rect 43625 24157 43637 24191
rect 43671 24188 43683 24191
rect 43806 24188 43812 24200
rect 43671 24160 43812 24188
rect 43671 24157 43683 24160
rect 43625 24151 43683 24157
rect 43806 24148 43812 24160
rect 43864 24148 43870 24200
rect 44174 24148 44180 24200
rect 44232 24188 44238 24200
rect 45296 24197 45324 24228
rect 48869 24225 48881 24259
rect 48915 24256 48927 24259
rect 49234 24256 49240 24268
rect 48915 24228 49240 24256
rect 48915 24225 48927 24228
rect 48869 24219 48927 24225
rect 49234 24216 49240 24228
rect 49292 24216 49298 24268
rect 52822 24216 52828 24268
rect 52880 24256 52886 24268
rect 53101 24259 53159 24265
rect 53101 24256 53113 24259
rect 52880 24228 53113 24256
rect 52880 24216 52886 24228
rect 53101 24225 53113 24228
rect 53147 24225 53159 24259
rect 53101 24219 53159 24225
rect 57882 24216 57888 24268
rect 57940 24256 57946 24268
rect 57940 24228 58204 24256
rect 57940 24216 57946 24228
rect 45005 24191 45063 24197
rect 45005 24188 45017 24191
rect 44232 24160 45017 24188
rect 44232 24148 44238 24160
rect 45005 24157 45017 24160
rect 45051 24157 45063 24191
rect 45005 24151 45063 24157
rect 45189 24191 45247 24197
rect 45189 24157 45201 24191
rect 45235 24157 45247 24191
rect 45189 24151 45247 24157
rect 45281 24191 45339 24197
rect 45281 24157 45293 24191
rect 45327 24157 45339 24191
rect 45281 24151 45339 24157
rect 41923 24092 42196 24120
rect 43901 24123 43959 24129
rect 41923 24089 41935 24092
rect 41877 24083 41935 24089
rect 43901 24089 43913 24123
rect 43947 24120 43959 24123
rect 43990 24120 43996 24132
rect 43947 24092 43996 24120
rect 43947 24089 43959 24092
rect 43901 24083 43959 24089
rect 43990 24080 43996 24092
rect 44048 24080 44054 24132
rect 44542 24080 44548 24132
rect 44600 24120 44606 24132
rect 45204 24120 45232 24151
rect 45370 24148 45376 24200
rect 45428 24188 45434 24200
rect 47854 24188 47860 24200
rect 45428 24160 45473 24188
rect 47815 24160 47860 24188
rect 45428 24148 45434 24160
rect 47854 24148 47860 24160
rect 47912 24148 47918 24200
rect 48038 24188 48044 24200
rect 47999 24160 48044 24188
rect 48038 24148 48044 24160
rect 48096 24148 48102 24200
rect 52270 24148 52276 24200
rect 52328 24188 52334 24200
rect 52641 24191 52699 24197
rect 52641 24188 52653 24191
rect 52328 24160 52653 24188
rect 52328 24148 52334 24160
rect 52641 24157 52653 24160
rect 52687 24157 52699 24191
rect 52641 24151 52699 24157
rect 52730 24148 52736 24200
rect 52788 24188 52794 24200
rect 52917 24191 52975 24197
rect 52917 24188 52929 24191
rect 52788 24160 52929 24188
rect 52788 24148 52794 24160
rect 52917 24157 52929 24160
rect 52963 24157 52975 24191
rect 52917 24151 52975 24157
rect 53285 24191 53343 24197
rect 53285 24157 53297 24191
rect 53331 24188 53343 24191
rect 53650 24188 53656 24200
rect 53331 24160 53656 24188
rect 53331 24157 53343 24160
rect 53285 24151 53343 24157
rect 53650 24148 53656 24160
rect 53708 24148 53714 24200
rect 55306 24188 55312 24200
rect 55267 24160 55312 24188
rect 55306 24148 55312 24160
rect 55364 24148 55370 24200
rect 55398 24148 55404 24200
rect 55456 24188 55462 24200
rect 55582 24188 55588 24200
rect 55456 24160 55501 24188
rect 55543 24160 55588 24188
rect 55456 24148 55462 24160
rect 55582 24148 55588 24160
rect 55640 24148 55646 24200
rect 55674 24148 55680 24200
rect 55732 24188 55738 24200
rect 58176 24197 58204 24228
rect 58161 24191 58219 24197
rect 55732 24160 55777 24188
rect 55732 24148 55738 24160
rect 58161 24157 58173 24191
rect 58207 24157 58219 24191
rect 58161 24151 58219 24157
rect 44600 24092 45232 24120
rect 55324 24120 55352 24148
rect 56505 24123 56563 24129
rect 56505 24120 56517 24123
rect 55324 24092 56517 24120
rect 44600 24080 44606 24092
rect 56505 24089 56517 24092
rect 56551 24089 56563 24123
rect 56686 24120 56692 24132
rect 56647 24092 56692 24120
rect 56505 24083 56563 24089
rect 56686 24080 56692 24092
rect 56744 24080 56750 24132
rect 56778 24080 56784 24132
rect 56836 24120 56842 24132
rect 57885 24123 57943 24129
rect 57885 24120 57897 24123
rect 56836 24092 57897 24120
rect 56836 24080 56842 24092
rect 57885 24089 57897 24092
rect 57931 24089 57943 24123
rect 57885 24083 57943 24089
rect 34388 24024 35020 24052
rect 34388 24012 34394 24024
rect 37366 24012 37372 24064
rect 37424 24052 37430 24064
rect 38378 24052 38384 24064
rect 37424 24024 38384 24052
rect 37424 24012 37430 24024
rect 38378 24012 38384 24024
rect 38436 24012 38442 24064
rect 43530 24012 43536 24064
rect 43588 24052 43594 24064
rect 43717 24055 43775 24061
rect 43717 24052 43729 24055
rect 43588 24024 43729 24052
rect 43588 24012 43594 24024
rect 43717 24021 43729 24024
rect 43763 24021 43775 24055
rect 43717 24015 43775 24021
rect 55861 24055 55919 24061
rect 55861 24021 55873 24055
rect 55907 24052 55919 24055
rect 56318 24052 56324 24064
rect 55907 24024 56324 24052
rect 55907 24021 55919 24024
rect 55861 24015 55919 24021
rect 56318 24012 56324 24024
rect 56376 24012 56382 24064
rect 1104 23962 58880 23984
rect 1104 23910 19574 23962
rect 19626 23910 19638 23962
rect 19690 23910 19702 23962
rect 19754 23910 19766 23962
rect 19818 23910 19830 23962
rect 19882 23910 50294 23962
rect 50346 23910 50358 23962
rect 50410 23910 50422 23962
rect 50474 23910 50486 23962
rect 50538 23910 50550 23962
rect 50602 23910 58880 23962
rect 1104 23888 58880 23910
rect 7009 23851 7067 23857
rect 7009 23817 7021 23851
rect 7055 23817 7067 23851
rect 9398 23848 9404 23860
rect 9359 23820 9404 23848
rect 7009 23811 7067 23817
rect 2590 23780 2596 23792
rect 2240 23752 2596 23780
rect 2240 23721 2268 23752
rect 2590 23740 2596 23752
rect 2648 23740 2654 23792
rect 3881 23783 3939 23789
rect 3881 23749 3893 23783
rect 3927 23780 3939 23783
rect 4062 23780 4068 23792
rect 3927 23752 4068 23780
rect 3927 23749 3939 23752
rect 3881 23743 3939 23749
rect 4062 23740 4068 23752
rect 4120 23740 4126 23792
rect 7024 23780 7052 23811
rect 9398 23808 9404 23820
rect 9456 23808 9462 23860
rect 10318 23848 10324 23860
rect 10279 23820 10324 23848
rect 10318 23808 10324 23820
rect 10376 23808 10382 23860
rect 10778 23848 10784 23860
rect 10739 23820 10784 23848
rect 10778 23808 10784 23820
rect 10836 23808 10842 23860
rect 12802 23808 12808 23860
rect 12860 23808 12866 23860
rect 13817 23851 13875 23857
rect 13817 23817 13829 23851
rect 13863 23848 13875 23851
rect 14550 23848 14556 23860
rect 13863 23820 14556 23848
rect 13863 23817 13875 23820
rect 13817 23811 13875 23817
rect 14550 23808 14556 23820
rect 14608 23808 14614 23860
rect 17218 23848 17224 23860
rect 17179 23820 17224 23848
rect 17218 23808 17224 23820
rect 17276 23808 17282 23860
rect 18049 23851 18107 23857
rect 18049 23817 18061 23851
rect 18095 23848 18107 23851
rect 18138 23848 18144 23860
rect 18095 23820 18144 23848
rect 18095 23817 18107 23820
rect 18049 23811 18107 23817
rect 18138 23808 18144 23820
rect 18196 23848 18202 23860
rect 19242 23848 19248 23860
rect 18196 23820 19248 23848
rect 18196 23808 18202 23820
rect 19242 23808 19248 23820
rect 19300 23808 19306 23860
rect 19334 23808 19340 23860
rect 19392 23848 19398 23860
rect 19705 23851 19763 23857
rect 19705 23848 19717 23851
rect 19392 23820 19717 23848
rect 19392 23808 19398 23820
rect 19705 23817 19717 23820
rect 19751 23817 19763 23851
rect 19705 23811 19763 23817
rect 20162 23808 20168 23860
rect 20220 23848 20226 23860
rect 20346 23848 20352 23860
rect 20220 23820 20352 23848
rect 20220 23808 20226 23820
rect 20346 23808 20352 23820
rect 20404 23808 20410 23860
rect 20530 23808 20536 23860
rect 20588 23848 20594 23860
rect 20588 23820 20668 23848
rect 20588 23808 20594 23820
rect 7650 23780 7656 23792
rect 7024 23752 7656 23780
rect 2225 23715 2283 23721
rect 2225 23681 2237 23715
rect 2271 23681 2283 23715
rect 2498 23712 2504 23724
rect 2459 23684 2504 23712
rect 2225 23675 2283 23681
rect 2498 23672 2504 23684
rect 2556 23672 2562 23724
rect 5442 23712 5448 23724
rect 5403 23684 5448 23712
rect 5442 23672 5448 23684
rect 5500 23672 5506 23724
rect 7576 23721 7604 23752
rect 7650 23740 7656 23752
rect 7708 23740 7714 23792
rect 9950 23780 9956 23792
rect 9911 23752 9956 23780
rect 9950 23740 9956 23752
rect 10008 23740 10014 23792
rect 10183 23749 10241 23755
rect 10183 23724 10195 23749
rect 6825 23715 6883 23721
rect 6825 23681 6837 23715
rect 6871 23681 6883 23715
rect 6825 23675 6883 23681
rect 7561 23715 7619 23721
rect 7561 23681 7573 23715
rect 7607 23681 7619 23715
rect 7742 23712 7748 23724
rect 7703 23684 7748 23712
rect 7561 23675 7619 23681
rect 5353 23647 5411 23653
rect 5353 23644 5365 23647
rect 4816 23616 5365 23644
rect 4816 23520 4844 23616
rect 5353 23613 5365 23616
rect 5399 23613 5411 23647
rect 5353 23607 5411 23613
rect 5813 23647 5871 23653
rect 5813 23613 5825 23647
rect 5859 23644 5871 23647
rect 6840 23644 6868 23675
rect 7742 23672 7748 23684
rect 7800 23672 7806 23724
rect 8757 23715 8815 23721
rect 8757 23681 8769 23715
rect 8803 23712 8815 23715
rect 9217 23715 9275 23721
rect 9217 23712 9229 23715
rect 8803 23684 9229 23712
rect 8803 23681 8815 23684
rect 8757 23675 8815 23681
rect 9217 23681 9229 23684
rect 9263 23712 9275 23715
rect 9306 23712 9312 23724
rect 9263 23684 9312 23712
rect 9263 23681 9275 23684
rect 9217 23675 9275 23681
rect 9306 23672 9312 23684
rect 9364 23672 9370 23724
rect 9493 23715 9551 23721
rect 9493 23681 9505 23715
rect 9539 23712 9551 23715
rect 10134 23712 10140 23724
rect 9539 23684 10140 23712
rect 9539 23681 9551 23684
rect 9493 23675 9551 23681
rect 10134 23672 10140 23684
rect 10192 23715 10195 23724
rect 10229 23715 10241 23749
rect 10192 23712 10241 23715
rect 12434 23712 12440 23724
rect 10192 23684 12440 23712
rect 10192 23672 10198 23684
rect 12434 23672 12440 23684
rect 12492 23672 12498 23724
rect 12820 23721 12848 23808
rect 16758 23780 16764 23792
rect 13372 23752 16764 23780
rect 12621 23715 12679 23721
rect 12621 23712 12633 23715
rect 12544 23684 12633 23712
rect 12544 23656 12572 23684
rect 12621 23681 12633 23684
rect 12667 23681 12679 23715
rect 12621 23675 12679 23681
rect 12709 23715 12767 23721
rect 12709 23681 12721 23715
rect 12755 23681 12767 23715
rect 12709 23675 12767 23681
rect 12805 23715 12863 23721
rect 12805 23681 12817 23715
rect 12851 23681 12863 23715
rect 12805 23675 12863 23681
rect 7006 23644 7012 23656
rect 5859 23616 7012 23644
rect 5859 23613 5871 23616
rect 5813 23607 5871 23613
rect 7006 23604 7012 23616
rect 7064 23604 7070 23656
rect 7929 23647 7987 23653
rect 7929 23613 7941 23647
rect 7975 23644 7987 23647
rect 12526 23644 12532 23656
rect 7975 23616 12532 23644
rect 7975 23613 7987 23616
rect 7929 23607 7987 23613
rect 12526 23604 12532 23616
rect 12584 23604 12590 23656
rect 9214 23576 9220 23588
rect 9175 23548 9220 23576
rect 9214 23536 9220 23548
rect 9272 23536 9278 23588
rect 12728 23576 12756 23675
rect 12986 23576 12992 23588
rect 10060 23548 12756 23576
rect 12947 23548 12992 23576
rect 4798 23508 4804 23520
rect 4759 23480 4804 23508
rect 4798 23468 4804 23480
rect 4856 23468 4862 23520
rect 8018 23468 8024 23520
rect 8076 23508 8082 23520
rect 10060 23508 10088 23548
rect 12986 23536 12992 23548
rect 13044 23536 13050 23588
rect 8076 23480 10088 23508
rect 10137 23511 10195 23517
rect 8076 23468 8082 23480
rect 10137 23477 10149 23511
rect 10183 23508 10195 23511
rect 10594 23508 10600 23520
rect 10183 23480 10600 23508
rect 10183 23477 10195 23480
rect 10137 23471 10195 23477
rect 10594 23468 10600 23480
rect 10652 23468 10658 23520
rect 12526 23468 12532 23520
rect 12584 23508 12590 23520
rect 13372 23508 13400 23752
rect 16758 23740 16764 23752
rect 16816 23780 16822 23792
rect 16853 23783 16911 23789
rect 16853 23780 16865 23783
rect 16816 23752 16865 23780
rect 16816 23740 16822 23752
rect 16853 23749 16865 23752
rect 16899 23749 16911 23783
rect 16853 23743 16911 23749
rect 17862 23740 17868 23792
rect 17920 23780 17926 23792
rect 20640 23780 20668 23820
rect 20714 23808 20720 23860
rect 20772 23808 20778 23860
rect 21174 23808 21180 23860
rect 21232 23848 21238 23860
rect 21358 23848 21364 23860
rect 21232 23820 21364 23848
rect 21232 23808 21238 23820
rect 21358 23808 21364 23820
rect 21416 23808 21422 23860
rect 23014 23848 23020 23860
rect 22975 23820 23020 23848
rect 23014 23808 23020 23820
rect 23072 23808 23078 23860
rect 23216 23820 26832 23848
rect 17920 23752 20300 23780
rect 17920 23740 17926 23752
rect 20272 23734 20300 23752
rect 20548 23752 20668 23780
rect 20431 23737 20489 23743
rect 20431 23734 20443 23737
rect 13630 23712 13636 23724
rect 13591 23684 13636 23712
rect 13630 23672 13636 23684
rect 13688 23672 13694 23724
rect 14550 23672 14556 23724
rect 14608 23712 14614 23724
rect 14608 23684 16528 23712
rect 14608 23672 14614 23684
rect 13449 23647 13507 23653
rect 13449 23613 13461 23647
rect 13495 23644 13507 23647
rect 13538 23644 13544 23656
rect 13495 23616 13544 23644
rect 13495 23613 13507 23616
rect 13449 23607 13507 23613
rect 13538 23604 13544 23616
rect 13596 23644 13602 23656
rect 16500 23644 16528 23684
rect 16574 23672 16580 23724
rect 16632 23712 16638 23724
rect 16669 23715 16727 23721
rect 16669 23712 16681 23715
rect 16632 23684 16681 23712
rect 16632 23672 16638 23684
rect 16669 23681 16681 23684
rect 16715 23681 16727 23715
rect 16942 23712 16948 23724
rect 16903 23684 16948 23712
rect 16669 23675 16727 23681
rect 16942 23672 16948 23684
rect 17000 23672 17006 23724
rect 17034 23672 17040 23724
rect 17092 23712 17098 23724
rect 17957 23715 18015 23721
rect 17092 23684 17137 23712
rect 17092 23672 17098 23684
rect 17957 23681 17969 23715
rect 18003 23681 18015 23715
rect 17957 23675 18015 23681
rect 17770 23644 17776 23656
rect 13596 23616 15884 23644
rect 16500 23616 17776 23644
rect 13596 23604 13602 23616
rect 12584 23480 13400 23508
rect 12584 23468 12590 23480
rect 14090 23468 14096 23520
rect 14148 23508 14154 23520
rect 14277 23511 14335 23517
rect 14277 23508 14289 23511
rect 14148 23480 14289 23508
rect 14148 23468 14154 23480
rect 14277 23477 14289 23480
rect 14323 23477 14335 23511
rect 15856 23508 15884 23616
rect 17770 23604 17776 23616
rect 17828 23644 17834 23656
rect 17972 23644 18000 23675
rect 18414 23672 18420 23724
rect 18472 23712 18478 23724
rect 18877 23715 18935 23721
rect 18877 23712 18889 23715
rect 18472 23684 18889 23712
rect 18472 23672 18478 23684
rect 18877 23681 18889 23684
rect 18923 23681 18935 23715
rect 18877 23675 18935 23681
rect 18966 23672 18972 23724
rect 19024 23712 19030 23724
rect 19426 23712 19432 23724
rect 19024 23684 19432 23712
rect 19024 23672 19030 23684
rect 19426 23672 19432 23684
rect 19484 23712 19490 23724
rect 19613 23715 19671 23721
rect 19613 23712 19625 23715
rect 19484 23684 19625 23712
rect 19484 23672 19490 23684
rect 19613 23681 19625 23684
rect 19659 23681 19671 23715
rect 19613 23675 19671 23681
rect 19797 23715 19855 23721
rect 19797 23681 19809 23715
rect 19843 23712 19855 23715
rect 20162 23712 20168 23724
rect 19843 23684 20168 23712
rect 19843 23681 19855 23684
rect 19797 23675 19855 23681
rect 20162 23672 20168 23684
rect 20220 23672 20226 23724
rect 20272 23706 20443 23734
rect 20431 23703 20443 23706
rect 20477 23703 20489 23737
rect 20548 23721 20576 23752
rect 20431 23697 20489 23703
rect 20533 23715 20591 23721
rect 20533 23681 20545 23715
rect 20579 23681 20591 23715
rect 20533 23675 20591 23681
rect 20644 23715 20702 23721
rect 20644 23681 20656 23715
rect 20690 23712 20702 23715
rect 20744 23712 20772 23808
rect 20898 23740 20904 23792
rect 20956 23780 20962 23792
rect 23216 23780 23244 23820
rect 20956 23752 23244 23780
rect 23477 23783 23535 23789
rect 20956 23740 20962 23752
rect 23477 23749 23489 23783
rect 23523 23780 23535 23783
rect 23566 23780 23572 23792
rect 23523 23752 23572 23780
rect 23523 23749 23535 23752
rect 23477 23743 23535 23749
rect 20690 23684 20772 23712
rect 20690 23681 20702 23684
rect 20732 23682 20772 23684
rect 20809 23715 20867 23721
rect 20644 23675 20702 23681
rect 20809 23681 20821 23715
rect 20855 23712 20867 23715
rect 20990 23712 20996 23724
rect 20855 23684 20996 23712
rect 20855 23681 20867 23684
rect 20809 23675 20867 23681
rect 20990 23672 20996 23684
rect 21048 23672 21054 23724
rect 17828 23616 18000 23644
rect 17828 23604 17834 23616
rect 18322 23604 18328 23656
rect 18380 23644 18386 23656
rect 19978 23644 19984 23656
rect 18380 23616 19984 23644
rect 18380 23604 18386 23616
rect 19978 23604 19984 23616
rect 20036 23644 20042 23656
rect 23492 23644 23520 23743
rect 23566 23740 23572 23752
rect 23624 23740 23630 23792
rect 24946 23780 24952 23792
rect 24907 23752 24952 23780
rect 24946 23740 24952 23752
rect 25004 23740 25010 23792
rect 25777 23783 25835 23789
rect 25777 23749 25789 23783
rect 25823 23749 25835 23783
rect 25958 23780 25964 23792
rect 25919 23752 25964 23780
rect 25777 23743 25835 23749
rect 23750 23672 23756 23724
rect 23808 23712 23814 23724
rect 23845 23715 23903 23721
rect 23845 23712 23857 23715
rect 23808 23684 23857 23712
rect 23808 23672 23814 23684
rect 23845 23681 23857 23684
rect 23891 23681 23903 23715
rect 23845 23675 23903 23681
rect 23934 23672 23940 23724
rect 23992 23712 23998 23724
rect 24588 23715 24646 23721
rect 24588 23713 24600 23715
rect 24504 23712 24600 23713
rect 23992 23684 24037 23712
rect 24136 23685 24600 23712
rect 24136 23684 24532 23685
rect 23992 23672 23998 23684
rect 20036 23616 23520 23644
rect 23569 23647 23627 23653
rect 20036 23604 20042 23616
rect 23569 23613 23581 23647
rect 23615 23644 23627 23647
rect 23658 23644 23664 23656
rect 23615 23616 23664 23644
rect 23615 23613 23627 23616
rect 23569 23607 23627 23613
rect 18046 23536 18052 23588
rect 18104 23576 18110 23588
rect 18414 23576 18420 23588
rect 18104 23548 18420 23576
rect 18104 23536 18110 23548
rect 18414 23536 18420 23548
rect 18472 23536 18478 23588
rect 20530 23536 20536 23588
rect 20588 23576 20594 23588
rect 20993 23579 21051 23585
rect 20588 23548 20668 23576
rect 20588 23536 20594 23548
rect 18966 23508 18972 23520
rect 15856 23480 18972 23508
rect 14277 23471 14335 23477
rect 18966 23468 18972 23480
rect 19024 23468 19030 23520
rect 19061 23511 19119 23517
rect 19061 23477 19073 23511
rect 19107 23508 19119 23511
rect 19334 23508 19340 23520
rect 19107 23480 19340 23508
rect 19107 23477 19119 23480
rect 19061 23471 19119 23477
rect 19334 23468 19340 23480
rect 19392 23468 19398 23520
rect 20640 23508 20668 23548
rect 20993 23545 21005 23579
rect 21039 23576 21051 23579
rect 21634 23576 21640 23588
rect 21039 23548 21640 23576
rect 21039 23545 21051 23548
rect 20993 23539 21051 23545
rect 21634 23536 21640 23548
rect 21692 23536 21698 23588
rect 23584 23576 23612 23607
rect 23658 23604 23664 23616
rect 23716 23604 23722 23656
rect 24136 23585 24164 23684
rect 24588 23681 24600 23685
rect 24634 23681 24646 23715
rect 24588 23675 24646 23681
rect 24674 23715 24732 23721
rect 24674 23681 24686 23715
rect 24720 23681 24732 23715
rect 24674 23675 24732 23681
rect 24857 23715 24915 23721
rect 24857 23681 24869 23715
rect 24903 23681 24915 23715
rect 24857 23675 24915 23681
rect 22066 23548 23612 23576
rect 24121 23579 24179 23585
rect 22066 23508 22094 23548
rect 24121 23545 24133 23579
rect 24167 23545 24179 23579
rect 24121 23539 24179 23545
rect 24302 23536 24308 23588
rect 24360 23576 24366 23588
rect 24688 23576 24716 23675
rect 24762 23604 24768 23656
rect 24820 23644 24826 23656
rect 24872 23644 24900 23675
rect 25038 23672 25044 23724
rect 25096 23721 25102 23724
rect 25096 23712 25104 23721
rect 25096 23684 25141 23712
rect 25096 23675 25104 23684
rect 25096 23672 25102 23675
rect 24820 23616 24900 23644
rect 24820 23604 24826 23616
rect 25792 23576 25820 23743
rect 25958 23740 25964 23752
rect 26016 23740 26022 23792
rect 26804 23780 26832 23820
rect 31294 23808 31300 23860
rect 31352 23848 31358 23860
rect 46937 23851 46995 23857
rect 31352 23820 44128 23848
rect 31352 23808 31358 23820
rect 34793 23783 34851 23789
rect 26804 23752 31754 23780
rect 30929 23715 30987 23721
rect 30929 23712 30941 23715
rect 30208 23684 30941 23712
rect 30208 23585 30236 23684
rect 30929 23681 30941 23684
rect 30975 23681 30987 23715
rect 30929 23675 30987 23681
rect 30745 23647 30803 23653
rect 30745 23644 30757 23647
rect 30300 23616 30757 23644
rect 30193 23579 30251 23585
rect 30193 23576 30205 23579
rect 24360 23548 24716 23576
rect 24780 23548 25820 23576
rect 28828 23548 30205 23576
rect 24360 23536 24366 23548
rect 20640 23480 22094 23508
rect 23566 23468 23572 23520
rect 23624 23508 23630 23520
rect 24780 23508 24808 23548
rect 28828 23520 28856 23548
rect 30193 23545 30205 23548
rect 30239 23545 30251 23579
rect 30193 23539 30251 23545
rect 23624 23480 24808 23508
rect 25225 23511 25283 23517
rect 23624 23468 23630 23480
rect 25225 23477 25237 23511
rect 25271 23508 25283 23511
rect 25406 23508 25412 23520
rect 25271 23480 25412 23508
rect 25271 23477 25283 23480
rect 25225 23471 25283 23477
rect 25406 23468 25412 23480
rect 25464 23468 25470 23520
rect 27706 23468 27712 23520
rect 27764 23508 27770 23520
rect 28353 23511 28411 23517
rect 28353 23508 28365 23511
rect 27764 23480 28365 23508
rect 27764 23468 27770 23480
rect 28353 23477 28365 23480
rect 28399 23508 28411 23511
rect 28810 23508 28816 23520
rect 28399 23480 28816 23508
rect 28399 23477 28411 23480
rect 28353 23471 28411 23477
rect 28810 23468 28816 23480
rect 28868 23468 28874 23520
rect 29638 23508 29644 23520
rect 29599 23480 29644 23508
rect 29638 23468 29644 23480
rect 29696 23508 29702 23520
rect 30300 23508 30328 23616
rect 30745 23613 30757 23616
rect 30791 23613 30803 23647
rect 30745 23607 30803 23613
rect 31110 23604 31116 23656
rect 31168 23644 31174 23656
rect 31297 23647 31355 23653
rect 31297 23644 31309 23647
rect 31168 23616 31309 23644
rect 31168 23604 31174 23616
rect 31297 23613 31309 23616
rect 31343 23613 31355 23647
rect 31726 23644 31754 23752
rect 34793 23749 34805 23783
rect 34839 23780 34851 23783
rect 35434 23780 35440 23792
rect 34839 23752 35440 23780
rect 34839 23749 34851 23752
rect 34793 23743 34851 23749
rect 35434 23740 35440 23752
rect 35492 23740 35498 23792
rect 37921 23783 37979 23789
rect 37292 23752 37872 23780
rect 37292 23724 37320 23752
rect 34609 23715 34667 23721
rect 34609 23681 34621 23715
rect 34655 23712 34667 23715
rect 34698 23712 34704 23724
rect 34655 23684 34704 23712
rect 34655 23681 34667 23684
rect 34609 23675 34667 23681
rect 34698 23672 34704 23684
rect 34756 23672 34762 23724
rect 34882 23672 34888 23724
rect 34940 23712 34946 23724
rect 37274 23712 37280 23724
rect 34940 23684 34985 23712
rect 37187 23684 37280 23712
rect 34940 23672 34946 23684
rect 37274 23672 37280 23684
rect 37332 23672 37338 23724
rect 37458 23712 37464 23724
rect 37419 23684 37464 23712
rect 37458 23672 37464 23684
rect 37516 23672 37522 23724
rect 37734 23712 37740 23724
rect 37695 23684 37740 23712
rect 37734 23672 37740 23684
rect 37792 23672 37798 23724
rect 37844 23712 37872 23752
rect 37921 23749 37933 23783
rect 37967 23780 37979 23783
rect 41046 23780 41052 23792
rect 37967 23752 41052 23780
rect 37967 23749 37979 23752
rect 37921 23743 37979 23749
rect 41046 23740 41052 23752
rect 41104 23740 41110 23792
rect 43530 23740 43536 23792
rect 43588 23780 43594 23792
rect 43990 23789 43996 23792
rect 43717 23783 43775 23789
rect 43717 23780 43729 23783
rect 43588 23752 43729 23780
rect 43588 23740 43594 23752
rect 43717 23749 43729 23752
rect 43763 23749 43775 23783
rect 43717 23743 43775 23749
rect 43933 23783 43996 23789
rect 43933 23749 43945 23783
rect 43979 23749 43996 23783
rect 43933 23743 43996 23749
rect 43990 23740 43996 23743
rect 44048 23740 44054 23792
rect 44100 23780 44128 23820
rect 46937 23817 46949 23851
rect 46983 23848 46995 23851
rect 47302 23848 47308 23860
rect 46983 23820 47308 23848
rect 46983 23817 46995 23820
rect 46937 23811 46995 23817
rect 47302 23808 47308 23820
rect 47360 23848 47366 23860
rect 47854 23848 47860 23860
rect 47360 23820 47860 23848
rect 47360 23808 47366 23820
rect 47854 23808 47860 23820
rect 47912 23808 47918 23860
rect 48038 23848 48044 23860
rect 47999 23820 48044 23848
rect 48038 23808 48044 23820
rect 48096 23808 48102 23860
rect 53190 23848 53196 23860
rect 53151 23820 53196 23848
rect 53190 23808 53196 23820
rect 53248 23808 53254 23860
rect 55766 23808 55772 23860
rect 55824 23848 55830 23860
rect 56045 23851 56103 23857
rect 56045 23848 56057 23851
rect 55824 23820 56057 23848
rect 55824 23808 55830 23820
rect 56045 23817 56057 23820
rect 56091 23817 56103 23851
rect 56045 23811 56103 23817
rect 46293 23783 46351 23789
rect 46293 23780 46305 23783
rect 44100 23752 46305 23780
rect 46293 23749 46305 23752
rect 46339 23780 46351 23783
rect 49510 23780 49516 23792
rect 46339 23752 49516 23780
rect 46339 23749 46351 23752
rect 46293 23743 46351 23749
rect 40126 23712 40132 23724
rect 37844 23684 40132 23712
rect 40126 23672 40132 23684
rect 40184 23672 40190 23724
rect 47044 23721 47072 23752
rect 49510 23740 49516 23752
rect 49568 23780 49574 23792
rect 49568 23752 51212 23780
rect 49568 23740 49574 23752
rect 46845 23715 46903 23721
rect 46845 23712 46857 23715
rect 41386 23684 46857 23712
rect 39393 23647 39451 23653
rect 39393 23644 39405 23647
rect 31726 23616 39405 23644
rect 31297 23607 31355 23613
rect 39393 23613 39405 23616
rect 39439 23644 39451 23647
rect 40037 23647 40095 23653
rect 40037 23644 40049 23647
rect 39439 23616 40049 23644
rect 39439 23613 39451 23616
rect 39393 23607 39451 23613
rect 40037 23613 40049 23616
rect 40083 23613 40095 23647
rect 40037 23607 40095 23613
rect 31205 23579 31263 23585
rect 31205 23545 31217 23579
rect 31251 23576 31263 23579
rect 41386 23576 41414 23684
rect 46845 23681 46857 23684
rect 46891 23681 46903 23715
rect 46845 23675 46903 23681
rect 47029 23715 47087 23721
rect 47029 23681 47041 23715
rect 47075 23681 47087 23715
rect 47029 23675 47087 23681
rect 50246 23672 50252 23724
rect 50304 23712 50310 23724
rect 50341 23715 50399 23721
rect 50341 23712 50353 23715
rect 50304 23684 50353 23712
rect 50304 23672 50310 23684
rect 50341 23681 50353 23684
rect 50387 23681 50399 23715
rect 50341 23675 50399 23681
rect 50525 23715 50583 23721
rect 50525 23681 50537 23715
rect 50571 23712 50583 23715
rect 50614 23712 50620 23724
rect 50571 23684 50620 23712
rect 50571 23681 50583 23684
rect 50525 23675 50583 23681
rect 50614 23672 50620 23684
rect 50672 23672 50678 23724
rect 50985 23715 51043 23721
rect 50985 23681 50997 23715
rect 51031 23712 51043 23715
rect 51074 23712 51080 23724
rect 51031 23684 51080 23712
rect 51031 23681 51043 23684
rect 50985 23675 51043 23681
rect 51074 23672 51080 23684
rect 51132 23672 51138 23724
rect 51184 23721 51212 23752
rect 55306 23740 55312 23792
rect 55364 23780 55370 23792
rect 55364 23752 56180 23780
rect 55364 23740 55370 23752
rect 51169 23715 51227 23721
rect 51169 23681 51181 23715
rect 51215 23712 51227 23715
rect 51629 23715 51687 23721
rect 51629 23712 51641 23715
rect 51215 23684 51641 23712
rect 51215 23681 51227 23684
rect 51169 23675 51227 23681
rect 51629 23681 51641 23684
rect 51675 23681 51687 23715
rect 51629 23675 51687 23681
rect 52270 23672 52276 23724
rect 52328 23712 52334 23724
rect 53009 23715 53067 23721
rect 53009 23712 53021 23715
rect 52328 23684 53021 23712
rect 52328 23672 52334 23684
rect 53009 23681 53021 23684
rect 53055 23681 53067 23715
rect 53009 23675 53067 23681
rect 55674 23672 55680 23724
rect 55732 23712 55738 23724
rect 56152 23721 56180 23752
rect 55953 23715 56011 23721
rect 55953 23712 55965 23715
rect 55732 23684 55965 23712
rect 55732 23672 55738 23684
rect 55953 23681 55965 23684
rect 55999 23681 56011 23715
rect 55953 23675 56011 23681
rect 56137 23715 56195 23721
rect 56137 23681 56149 23715
rect 56183 23681 56195 23715
rect 56137 23675 56195 23681
rect 47578 23644 47584 23656
rect 47539 23616 47584 23644
rect 47578 23604 47584 23616
rect 47636 23604 47642 23656
rect 52730 23644 52736 23656
rect 52691 23616 52736 23644
rect 52730 23604 52736 23616
rect 52788 23604 52794 23656
rect 31251 23548 41414 23576
rect 44085 23579 44143 23585
rect 31251 23545 31263 23548
rect 31205 23539 31263 23545
rect 44085 23545 44097 23579
rect 44131 23576 44143 23579
rect 45370 23576 45376 23588
rect 44131 23548 45376 23576
rect 44131 23545 44143 23548
rect 44085 23539 44143 23545
rect 45370 23536 45376 23548
rect 45428 23536 45434 23588
rect 47394 23536 47400 23588
rect 47452 23576 47458 23588
rect 47857 23579 47915 23585
rect 47857 23576 47869 23579
rect 47452 23548 47869 23576
rect 47452 23536 47458 23548
rect 47857 23545 47869 23548
rect 47903 23545 47915 23579
rect 47857 23539 47915 23545
rect 50433 23579 50491 23585
rect 50433 23545 50445 23579
rect 50479 23576 50491 23579
rect 52270 23576 52276 23588
rect 50479 23548 52276 23576
rect 50479 23545 50491 23548
rect 50433 23539 50491 23545
rect 52270 23536 52276 23548
rect 52328 23536 52334 23588
rect 29696 23480 30328 23508
rect 34609 23511 34667 23517
rect 29696 23468 29702 23480
rect 34609 23477 34621 23511
rect 34655 23508 34667 23511
rect 36538 23508 36544 23520
rect 34655 23480 36544 23508
rect 34655 23477 34667 23480
rect 34609 23471 34667 23477
rect 36538 23468 36544 23480
rect 36596 23468 36602 23520
rect 36722 23508 36728 23520
rect 36683 23480 36728 23508
rect 36722 23468 36728 23480
rect 36780 23508 36786 23520
rect 37458 23508 37464 23520
rect 36780 23480 37464 23508
rect 36780 23468 36786 23480
rect 37458 23468 37464 23480
rect 37516 23468 37522 23520
rect 40405 23511 40463 23517
rect 40405 23477 40417 23511
rect 40451 23508 40463 23511
rect 41598 23508 41604 23520
rect 40451 23480 41604 23508
rect 40451 23477 40463 23480
rect 40405 23471 40463 23477
rect 41598 23468 41604 23480
rect 41656 23468 41662 23520
rect 43898 23508 43904 23520
rect 43859 23480 43904 23508
rect 43898 23468 43904 23480
rect 43956 23468 43962 23520
rect 51077 23511 51135 23517
rect 51077 23477 51089 23511
rect 51123 23508 51135 23511
rect 52086 23508 52092 23520
rect 51123 23480 52092 23508
rect 51123 23477 51135 23480
rect 51077 23471 51135 23477
rect 52086 23468 52092 23480
rect 52144 23468 52150 23520
rect 52822 23508 52828 23520
rect 52783 23480 52828 23508
rect 52822 23468 52828 23480
rect 52880 23468 52886 23520
rect 57882 23468 57888 23520
rect 57940 23508 57946 23520
rect 58069 23511 58127 23517
rect 58069 23508 58081 23511
rect 57940 23480 58081 23508
rect 57940 23468 57946 23480
rect 58069 23477 58081 23480
rect 58115 23477 58127 23511
rect 58069 23471 58127 23477
rect 1104 23418 58880 23440
rect 1104 23366 4214 23418
rect 4266 23366 4278 23418
rect 4330 23366 4342 23418
rect 4394 23366 4406 23418
rect 4458 23366 4470 23418
rect 4522 23366 34934 23418
rect 34986 23366 34998 23418
rect 35050 23366 35062 23418
rect 35114 23366 35126 23418
rect 35178 23366 35190 23418
rect 35242 23366 58880 23418
rect 1104 23344 58880 23366
rect 4341 23307 4399 23313
rect 4341 23273 4353 23307
rect 4387 23304 4399 23307
rect 6822 23304 6828 23316
rect 4387 23276 6828 23304
rect 4387 23273 4399 23276
rect 4341 23267 4399 23273
rect 6822 23264 6828 23276
rect 6880 23264 6886 23316
rect 7282 23264 7288 23316
rect 7340 23304 7346 23316
rect 7340 23276 8248 23304
rect 7340 23264 7346 23276
rect 6457 23239 6515 23245
rect 6457 23205 6469 23239
rect 6503 23236 6515 23239
rect 7377 23239 7435 23245
rect 7377 23236 7389 23239
rect 6503 23208 7389 23236
rect 6503 23205 6515 23208
rect 6457 23199 6515 23205
rect 7377 23205 7389 23208
rect 7423 23236 7435 23239
rect 7742 23236 7748 23248
rect 7423 23208 7748 23236
rect 7423 23205 7435 23208
rect 7377 23199 7435 23205
rect 7742 23196 7748 23208
rect 7800 23196 7806 23248
rect 8220 23245 8248 23276
rect 9306 23264 9312 23316
rect 9364 23304 9370 23316
rect 9490 23304 9496 23316
rect 9364 23276 9496 23304
rect 9364 23264 9370 23276
rect 9490 23264 9496 23276
rect 9548 23304 9554 23316
rect 12989 23307 13047 23313
rect 12989 23304 13001 23307
rect 9548 23276 13001 23304
rect 9548 23264 9554 23276
rect 12989 23273 13001 23276
rect 13035 23304 13047 23307
rect 14277 23307 14335 23313
rect 14277 23304 14289 23307
rect 13035 23276 14289 23304
rect 13035 23273 13047 23276
rect 12989 23267 13047 23273
rect 14277 23273 14289 23276
rect 14323 23304 14335 23307
rect 15470 23304 15476 23316
rect 14323 23276 15476 23304
rect 14323 23273 14335 23276
rect 14277 23267 14335 23273
rect 15470 23264 15476 23276
rect 15528 23264 15534 23316
rect 20806 23264 20812 23316
rect 20864 23304 20870 23316
rect 23750 23304 23756 23316
rect 20864 23276 23756 23304
rect 20864 23264 20870 23276
rect 23750 23264 23756 23276
rect 23808 23264 23814 23316
rect 23845 23307 23903 23313
rect 23845 23273 23857 23307
rect 23891 23304 23903 23307
rect 24486 23304 24492 23316
rect 23891 23276 24492 23304
rect 23891 23273 23903 23276
rect 23845 23267 23903 23273
rect 24486 23264 24492 23276
rect 24544 23264 24550 23316
rect 30377 23307 30435 23313
rect 30377 23273 30389 23307
rect 30423 23304 30435 23307
rect 31110 23304 31116 23316
rect 30423 23276 31116 23304
rect 30423 23273 30435 23276
rect 30377 23267 30435 23273
rect 31110 23264 31116 23276
rect 31168 23264 31174 23316
rect 34977 23307 35035 23313
rect 34977 23273 34989 23307
rect 35023 23304 35035 23307
rect 35434 23304 35440 23316
rect 35023 23276 35440 23304
rect 35023 23273 35035 23276
rect 34977 23267 35035 23273
rect 35434 23264 35440 23276
rect 35492 23264 35498 23316
rect 54757 23307 54815 23313
rect 54757 23273 54769 23307
rect 54803 23304 54815 23307
rect 55306 23304 55312 23316
rect 54803 23276 55312 23304
rect 54803 23273 54815 23276
rect 54757 23267 54815 23273
rect 55306 23264 55312 23276
rect 55364 23264 55370 23316
rect 55490 23304 55496 23316
rect 55451 23276 55496 23304
rect 55490 23264 55496 23276
rect 55548 23264 55554 23316
rect 8205 23239 8263 23245
rect 8205 23205 8217 23239
rect 8251 23236 8263 23239
rect 12802 23236 12808 23248
rect 8251 23208 12808 23236
rect 8251 23205 8263 23208
rect 8205 23199 8263 23205
rect 12802 23196 12808 23208
rect 12860 23196 12866 23248
rect 13814 23196 13820 23248
rect 13872 23236 13878 23248
rect 13872 23208 15148 23236
rect 13872 23196 13878 23208
rect 6178 23168 6184 23180
rect 6139 23140 6184 23168
rect 6178 23128 6184 23140
rect 6236 23128 6242 23180
rect 7006 23168 7012 23180
rect 6967 23140 7012 23168
rect 7006 23128 7012 23140
rect 7064 23128 7070 23180
rect 7469 23171 7527 23177
rect 7469 23137 7481 23171
rect 7515 23168 7527 23171
rect 12820 23168 12848 23196
rect 15010 23168 15016 23180
rect 7515 23140 12434 23168
rect 12820 23140 15016 23168
rect 7515 23137 7527 23140
rect 7469 23131 7527 23137
rect 1854 23100 1860 23112
rect 1815 23072 1860 23100
rect 1854 23060 1860 23072
rect 1912 23060 1918 23112
rect 4249 23103 4307 23109
rect 4249 23069 4261 23103
rect 4295 23100 4307 23103
rect 4614 23100 4620 23112
rect 4295 23072 4620 23100
rect 4295 23069 4307 23072
rect 4249 23063 4307 23069
rect 4614 23060 4620 23072
rect 4672 23060 4678 23112
rect 6089 23103 6147 23109
rect 6089 23069 6101 23103
rect 6135 23069 6147 23103
rect 8018 23100 8024 23112
rect 7979 23072 8024 23100
rect 6089 23063 6147 23069
rect 2038 23032 2044 23044
rect 1999 23004 2044 23032
rect 2038 22992 2044 23004
rect 2096 22992 2102 23044
rect 4798 22992 4804 23044
rect 4856 23032 4862 23044
rect 5353 23035 5411 23041
rect 5353 23032 5365 23035
rect 4856 23004 5365 23032
rect 4856 22992 4862 23004
rect 5353 23001 5365 23004
rect 5399 23032 5411 23035
rect 6104 23032 6132 23063
rect 8018 23060 8024 23072
rect 8076 23060 8082 23112
rect 9858 23100 9864 23112
rect 9819 23072 9864 23100
rect 9858 23060 9864 23072
rect 9916 23060 9922 23112
rect 10134 23100 10140 23112
rect 10095 23072 10140 23100
rect 10134 23060 10140 23072
rect 10192 23060 10198 23112
rect 12406 23100 12434 23140
rect 12618 23100 12624 23112
rect 12406 23072 12624 23100
rect 12618 23060 12624 23072
rect 12676 23100 12682 23112
rect 13630 23100 13636 23112
rect 12676 23072 13636 23100
rect 12676 23060 12682 23072
rect 13630 23060 13636 23072
rect 13688 23060 13694 23112
rect 5399 23004 6132 23032
rect 14093 23035 14151 23041
rect 5399 23001 5411 23004
rect 5353 22995 5411 23001
rect 14093 23001 14105 23035
rect 14139 23001 14151 23035
rect 14200 23032 14228 23140
rect 15010 23128 15016 23140
rect 15068 23128 15074 23180
rect 15120 23100 15148 23208
rect 20254 23196 20260 23248
rect 20312 23236 20318 23248
rect 21634 23236 21640 23248
rect 20312 23208 21640 23236
rect 20312 23196 20318 23208
rect 21634 23196 21640 23208
rect 21692 23196 21698 23248
rect 23014 23196 23020 23248
rect 23072 23236 23078 23248
rect 23201 23239 23259 23245
rect 23201 23236 23213 23239
rect 23072 23208 23213 23236
rect 23072 23196 23078 23208
rect 23201 23205 23213 23208
rect 23247 23236 23259 23239
rect 24762 23236 24768 23248
rect 23247 23208 24768 23236
rect 23247 23205 23259 23208
rect 23201 23199 23259 23205
rect 24762 23196 24768 23208
rect 24820 23196 24826 23248
rect 35161 23239 35219 23245
rect 35161 23205 35173 23239
rect 35207 23236 35219 23239
rect 37734 23236 37740 23248
rect 35207 23208 37740 23236
rect 35207 23205 35219 23208
rect 35161 23199 35219 23205
rect 37734 23196 37740 23208
rect 37792 23196 37798 23248
rect 52730 23196 52736 23248
rect 52788 23236 52794 23248
rect 53469 23239 53527 23245
rect 53469 23236 53481 23239
rect 52788 23208 53481 23236
rect 52788 23196 52794 23208
rect 53469 23205 53481 23208
rect 53515 23205 53527 23239
rect 53469 23199 53527 23205
rect 16482 23128 16488 23180
rect 16540 23168 16546 23180
rect 16577 23171 16635 23177
rect 16577 23168 16589 23171
rect 16540 23140 16589 23168
rect 16540 23128 16546 23140
rect 16577 23137 16589 23140
rect 16623 23168 16635 23171
rect 18322 23168 18328 23180
rect 16623 23140 18328 23168
rect 16623 23137 16635 23140
rect 16577 23131 16635 23137
rect 15028 23072 15148 23100
rect 15028 23041 15056 23072
rect 15378 23060 15384 23112
rect 15436 23100 15442 23112
rect 16390 23100 16396 23112
rect 15436 23072 16396 23100
rect 15436 23060 15442 23072
rect 16390 23060 16396 23072
rect 16448 23100 16454 23112
rect 17512 23109 17540 23140
rect 18322 23128 18328 23140
rect 18380 23128 18386 23180
rect 19978 23128 19984 23180
rect 20036 23168 20042 23180
rect 26697 23171 26755 23177
rect 26697 23168 26709 23171
rect 20036 23140 26709 23168
rect 20036 23128 20042 23140
rect 26697 23137 26709 23140
rect 26743 23137 26755 23171
rect 29549 23171 29607 23177
rect 29549 23168 29561 23171
rect 26697 23131 26755 23137
rect 28828 23140 29561 23168
rect 28828 23112 28856 23140
rect 29549 23137 29561 23140
rect 29595 23137 29607 23171
rect 32401 23171 32459 23177
rect 29549 23131 29607 23137
rect 30852 23140 31616 23168
rect 17313 23103 17371 23109
rect 17313 23100 17325 23103
rect 16448 23072 17325 23100
rect 16448 23060 16454 23072
rect 17313 23069 17325 23072
rect 17359 23069 17371 23103
rect 17313 23063 17371 23069
rect 17497 23103 17555 23109
rect 17497 23069 17509 23103
rect 17543 23069 17555 23103
rect 17497 23063 17555 23069
rect 17678 23060 17684 23112
rect 17736 23100 17742 23112
rect 20070 23100 20076 23112
rect 17736 23072 17829 23100
rect 19306 23072 20076 23100
rect 17736 23060 17742 23072
rect 14293 23035 14351 23041
rect 14293 23032 14305 23035
rect 14200 23004 14305 23032
rect 14093 22995 14151 23001
rect 14293 23001 14305 23004
rect 14339 23001 14351 23035
rect 14293 22995 14351 23001
rect 15013 23035 15071 23041
rect 15013 23001 15025 23035
rect 15059 23001 15071 23035
rect 15013 22995 15071 23001
rect 15197 23035 15255 23041
rect 15197 23001 15209 23035
rect 15243 23032 15255 23035
rect 16114 23032 16120 23044
rect 15243 23004 16120 23032
rect 15243 23001 15255 23004
rect 15197 22995 15255 23001
rect 11514 22924 11520 22976
rect 11572 22964 11578 22976
rect 13449 22967 13507 22973
rect 13449 22964 13461 22967
rect 11572 22936 13461 22964
rect 11572 22924 11578 22936
rect 13449 22933 13461 22936
rect 13495 22964 13507 22967
rect 13722 22964 13728 22976
rect 13495 22936 13728 22964
rect 13495 22933 13507 22936
rect 13449 22927 13507 22933
rect 13722 22924 13728 22936
rect 13780 22964 13786 22976
rect 14108 22964 14136 22995
rect 16114 22992 16120 23004
rect 16172 22992 16178 23044
rect 16758 23032 16764 23044
rect 16719 23004 16764 23032
rect 16758 22992 16764 23004
rect 16816 22992 16822 23044
rect 17586 23032 17592 23044
rect 17547 23004 17592 23032
rect 17586 22992 17592 23004
rect 17644 22992 17650 23044
rect 17696 23032 17724 23060
rect 19306 23032 19334 23072
rect 20070 23060 20076 23072
rect 20128 23060 20134 23112
rect 20990 23060 20996 23112
rect 21048 23100 21054 23112
rect 23017 23103 23075 23109
rect 23017 23100 23029 23103
rect 21048 23072 23029 23100
rect 21048 23060 21054 23072
rect 23017 23069 23029 23072
rect 23063 23069 23075 23103
rect 23017 23063 23075 23069
rect 23474 23060 23480 23112
rect 23532 23100 23538 23112
rect 23661 23103 23719 23109
rect 23661 23100 23673 23103
rect 23532 23072 23673 23100
rect 23532 23060 23538 23072
rect 23661 23069 23673 23072
rect 23707 23069 23719 23103
rect 23661 23063 23719 23069
rect 23750 23060 23756 23112
rect 23808 23100 23814 23112
rect 23845 23103 23903 23109
rect 23845 23100 23857 23103
rect 23808 23072 23857 23100
rect 23808 23060 23814 23072
rect 23845 23069 23857 23072
rect 23891 23069 23903 23103
rect 24854 23100 24860 23112
rect 24815 23072 24860 23100
rect 23845 23063 23903 23069
rect 24854 23060 24860 23072
rect 24912 23060 24918 23112
rect 26418 23060 26424 23112
rect 26476 23100 26482 23112
rect 26786 23100 26792 23112
rect 26476 23072 26792 23100
rect 26476 23060 26482 23072
rect 26786 23060 26792 23072
rect 26844 23060 26850 23112
rect 27617 23103 27675 23109
rect 27617 23069 27629 23103
rect 27663 23100 27675 23103
rect 27798 23100 27804 23112
rect 27663 23072 27804 23100
rect 27663 23069 27675 23072
rect 27617 23063 27675 23069
rect 27798 23060 27804 23072
rect 27856 23060 27862 23112
rect 28810 23100 28816 23112
rect 28771 23072 28816 23100
rect 28810 23060 28816 23072
rect 28868 23060 28874 23112
rect 28997 23103 29055 23109
rect 28997 23069 29009 23103
rect 29043 23100 29055 23103
rect 29733 23103 29791 23109
rect 29733 23100 29745 23103
rect 29043 23072 29745 23100
rect 29043 23069 29055 23072
rect 28997 23063 29055 23069
rect 29733 23069 29745 23072
rect 29779 23069 29791 23103
rect 29733 23063 29791 23069
rect 29917 23103 29975 23109
rect 29917 23069 29929 23103
rect 29963 23100 29975 23103
rect 30374 23100 30380 23112
rect 29963 23072 30380 23100
rect 29963 23069 29975 23072
rect 29917 23063 29975 23069
rect 17696 23004 19334 23032
rect 20162 22992 20168 23044
rect 20220 23032 20226 23044
rect 20441 23035 20499 23041
rect 20441 23032 20453 23035
rect 20220 23004 20453 23032
rect 20220 22992 20226 23004
rect 20441 23001 20453 23004
rect 20487 23032 20499 23035
rect 21450 23032 21456 23044
rect 20487 23004 21456 23032
rect 20487 23001 20499 23004
rect 20441 22995 20499 23001
rect 21450 22992 21456 23004
rect 21508 22992 21514 23044
rect 29012 23032 29040 23063
rect 30374 23060 30380 23072
rect 30432 23100 30438 23112
rect 30852 23109 30880 23140
rect 31588 23112 31616 23140
rect 32401 23137 32413 23171
rect 32447 23168 32459 23171
rect 43990 23168 43996 23180
rect 32447 23140 43996 23168
rect 32447 23137 32459 23140
rect 32401 23131 32459 23137
rect 43990 23128 43996 23140
rect 44048 23128 44054 23180
rect 44177 23171 44235 23177
rect 44177 23137 44189 23171
rect 44223 23168 44235 23171
rect 46477 23171 46535 23177
rect 44223 23140 46336 23168
rect 44223 23137 44235 23140
rect 44177 23131 44235 23137
rect 46308 23112 46336 23140
rect 46477 23137 46489 23171
rect 46523 23168 46535 23171
rect 46523 23140 47440 23168
rect 46523 23137 46535 23140
rect 46477 23131 46535 23137
rect 47412 23112 47440 23140
rect 51074 23128 51080 23180
rect 51132 23168 51138 23180
rect 51169 23171 51227 23177
rect 51169 23168 51181 23171
rect 51132 23140 51181 23168
rect 51132 23128 51138 23140
rect 51169 23137 51181 23140
rect 51215 23137 51227 23171
rect 52086 23168 52092 23180
rect 52047 23140 52092 23168
rect 51169 23131 51227 23137
rect 52086 23128 52092 23140
rect 52144 23128 52150 23180
rect 53282 23128 53288 23180
rect 53340 23128 53346 23180
rect 30561 23103 30619 23109
rect 30561 23100 30573 23103
rect 30432 23072 30573 23100
rect 30432 23060 30438 23072
rect 30561 23069 30573 23072
rect 30607 23069 30619 23103
rect 30561 23063 30619 23069
rect 30837 23103 30895 23109
rect 30837 23069 30849 23103
rect 30883 23069 30895 23103
rect 30837 23063 30895 23069
rect 31389 23103 31447 23109
rect 31389 23069 31401 23103
rect 31435 23069 31447 23103
rect 31389 23063 31447 23069
rect 27172 23004 29040 23032
rect 14458 22964 14464 22976
rect 13780 22936 14136 22964
rect 14419 22936 14464 22964
rect 13780 22924 13786 22936
rect 14458 22924 14464 22936
rect 14516 22924 14522 22976
rect 17865 22967 17923 22973
rect 17865 22933 17877 22967
rect 17911 22964 17923 22967
rect 19150 22964 19156 22976
rect 17911 22936 19156 22964
rect 17911 22933 17923 22936
rect 17865 22927 17923 22933
rect 19150 22924 19156 22936
rect 19208 22924 19214 22976
rect 20070 22924 20076 22976
rect 20128 22964 20134 22976
rect 20898 22964 20904 22976
rect 20128 22936 20904 22964
rect 20128 22924 20134 22936
rect 20898 22924 20904 22936
rect 20956 22924 20962 22976
rect 24946 22964 24952 22976
rect 24907 22936 24952 22964
rect 24946 22924 24952 22936
rect 25004 22924 25010 22976
rect 27172 22973 27200 23004
rect 30282 22992 30288 23044
rect 30340 23032 30346 23044
rect 30745 23035 30803 23041
rect 30745 23032 30757 23035
rect 30340 23004 30757 23032
rect 30340 22992 30346 23004
rect 30745 23001 30757 23004
rect 30791 23032 30803 23035
rect 31404 23032 31432 23063
rect 31570 23060 31576 23112
rect 31628 23060 31634 23112
rect 42794 23060 42800 23112
rect 42852 23100 42858 23112
rect 43898 23100 43904 23112
rect 42852 23072 43904 23100
rect 42852 23060 42858 23072
rect 43898 23060 43904 23072
rect 43956 23060 43962 23112
rect 46014 23100 46020 23112
rect 45975 23072 46020 23100
rect 46014 23060 46020 23072
rect 46072 23060 46078 23112
rect 46290 23100 46296 23112
rect 46203 23072 46296 23100
rect 46290 23060 46296 23072
rect 46348 23060 46354 23112
rect 47302 23100 47308 23112
rect 47263 23072 47308 23100
rect 47302 23060 47308 23072
rect 47360 23060 47366 23112
rect 47394 23060 47400 23112
rect 47452 23100 47458 23112
rect 47578 23100 47584 23112
rect 47452 23072 47497 23100
rect 47539 23072 47584 23100
rect 47452 23060 47458 23072
rect 47578 23060 47584 23072
rect 47636 23060 47642 23112
rect 47765 23103 47823 23109
rect 47765 23069 47777 23103
rect 47811 23100 47823 23103
rect 50246 23100 50252 23112
rect 47811 23072 50252 23100
rect 47811 23069 47823 23072
rect 47765 23063 47823 23069
rect 50246 23060 50252 23072
rect 50304 23060 50310 23112
rect 50614 23060 50620 23112
rect 50672 23060 50678 23112
rect 52270 23060 52276 23112
rect 52328 23100 52334 23112
rect 52457 23103 52515 23109
rect 52457 23100 52469 23103
rect 52328 23072 52469 23100
rect 52328 23060 52334 23072
rect 52457 23069 52469 23072
rect 52503 23069 52515 23103
rect 52457 23063 52515 23069
rect 53006 23060 53012 23112
rect 53064 23100 53070 23112
rect 53101 23103 53159 23109
rect 53101 23100 53113 23103
rect 53064 23072 53113 23100
rect 53064 23060 53070 23072
rect 53101 23069 53113 23072
rect 53147 23069 53159 23103
rect 53101 23063 53159 23069
rect 30791 23004 31432 23032
rect 30791 23001 30803 23004
rect 30745 22995 30803 23001
rect 34698 22992 34704 23044
rect 34756 23032 34762 23044
rect 34793 23035 34851 23041
rect 34793 23032 34805 23035
rect 34756 23004 34805 23032
rect 34756 22992 34762 23004
rect 34793 23001 34805 23004
rect 34839 23001 34851 23035
rect 34793 22995 34851 23001
rect 34882 22992 34888 23044
rect 34940 23032 34946 23044
rect 34993 23035 35051 23041
rect 34993 23032 35005 23035
rect 34940 23004 35005 23032
rect 34940 22992 34946 23004
rect 34993 23001 35005 23004
rect 35039 23001 35051 23035
rect 53484 23032 53512 23199
rect 54478 23100 54484 23112
rect 54439 23072 54484 23100
rect 54478 23060 54484 23072
rect 54536 23060 54542 23112
rect 54573 23103 54631 23109
rect 54573 23069 54585 23103
rect 54619 23100 54631 23103
rect 55490 23100 55496 23112
rect 54619 23072 55496 23100
rect 54619 23069 54631 23072
rect 54573 23063 54631 23069
rect 55490 23060 55496 23072
rect 55548 23060 55554 23112
rect 56502 23100 56508 23112
rect 56463 23072 56508 23100
rect 56502 23060 56508 23072
rect 56560 23060 56566 23112
rect 57054 23100 57060 23112
rect 57015 23072 57060 23100
rect 57054 23060 57060 23072
rect 57112 23060 57118 23112
rect 53742 23032 53748 23044
rect 53484 23004 53748 23032
rect 34993 22995 35051 23001
rect 53742 22992 53748 23004
rect 53800 23032 53806 23044
rect 54757 23035 54815 23041
rect 54757 23032 54769 23035
rect 53800 23004 54769 23032
rect 53800 22992 53806 23004
rect 54757 23001 54769 23004
rect 54803 23032 54815 23035
rect 55309 23035 55367 23041
rect 55309 23032 55321 23035
rect 54803 23004 55321 23032
rect 54803 23001 54815 23004
rect 54757 22995 54815 23001
rect 55309 23001 55321 23004
rect 55355 23001 55367 23035
rect 55309 22995 55367 23001
rect 57698 22992 57704 23044
rect 57756 22992 57762 23044
rect 27157 22967 27215 22973
rect 27157 22933 27169 22967
rect 27203 22933 27215 22967
rect 27157 22927 27215 22933
rect 27706 22924 27712 22976
rect 27764 22964 27770 22976
rect 27801 22967 27859 22973
rect 27801 22964 27813 22967
rect 27764 22936 27813 22964
rect 27764 22924 27770 22936
rect 27801 22933 27813 22936
rect 27847 22933 27859 22967
rect 27801 22927 27859 22933
rect 28905 22967 28963 22973
rect 28905 22933 28917 22967
rect 28951 22964 28963 22967
rect 29822 22964 29828 22976
rect 28951 22936 29828 22964
rect 28951 22933 28963 22936
rect 28905 22927 28963 22933
rect 29822 22924 29828 22936
rect 29880 22924 29886 22976
rect 33502 22964 33508 22976
rect 33463 22936 33508 22964
rect 33502 22924 33508 22936
rect 33560 22924 33566 22976
rect 34149 22967 34207 22973
rect 34149 22933 34161 22967
rect 34195 22964 34207 22967
rect 34606 22964 34612 22976
rect 34195 22936 34612 22964
rect 34195 22933 34207 22936
rect 34149 22927 34207 22933
rect 34606 22924 34612 22936
rect 34664 22924 34670 22976
rect 35618 22964 35624 22976
rect 35579 22936 35624 22964
rect 35618 22924 35624 22936
rect 35676 22924 35682 22976
rect 43530 22964 43536 22976
rect 43491 22936 43536 22964
rect 43530 22924 43536 22936
rect 43588 22924 43594 22976
rect 46106 22964 46112 22976
rect 46067 22936 46112 22964
rect 46106 22924 46112 22936
rect 46164 22924 46170 22976
rect 54478 22924 54484 22976
rect 54536 22964 54542 22976
rect 55509 22967 55567 22973
rect 55509 22964 55521 22967
rect 54536 22936 55521 22964
rect 54536 22924 54542 22936
rect 55509 22933 55521 22936
rect 55555 22933 55567 22967
rect 55674 22964 55680 22976
rect 55635 22936 55680 22964
rect 55509 22927 55567 22933
rect 55674 22924 55680 22936
rect 55732 22924 55738 22976
rect 1104 22874 58880 22896
rect 1104 22822 19574 22874
rect 19626 22822 19638 22874
rect 19690 22822 19702 22874
rect 19754 22822 19766 22874
rect 19818 22822 19830 22874
rect 19882 22822 50294 22874
rect 50346 22822 50358 22874
rect 50410 22822 50422 22874
rect 50474 22822 50486 22874
rect 50538 22822 50550 22874
rect 50602 22822 58880 22874
rect 1104 22800 58880 22822
rect 1673 22763 1731 22769
rect 1673 22729 1685 22763
rect 1719 22760 1731 22763
rect 1854 22760 1860 22772
rect 1719 22732 1860 22760
rect 1719 22729 1731 22732
rect 1673 22723 1731 22729
rect 1854 22720 1860 22732
rect 1912 22720 1918 22772
rect 4614 22720 4620 22772
rect 4672 22760 4678 22772
rect 5077 22763 5135 22769
rect 5077 22760 5089 22763
rect 4672 22732 5089 22760
rect 4672 22720 4678 22732
rect 5077 22729 5089 22732
rect 5123 22760 5135 22763
rect 5258 22760 5264 22772
rect 5123 22732 5264 22760
rect 5123 22729 5135 22732
rect 5077 22723 5135 22729
rect 5258 22720 5264 22732
rect 5316 22720 5322 22772
rect 6178 22720 6184 22772
rect 6236 22760 6242 22772
rect 6641 22763 6699 22769
rect 6641 22760 6653 22763
rect 6236 22732 6653 22760
rect 6236 22720 6242 22732
rect 6641 22729 6653 22732
rect 6687 22760 6699 22763
rect 8478 22760 8484 22772
rect 6687 22732 8484 22760
rect 6687 22729 6699 22732
rect 6641 22723 6699 22729
rect 8478 22720 8484 22732
rect 8536 22720 8542 22772
rect 9401 22763 9459 22769
rect 9401 22760 9413 22763
rect 8772 22732 9413 22760
rect 8772 22704 8800 22732
rect 9401 22729 9413 22732
rect 9447 22729 9459 22763
rect 9401 22723 9459 22729
rect 11701 22763 11759 22769
rect 11701 22729 11713 22763
rect 11747 22760 11759 22763
rect 15197 22763 15255 22769
rect 11747 22732 13308 22760
rect 11747 22729 11759 22732
rect 11701 22723 11759 22729
rect 4062 22692 4068 22704
rect 3528 22664 4068 22692
rect 3528 22633 3556 22664
rect 4062 22652 4068 22664
rect 4120 22652 4126 22704
rect 8754 22692 8760 22704
rect 8715 22664 8760 22692
rect 8754 22652 8760 22664
rect 8812 22652 8818 22704
rect 8941 22695 8999 22701
rect 8941 22661 8953 22695
rect 8987 22692 8999 22695
rect 9858 22692 9864 22704
rect 8987 22664 9864 22692
rect 8987 22661 8999 22664
rect 8941 22655 8999 22661
rect 9858 22652 9864 22664
rect 9916 22652 9922 22704
rect 12894 22692 12900 22704
rect 9968 22664 12900 22692
rect 3513 22627 3571 22633
rect 3513 22593 3525 22627
rect 3559 22593 3571 22627
rect 3513 22587 3571 22593
rect 3602 22584 3608 22636
rect 3660 22624 3666 22636
rect 3789 22627 3847 22633
rect 3789 22624 3801 22627
rect 3660 22596 3801 22624
rect 3660 22584 3666 22596
rect 3789 22593 3801 22596
rect 3835 22593 3847 22627
rect 3789 22587 3847 22593
rect 6822 22584 6828 22636
rect 6880 22624 6886 22636
rect 7650 22624 7656 22636
rect 6880 22596 7656 22624
rect 6880 22584 6886 22596
rect 7650 22584 7656 22596
rect 7708 22584 7714 22636
rect 7837 22627 7895 22633
rect 7837 22593 7849 22627
rect 7883 22624 7895 22627
rect 8294 22624 8300 22636
rect 7883 22596 8300 22624
rect 7883 22593 7895 22596
rect 7837 22587 7895 22593
rect 8294 22584 8300 22596
rect 8352 22624 8358 22636
rect 9968 22624 9996 22664
rect 12894 22652 12900 22664
rect 12952 22692 12958 22704
rect 13081 22695 13139 22701
rect 13081 22692 13093 22695
rect 12952 22664 13093 22692
rect 12952 22652 12958 22664
rect 13081 22661 13093 22664
rect 13127 22661 13139 22695
rect 13081 22655 13139 22661
rect 8352 22596 9996 22624
rect 8352 22584 8358 22596
rect 10594 22584 10600 22636
rect 10652 22624 10658 22636
rect 11517 22627 11575 22633
rect 11517 22624 11529 22627
rect 10652 22596 11529 22624
rect 10652 22584 10658 22596
rect 11517 22593 11529 22596
rect 11563 22593 11575 22627
rect 12802 22624 12808 22636
rect 12763 22596 12808 22624
rect 11517 22587 11575 22593
rect 12802 22584 12808 22596
rect 12860 22584 12866 22636
rect 12986 22624 12992 22636
rect 12947 22596 12992 22624
rect 12986 22584 12992 22596
rect 13044 22584 13050 22636
rect 13173 22627 13231 22633
rect 13173 22593 13185 22627
rect 13219 22593 13231 22627
rect 13173 22587 13231 22593
rect 12345 22559 12403 22565
rect 12345 22525 12357 22559
rect 12391 22556 12403 22559
rect 13078 22556 13084 22568
rect 12391 22528 13084 22556
rect 12391 22525 12403 22528
rect 12345 22519 12403 22525
rect 13078 22516 13084 22528
rect 13136 22556 13142 22568
rect 13188 22556 13216 22587
rect 13136 22528 13216 22556
rect 13136 22516 13142 22528
rect 4614 22420 4620 22432
rect 4575 22392 4620 22420
rect 4614 22380 4620 22392
rect 4672 22380 4678 22432
rect 9766 22380 9772 22432
rect 9824 22420 9830 22432
rect 10229 22423 10287 22429
rect 10229 22420 10241 22423
rect 9824 22392 10241 22420
rect 9824 22380 9830 22392
rect 10229 22389 10241 22392
rect 10275 22389 10287 22423
rect 13280 22420 13308 22732
rect 15197 22729 15209 22763
rect 15243 22760 15255 22763
rect 15378 22760 15384 22772
rect 15243 22732 15384 22760
rect 15243 22729 15255 22732
rect 15197 22723 15255 22729
rect 15378 22720 15384 22732
rect 15436 22720 15442 22772
rect 17221 22763 17279 22769
rect 17221 22729 17233 22763
rect 17267 22760 17279 22763
rect 17494 22760 17500 22772
rect 17267 22732 17500 22760
rect 17267 22729 17279 22732
rect 17221 22723 17279 22729
rect 17494 22720 17500 22732
rect 17552 22720 17558 22772
rect 19242 22720 19248 22772
rect 19300 22760 19306 22772
rect 19797 22763 19855 22769
rect 19300 22732 19661 22760
rect 19300 22720 19306 22732
rect 14458 22652 14464 22704
rect 14516 22692 14522 22704
rect 18693 22695 18751 22701
rect 18693 22692 18705 22695
rect 14516 22664 16804 22692
rect 14516 22652 14522 22664
rect 13998 22633 14004 22636
rect 13817 22627 13875 22633
rect 13817 22624 13829 22627
rect 13372 22596 13829 22624
rect 13372 22497 13400 22596
rect 13817 22593 13829 22596
rect 13863 22593 13875 22627
rect 13817 22587 13875 22593
rect 13965 22627 14004 22633
rect 13965 22593 13977 22627
rect 13965 22587 14004 22593
rect 13998 22584 14004 22587
rect 14056 22584 14062 22636
rect 14093 22627 14151 22633
rect 14093 22593 14105 22627
rect 14139 22593 14151 22627
rect 14093 22587 14151 22593
rect 14108 22556 14136 22587
rect 14182 22584 14188 22636
rect 14240 22624 14246 22636
rect 14323 22627 14381 22633
rect 14240 22596 14285 22624
rect 14240 22584 14246 22596
rect 14323 22593 14335 22627
rect 14369 22624 14381 22627
rect 14918 22624 14924 22636
rect 14369 22596 14924 22624
rect 14369 22593 14381 22596
rect 14323 22587 14381 22593
rect 14918 22584 14924 22596
rect 14976 22584 14982 22636
rect 15010 22584 15016 22636
rect 15068 22624 15074 22636
rect 15105 22627 15163 22633
rect 15105 22624 15117 22627
rect 15068 22596 15117 22624
rect 15068 22584 15074 22596
rect 15105 22593 15117 22596
rect 15151 22593 15163 22627
rect 15105 22587 15163 22593
rect 16482 22584 16488 22636
rect 16540 22624 16546 22636
rect 16776 22633 16804 22664
rect 16868 22664 18705 22692
rect 16669 22627 16727 22633
rect 16669 22624 16681 22627
rect 16540 22596 16681 22624
rect 16540 22584 16546 22596
rect 16669 22593 16681 22596
rect 16715 22593 16727 22627
rect 16669 22587 16727 22593
rect 16761 22627 16819 22633
rect 16761 22593 16773 22627
rect 16807 22593 16819 22627
rect 16761 22587 16819 22593
rect 16868 22556 16896 22664
rect 18693 22661 18705 22664
rect 18739 22692 18751 22695
rect 19429 22695 19487 22701
rect 19429 22692 19441 22695
rect 18739 22664 19441 22692
rect 18739 22661 18751 22664
rect 18693 22655 18751 22661
rect 19429 22661 19441 22664
rect 19475 22661 19487 22695
rect 19429 22655 19487 22661
rect 16945 22627 17003 22633
rect 16945 22593 16957 22627
rect 16991 22593 17003 22627
rect 16945 22587 17003 22593
rect 14108 22528 16896 22556
rect 14292 22500 14320 22528
rect 13357 22491 13415 22497
rect 13357 22457 13369 22491
rect 13403 22457 13415 22491
rect 13357 22451 13415 22457
rect 14274 22448 14280 22500
rect 14332 22448 14338 22500
rect 14458 22488 14464 22500
rect 14419 22460 14464 22488
rect 14458 22448 14464 22460
rect 14516 22448 14522 22500
rect 15102 22448 15108 22500
rect 15160 22488 15166 22500
rect 16025 22491 16083 22497
rect 16025 22488 16037 22491
rect 15160 22460 16037 22488
rect 15160 22448 15166 22460
rect 16025 22457 16037 22460
rect 16071 22488 16083 22491
rect 16960 22488 16988 22587
rect 17034 22584 17040 22636
rect 17092 22624 17098 22636
rect 19150 22624 19156 22636
rect 17092 22596 18828 22624
rect 19111 22596 19156 22624
rect 17092 22584 17098 22596
rect 18800 22556 18828 22596
rect 19150 22584 19156 22596
rect 19208 22584 19214 22636
rect 19334 22633 19340 22636
rect 19301 22627 19340 22633
rect 19301 22593 19313 22627
rect 19301 22587 19340 22593
rect 19334 22584 19340 22587
rect 19392 22584 19398 22636
rect 19633 22633 19661 22732
rect 19797 22729 19809 22763
rect 19843 22760 19855 22763
rect 19978 22760 19984 22772
rect 19843 22732 19984 22760
rect 19843 22729 19855 22732
rect 19797 22723 19855 22729
rect 19978 22720 19984 22732
rect 20036 22720 20042 22772
rect 20714 22720 20720 22772
rect 20772 22760 20778 22772
rect 23385 22763 23443 22769
rect 20772 22732 22140 22760
rect 20772 22720 20778 22732
rect 20806 22652 20812 22704
rect 20864 22692 20870 22704
rect 21177 22695 21235 22701
rect 21177 22692 21189 22695
rect 20864 22664 21189 22692
rect 20864 22652 20870 22664
rect 21177 22661 21189 22664
rect 21223 22661 21235 22695
rect 21177 22655 21235 22661
rect 19521 22627 19579 22633
rect 19521 22593 19533 22627
rect 19567 22593 19579 22627
rect 19633 22627 19717 22633
rect 19633 22596 19671 22627
rect 19521 22587 19579 22593
rect 19659 22593 19671 22596
rect 19705 22624 19717 22627
rect 20990 22624 20996 22636
rect 19705 22596 20996 22624
rect 19705 22593 19717 22596
rect 19659 22587 19717 22593
rect 19536 22556 19564 22587
rect 20990 22584 20996 22596
rect 21048 22584 21054 22636
rect 21818 22624 21824 22636
rect 21779 22596 21824 22624
rect 21818 22584 21824 22596
rect 21876 22584 21882 22636
rect 22112 22633 22140 22732
rect 23385 22729 23397 22763
rect 23431 22760 23443 22763
rect 23474 22760 23480 22772
rect 23431 22732 23480 22760
rect 23431 22729 23443 22732
rect 23385 22723 23443 22729
rect 23474 22720 23480 22732
rect 23532 22720 23538 22772
rect 28445 22763 28503 22769
rect 28445 22729 28457 22763
rect 28491 22760 28503 22763
rect 28810 22760 28816 22772
rect 28491 22732 28816 22760
rect 28491 22729 28503 22732
rect 28445 22723 28503 22729
rect 28810 22720 28816 22732
rect 28868 22720 28874 22772
rect 30282 22760 30288 22772
rect 30243 22732 30288 22760
rect 30282 22720 30288 22732
rect 30340 22720 30346 22772
rect 34057 22763 34115 22769
rect 34057 22729 34069 22763
rect 34103 22760 34115 22763
rect 34698 22760 34704 22772
rect 34103 22732 34704 22760
rect 34103 22729 34115 22732
rect 34057 22723 34115 22729
rect 34698 22720 34704 22732
rect 34756 22720 34762 22772
rect 34790 22720 34796 22772
rect 34848 22760 34854 22772
rect 34977 22763 35035 22769
rect 34977 22760 34989 22763
rect 34848 22732 34989 22760
rect 34848 22720 34854 22732
rect 34977 22729 34989 22732
rect 35023 22729 35035 22763
rect 35434 22760 35440 22772
rect 35395 22732 35440 22760
rect 34977 22723 35035 22729
rect 35434 22720 35440 22732
rect 35492 22720 35498 22772
rect 37829 22763 37887 22769
rect 37829 22729 37841 22763
rect 37875 22760 37887 22763
rect 38102 22760 38108 22772
rect 37875 22732 38108 22760
rect 37875 22729 37887 22732
rect 37829 22723 37887 22729
rect 38102 22720 38108 22732
rect 38160 22720 38166 22772
rect 43073 22763 43131 22769
rect 43073 22729 43085 22763
rect 43119 22760 43131 22763
rect 43530 22760 43536 22772
rect 43119 22732 43536 22760
rect 43119 22729 43131 22732
rect 43073 22723 43131 22729
rect 43530 22720 43536 22732
rect 43588 22720 43594 22772
rect 46014 22720 46020 22772
rect 46072 22760 46078 22772
rect 46493 22763 46551 22769
rect 46493 22760 46505 22763
rect 46072 22732 46505 22760
rect 46072 22720 46078 22732
rect 46493 22729 46505 22732
rect 46539 22729 46551 22763
rect 46493 22723 46551 22729
rect 46661 22763 46719 22769
rect 46661 22729 46673 22763
rect 46707 22760 46719 22763
rect 47578 22760 47584 22772
rect 46707 22732 47584 22760
rect 46707 22729 46719 22732
rect 46661 22723 46719 22729
rect 47578 22720 47584 22732
rect 47636 22720 47642 22772
rect 52822 22720 52828 22772
rect 52880 22760 52886 22772
rect 53377 22763 53435 22769
rect 53377 22760 53389 22763
rect 52880 22732 53389 22760
rect 52880 22720 52886 22732
rect 53377 22729 53389 22732
rect 53423 22729 53435 22763
rect 57054 22760 57060 22772
rect 57015 22732 57060 22760
rect 53377 22723 53435 22729
rect 57054 22720 57060 22732
rect 57112 22720 57118 22772
rect 24581 22695 24639 22701
rect 24581 22692 24593 22695
rect 24044 22664 24593 22692
rect 24044 22636 24072 22664
rect 24581 22661 24593 22664
rect 24627 22661 24639 22695
rect 24581 22655 24639 22661
rect 33502 22652 33508 22704
rect 33560 22692 33566 22704
rect 35618 22692 35624 22704
rect 33560 22664 35624 22692
rect 33560 22652 33566 22664
rect 21913 22627 21971 22633
rect 21913 22593 21925 22627
rect 21959 22593 21971 22627
rect 21913 22587 21971 22593
rect 22097 22627 22155 22633
rect 22097 22593 22109 22627
rect 22143 22593 22155 22627
rect 22097 22587 22155 22593
rect 20346 22556 20352 22568
rect 18800 22528 20352 22556
rect 20346 22516 20352 22528
rect 20404 22516 20410 22568
rect 20622 22516 20628 22568
rect 20680 22556 20686 22568
rect 21928 22556 21956 22587
rect 22186 22584 22192 22636
rect 22244 22624 22250 22636
rect 22244 22596 22289 22624
rect 22244 22584 22250 22596
rect 23566 22584 23572 22636
rect 23624 22624 23630 22636
rect 23845 22627 23903 22633
rect 23845 22624 23857 22627
rect 23624 22596 23857 22624
rect 23624 22584 23630 22596
rect 23845 22593 23857 22596
rect 23891 22593 23903 22627
rect 23845 22587 23903 22593
rect 23937 22627 23995 22633
rect 23937 22593 23949 22627
rect 23983 22624 23995 22627
rect 24026 22624 24032 22636
rect 23983 22596 24032 22624
rect 23983 22593 23995 22596
rect 23937 22587 23995 22593
rect 24026 22584 24032 22596
rect 24084 22584 24090 22636
rect 24121 22627 24179 22633
rect 24121 22593 24133 22627
rect 24167 22624 24179 22627
rect 24210 22624 24216 22636
rect 24167 22596 24216 22624
rect 24167 22593 24179 22596
rect 24121 22587 24179 22593
rect 24210 22584 24216 22596
rect 24268 22624 24274 22636
rect 24486 22624 24492 22636
rect 24268 22596 24492 22624
rect 24268 22584 24274 22596
rect 24486 22584 24492 22596
rect 24544 22624 24550 22636
rect 25133 22627 25191 22633
rect 25133 22624 25145 22627
rect 24544 22596 25145 22624
rect 24544 22584 24550 22596
rect 25133 22593 25145 22596
rect 25179 22593 25191 22627
rect 25133 22587 25191 22593
rect 28077 22627 28135 22633
rect 28077 22593 28089 22627
rect 28123 22593 28135 22627
rect 28077 22587 28135 22593
rect 20680 22528 21956 22556
rect 22373 22559 22431 22565
rect 20680 22516 20686 22528
rect 22373 22525 22385 22559
rect 22419 22556 22431 22559
rect 27985 22559 28043 22565
rect 27985 22556 27997 22559
rect 22419 22528 27997 22556
rect 22419 22525 22431 22528
rect 22373 22519 22431 22525
rect 27985 22525 27997 22528
rect 28031 22525 28043 22559
rect 27985 22519 28043 22525
rect 23658 22488 23664 22500
rect 16071 22460 23664 22488
rect 16071 22457 16083 22460
rect 16025 22451 16083 22457
rect 23658 22448 23664 22460
rect 23716 22448 23722 22500
rect 28092 22488 28120 22587
rect 29822 22584 29828 22636
rect 29880 22624 29886 22636
rect 30193 22627 30251 22633
rect 30193 22624 30205 22627
rect 29880 22596 30205 22624
rect 29880 22584 29886 22596
rect 30193 22593 30205 22596
rect 30239 22593 30251 22627
rect 30374 22624 30380 22636
rect 30335 22596 30380 22624
rect 30193 22587 30251 22593
rect 30374 22584 30380 22596
rect 30432 22584 30438 22636
rect 32950 22584 32956 22636
rect 33008 22624 33014 22636
rect 34532 22633 34560 22664
rect 35618 22652 35624 22664
rect 35676 22692 35682 22704
rect 35713 22695 35771 22701
rect 35713 22692 35725 22695
rect 35676 22664 35725 22692
rect 35676 22652 35682 22664
rect 35713 22661 35725 22664
rect 35759 22661 35771 22695
rect 46290 22692 46296 22704
rect 46251 22664 46296 22692
rect 35713 22655 35771 22661
rect 46290 22652 46296 22664
rect 46348 22652 46354 22704
rect 50341 22695 50399 22701
rect 50341 22661 50353 22695
rect 50387 22692 50399 22695
rect 50614 22692 50620 22704
rect 50387 22664 50620 22692
rect 50387 22661 50399 22664
rect 50341 22655 50399 22661
rect 50614 22652 50620 22664
rect 50672 22652 50678 22704
rect 52270 22652 52276 22704
rect 52328 22692 52334 22704
rect 52328 22664 52960 22692
rect 52328 22652 52334 22664
rect 33045 22627 33103 22633
rect 33045 22624 33057 22627
rect 33008 22596 33057 22624
rect 33008 22584 33014 22596
rect 33045 22593 33057 22596
rect 33091 22624 33103 22627
rect 33689 22627 33747 22633
rect 33689 22624 33701 22627
rect 33091 22596 33701 22624
rect 33091 22593 33103 22596
rect 33045 22587 33103 22593
rect 33689 22593 33701 22596
rect 33735 22593 33747 22627
rect 33689 22587 33747 22593
rect 34517 22627 34575 22633
rect 34517 22593 34529 22627
rect 34563 22593 34575 22627
rect 34517 22587 34575 22593
rect 34606 22584 34612 22636
rect 34664 22624 34670 22636
rect 34793 22627 34851 22633
rect 34664 22596 34709 22624
rect 34664 22584 34670 22596
rect 34793 22593 34805 22627
rect 34839 22593 34851 22627
rect 35434 22624 35440 22636
rect 35395 22596 35440 22624
rect 34793 22587 34851 22593
rect 33318 22516 33324 22568
rect 33376 22556 33382 22568
rect 33597 22559 33655 22565
rect 33597 22556 33609 22559
rect 33376 22528 33609 22556
rect 33376 22516 33382 22528
rect 33597 22525 33609 22528
rect 33643 22525 33655 22559
rect 34808 22556 34836 22587
rect 35434 22584 35440 22596
rect 35492 22584 35498 22636
rect 35529 22627 35587 22633
rect 35529 22593 35541 22627
rect 35575 22624 35587 22627
rect 35575 22596 35756 22624
rect 35575 22593 35587 22596
rect 35529 22587 35587 22593
rect 33597 22519 33655 22525
rect 34532 22528 34836 22556
rect 33502 22488 33508 22500
rect 28092 22460 33508 22488
rect 33502 22448 33508 22460
rect 33560 22448 33566 22500
rect 15930 22420 15936 22432
rect 13280 22392 15936 22420
rect 10229 22383 10287 22389
rect 15930 22380 15936 22392
rect 15988 22380 15994 22432
rect 21085 22423 21143 22429
rect 21085 22389 21097 22423
rect 21131 22420 21143 22423
rect 22002 22420 22008 22432
rect 21131 22392 22008 22420
rect 21131 22389 21143 22392
rect 21085 22383 21143 22389
rect 22002 22380 22008 22392
rect 22060 22380 22066 22432
rect 24121 22423 24179 22429
rect 24121 22389 24133 22423
rect 24167 22420 24179 22423
rect 24394 22420 24400 22432
rect 24167 22392 24400 22420
rect 24167 22389 24179 22392
rect 24121 22383 24179 22389
rect 24394 22380 24400 22392
rect 24452 22380 24458 22432
rect 33612 22420 33640 22519
rect 34532 22500 34560 22528
rect 34514 22448 34520 22500
rect 34572 22448 34578 22500
rect 34606 22448 34612 22500
rect 34664 22488 34670 22500
rect 35728 22488 35756 22596
rect 35802 22584 35808 22636
rect 35860 22624 35866 22636
rect 37461 22627 37519 22633
rect 37461 22624 37473 22627
rect 35860 22596 37473 22624
rect 35860 22584 35866 22596
rect 37461 22593 37473 22596
rect 37507 22624 37519 22627
rect 38930 22624 38936 22636
rect 37507 22596 38936 22624
rect 37507 22593 37519 22596
rect 37461 22587 37519 22593
rect 38930 22584 38936 22596
rect 38988 22584 38994 22636
rect 40218 22624 40224 22636
rect 40179 22596 40224 22624
rect 40218 22584 40224 22596
rect 40276 22584 40282 22636
rect 42518 22624 42524 22636
rect 42479 22596 42524 22624
rect 42518 22584 42524 22596
rect 42576 22584 42582 22636
rect 42889 22627 42947 22633
rect 42889 22593 42901 22627
rect 42935 22624 42947 22627
rect 42978 22624 42984 22636
rect 42935 22596 42984 22624
rect 42935 22593 42947 22596
rect 42889 22587 42947 22593
rect 42978 22584 42984 22596
rect 43036 22584 43042 22636
rect 49326 22624 49332 22636
rect 49287 22596 49332 22624
rect 49326 22584 49332 22596
rect 49384 22584 49390 22636
rect 49694 22584 49700 22636
rect 49752 22584 49758 22636
rect 52086 22584 52092 22636
rect 52144 22624 52150 22636
rect 52932 22633 52960 22664
rect 53742 22652 53748 22704
rect 53800 22692 53806 22704
rect 54481 22695 54539 22701
rect 54481 22692 54493 22695
rect 53800 22664 54493 22692
rect 53800 22652 53806 22664
rect 54481 22661 54493 22664
rect 54527 22661 54539 22695
rect 56502 22692 56508 22704
rect 56463 22664 56508 22692
rect 54481 22655 54539 22661
rect 56502 22652 56508 22664
rect 56560 22652 56566 22704
rect 52733 22627 52791 22633
rect 52733 22624 52745 22627
rect 52144 22596 52745 22624
rect 52144 22584 52150 22596
rect 52733 22593 52745 22596
rect 52779 22593 52791 22627
rect 52733 22587 52791 22593
rect 52917 22627 52975 22633
rect 52917 22593 52929 22627
rect 52963 22593 52975 22627
rect 52917 22587 52975 22593
rect 53006 22584 53012 22636
rect 53064 22624 53070 22636
rect 53147 22627 53205 22633
rect 53064 22596 53109 22624
rect 53064 22584 53070 22596
rect 53147 22593 53159 22627
rect 53193 22624 53205 22627
rect 53282 22624 53288 22636
rect 53193 22596 53288 22624
rect 53193 22593 53205 22596
rect 53147 22587 53205 22593
rect 53282 22584 53288 22596
rect 53340 22584 53346 22636
rect 53650 22584 53656 22636
rect 53708 22624 53714 22636
rect 54757 22627 54815 22633
rect 54757 22624 54769 22627
rect 53708 22596 54769 22624
rect 53708 22584 53714 22596
rect 54757 22593 54769 22596
rect 54803 22593 54815 22627
rect 54757 22587 54815 22593
rect 55125 22627 55183 22633
rect 55125 22593 55137 22627
rect 55171 22593 55183 22627
rect 55125 22587 55183 22593
rect 55217 22627 55275 22633
rect 55217 22593 55229 22627
rect 55263 22624 55275 22627
rect 56226 22624 56232 22636
rect 55263 22596 56232 22624
rect 55263 22593 55275 22596
rect 55217 22587 55275 22593
rect 37369 22559 37427 22565
rect 37369 22525 37381 22559
rect 37415 22525 37427 22559
rect 40126 22556 40132 22568
rect 40087 22528 40132 22556
rect 37369 22519 37427 22525
rect 36630 22488 36636 22500
rect 34664 22460 35756 22488
rect 36591 22460 36636 22488
rect 34664 22448 34670 22460
rect 36630 22448 36636 22460
rect 36688 22488 36694 22500
rect 37384 22488 37412 22519
rect 40126 22516 40132 22528
rect 40184 22516 40190 22568
rect 40586 22556 40592 22568
rect 40547 22528 40592 22556
rect 40586 22516 40592 22528
rect 40644 22516 40650 22568
rect 55140 22556 55168 22587
rect 56226 22584 56232 22596
rect 56284 22584 56290 22636
rect 56318 22584 56324 22636
rect 56376 22624 56382 22636
rect 56376 22596 56421 22624
rect 56376 22584 56382 22596
rect 56686 22584 56692 22636
rect 56744 22624 56750 22636
rect 56965 22627 57023 22633
rect 56965 22624 56977 22627
rect 56744 22596 56977 22624
rect 56744 22584 56750 22596
rect 56965 22593 56977 22596
rect 57011 22593 57023 22627
rect 57146 22624 57152 22636
rect 57107 22596 57152 22624
rect 56965 22587 57023 22593
rect 57146 22584 57152 22596
rect 57204 22584 57210 22636
rect 55490 22556 55496 22568
rect 55140 22528 55496 22556
rect 55490 22516 55496 22528
rect 55548 22516 55554 22568
rect 36688 22460 37412 22488
rect 36688 22448 36694 22460
rect 54478 22448 54484 22500
rect 54536 22488 54542 22500
rect 55309 22491 55367 22497
rect 55309 22488 55321 22491
rect 54536 22460 55321 22488
rect 54536 22448 54542 22460
rect 55309 22457 55321 22460
rect 55355 22457 55367 22491
rect 55309 22451 55367 22457
rect 36722 22420 36728 22432
rect 33612 22392 36728 22420
rect 36722 22380 36728 22392
rect 36780 22380 36786 22432
rect 42886 22420 42892 22432
rect 42847 22392 42892 22420
rect 42886 22380 42892 22392
rect 42944 22380 42950 22432
rect 46106 22380 46112 22432
rect 46164 22420 46170 22432
rect 46477 22423 46535 22429
rect 46477 22420 46489 22423
rect 46164 22392 46489 22420
rect 46164 22380 46170 22392
rect 46477 22389 46489 22392
rect 46523 22420 46535 22423
rect 46566 22420 46572 22432
rect 46523 22392 46572 22420
rect 46523 22389 46535 22392
rect 46477 22383 46535 22389
rect 46566 22380 46572 22392
rect 46624 22380 46630 22432
rect 1104 22330 58880 22352
rect 1104 22278 4214 22330
rect 4266 22278 4278 22330
rect 4330 22278 4342 22330
rect 4394 22278 4406 22330
rect 4458 22278 4470 22330
rect 4522 22278 34934 22330
rect 34986 22278 34998 22330
rect 35050 22278 35062 22330
rect 35114 22278 35126 22330
rect 35178 22278 35190 22330
rect 35242 22278 58880 22330
rect 1104 22256 58880 22278
rect 9309 22219 9367 22225
rect 9309 22185 9321 22219
rect 9355 22216 9367 22219
rect 10594 22216 10600 22228
rect 9355 22188 10600 22216
rect 9355 22185 9367 22188
rect 9309 22179 9367 22185
rect 10594 22176 10600 22188
rect 10652 22176 10658 22228
rect 13078 22176 13084 22228
rect 13136 22216 13142 22228
rect 13354 22216 13360 22228
rect 13136 22188 13360 22216
rect 13136 22176 13142 22188
rect 13354 22176 13360 22188
rect 13412 22176 13418 22228
rect 13722 22176 13728 22228
rect 13780 22216 13786 22228
rect 15746 22216 15752 22228
rect 13780 22188 15752 22216
rect 13780 22176 13786 22188
rect 15746 22176 15752 22188
rect 15804 22176 15810 22228
rect 16482 22176 16488 22228
rect 16540 22216 16546 22228
rect 16577 22219 16635 22225
rect 16577 22216 16589 22219
rect 16540 22188 16589 22216
rect 16540 22176 16546 22188
rect 16577 22185 16589 22188
rect 16623 22185 16635 22219
rect 16577 22179 16635 22185
rect 20622 22176 20628 22228
rect 20680 22216 20686 22228
rect 20717 22219 20775 22225
rect 20717 22216 20729 22219
rect 20680 22188 20729 22216
rect 20680 22176 20686 22188
rect 20717 22185 20729 22188
rect 20763 22185 20775 22219
rect 20717 22179 20775 22185
rect 21729 22219 21787 22225
rect 21729 22185 21741 22219
rect 21775 22216 21787 22219
rect 21818 22216 21824 22228
rect 21775 22188 21824 22216
rect 21775 22185 21787 22188
rect 21729 22179 21787 22185
rect 21818 22176 21824 22188
rect 21876 22176 21882 22228
rect 23106 22176 23112 22228
rect 23164 22216 23170 22228
rect 23661 22219 23719 22225
rect 23661 22216 23673 22219
rect 23164 22188 23673 22216
rect 23164 22176 23170 22188
rect 23661 22185 23673 22188
rect 23707 22185 23719 22219
rect 24949 22219 25007 22225
rect 23661 22179 23719 22185
rect 23768 22188 24164 22216
rect 7466 22148 7472 22160
rect 4264 22120 5212 22148
rect 7427 22120 7472 22148
rect 4264 22080 4292 22120
rect 5184 22080 5212 22120
rect 7466 22108 7472 22120
rect 7524 22108 7530 22160
rect 8389 22151 8447 22157
rect 8389 22117 8401 22151
rect 8435 22148 8447 22151
rect 8435 22120 9996 22148
rect 8435 22117 8447 22120
rect 8389 22111 8447 22117
rect 7285 22083 7343 22089
rect 7285 22080 7297 22083
rect 3068 22052 4292 22080
rect 4356 22052 5120 22080
rect 5184 22052 7297 22080
rect 1857 22015 1915 22021
rect 1857 21981 1869 22015
rect 1903 22012 1915 22015
rect 2130 22012 2136 22024
rect 1903 21984 2136 22012
rect 1903 21981 1915 21984
rect 1857 21975 1915 21981
rect 2130 21972 2136 21984
rect 2188 22012 2194 22024
rect 2317 22015 2375 22021
rect 2317 22012 2329 22015
rect 2188 21984 2329 22012
rect 2188 21972 2194 21984
rect 2317 21981 2329 21984
rect 2363 21981 2375 22015
rect 2317 21975 2375 21981
rect 2501 22015 2559 22021
rect 2501 21981 2513 22015
rect 2547 21981 2559 22015
rect 2501 21975 2559 21981
rect 2516 21944 2544 21975
rect 2774 21972 2780 22024
rect 2832 22012 2838 22024
rect 3068 22021 3096 22052
rect 4356 22021 4384 22052
rect 5092 22024 5120 22052
rect 7285 22049 7297 22052
rect 7331 22080 7343 22083
rect 9858 22080 9864 22092
rect 7331 22052 9864 22080
rect 7331 22049 7343 22052
rect 7285 22043 7343 22049
rect 9858 22040 9864 22052
rect 9916 22040 9922 22092
rect 9968 22080 9996 22120
rect 12894 22108 12900 22160
rect 12952 22148 12958 22160
rect 17586 22148 17592 22160
rect 12952 22120 17592 22148
rect 12952 22108 12958 22120
rect 17586 22108 17592 22120
rect 17644 22108 17650 22160
rect 19426 22108 19432 22160
rect 19484 22148 19490 22160
rect 23768 22148 23796 22188
rect 19484 22120 23796 22148
rect 23845 22151 23903 22157
rect 19484 22108 19490 22120
rect 23845 22117 23857 22151
rect 23891 22117 23903 22151
rect 24136 22148 24164 22188
rect 24949 22185 24961 22219
rect 24995 22216 25007 22219
rect 33594 22216 33600 22228
rect 24995 22188 33600 22216
rect 24995 22185 25007 22188
rect 24949 22179 25007 22185
rect 33594 22176 33600 22188
rect 33652 22176 33658 22228
rect 34885 22219 34943 22225
rect 34885 22185 34897 22219
rect 34931 22216 34943 22219
rect 35434 22216 35440 22228
rect 34931 22188 35440 22216
rect 34931 22185 34943 22188
rect 34885 22179 34943 22185
rect 35434 22176 35440 22188
rect 35492 22216 35498 22228
rect 35802 22216 35808 22228
rect 35492 22188 35808 22216
rect 35492 22176 35498 22188
rect 35802 22176 35808 22188
rect 35860 22176 35866 22228
rect 37182 22216 37188 22228
rect 37143 22188 37188 22216
rect 37182 22176 37188 22188
rect 37240 22176 37246 22228
rect 40126 22176 40132 22228
rect 40184 22176 40190 22228
rect 42518 22216 42524 22228
rect 42479 22188 42524 22216
rect 42518 22176 42524 22188
rect 42576 22176 42582 22228
rect 42794 22216 42800 22228
rect 42755 22188 42800 22216
rect 42794 22176 42800 22188
rect 42852 22176 42858 22228
rect 46014 22176 46020 22228
rect 46072 22216 46078 22228
rect 46109 22219 46167 22225
rect 46109 22216 46121 22219
rect 46072 22188 46121 22216
rect 46072 22176 46078 22188
rect 46109 22185 46121 22188
rect 46155 22185 46167 22219
rect 46566 22216 46572 22228
rect 46527 22188 46572 22216
rect 46109 22179 46167 22185
rect 46566 22176 46572 22188
rect 46624 22176 46630 22228
rect 27798 22148 27804 22160
rect 24136 22120 27804 22148
rect 23845 22111 23903 22117
rect 10870 22080 10876 22092
rect 9968 22052 10876 22080
rect 3053 22015 3111 22021
rect 3053 22012 3065 22015
rect 2832 21984 3065 22012
rect 2832 21972 2838 21984
rect 3053 21981 3065 21984
rect 3099 21981 3111 22015
rect 3237 22015 3295 22021
rect 3237 22012 3249 22015
rect 3053 21975 3111 21981
rect 3160 21984 3249 22012
rect 2866 21944 2872 21956
rect 2516 21916 2872 21944
rect 2866 21904 2872 21916
rect 2924 21944 2930 21956
rect 3160 21944 3188 21984
rect 3237 21981 3249 21984
rect 3283 21981 3295 22015
rect 3237 21975 3295 21981
rect 4341 22015 4399 22021
rect 4341 21981 4353 22015
rect 4387 21981 4399 22015
rect 4341 21975 4399 21981
rect 4617 22015 4675 22021
rect 4617 21981 4629 22015
rect 4663 22012 4675 22015
rect 4890 22012 4896 22024
rect 4663 21984 4896 22012
rect 4663 21981 4675 21984
rect 4617 21975 4675 21981
rect 4890 21972 4896 21984
rect 4948 21972 4954 22024
rect 5074 21972 5080 22024
rect 5132 22012 5138 22024
rect 5261 22015 5319 22021
rect 5132 21984 5225 22012
rect 5132 21972 5138 21984
rect 5261 21981 5273 22015
rect 5307 21981 5319 22015
rect 5261 21975 5319 21981
rect 5276 21944 5304 21975
rect 7098 21972 7104 22024
rect 7156 22012 7162 22024
rect 7469 22015 7527 22021
rect 7469 22012 7481 22015
rect 7156 21984 7481 22012
rect 7156 21972 7162 21984
rect 7469 21981 7481 21984
rect 7515 22012 7527 22015
rect 7650 22012 7656 22024
rect 7515 21984 7656 22012
rect 7515 21981 7527 21984
rect 7469 21975 7527 21981
rect 7650 21972 7656 21984
rect 7708 21972 7714 22024
rect 7837 22015 7895 22021
rect 7837 21981 7849 22015
rect 7883 22012 7895 22015
rect 8018 22012 8024 22024
rect 7883 21984 8024 22012
rect 7883 21981 7895 21984
rect 7837 21975 7895 21981
rect 8018 21972 8024 21984
rect 8076 21972 8082 22024
rect 9398 21972 9404 22024
rect 9456 21972 9462 22024
rect 9950 22012 9956 22024
rect 9911 21984 9956 22012
rect 9950 21972 9956 21984
rect 10008 21972 10014 22024
rect 10042 21972 10048 22024
rect 10100 22012 10106 22024
rect 10244 22021 10272 22052
rect 10870 22040 10876 22052
rect 10928 22040 10934 22092
rect 12805 22083 12863 22089
rect 12805 22049 12817 22083
rect 12851 22080 12863 22083
rect 14274 22080 14280 22092
rect 12851 22052 14280 22080
rect 12851 22049 12863 22052
rect 12805 22043 12863 22049
rect 14274 22040 14280 22052
rect 14332 22040 14338 22092
rect 14645 22083 14703 22089
rect 14645 22049 14657 22083
rect 14691 22080 14703 22083
rect 14918 22080 14924 22092
rect 14691 22052 14924 22080
rect 14691 22049 14703 22052
rect 14645 22043 14703 22049
rect 14918 22040 14924 22052
rect 14976 22040 14982 22092
rect 15010 22040 15016 22092
rect 15068 22080 15074 22092
rect 21818 22080 21824 22092
rect 15068 22052 21824 22080
rect 15068 22040 15074 22052
rect 21818 22040 21824 22052
rect 21876 22040 21882 22092
rect 23860 22080 23888 22111
rect 27798 22108 27804 22120
rect 27856 22108 27862 22160
rect 33502 22108 33508 22160
rect 33560 22148 33566 22160
rect 34790 22148 34796 22160
rect 33560 22120 34796 22148
rect 33560 22108 33566 22120
rect 34790 22108 34796 22120
rect 34848 22148 34854 22160
rect 35342 22148 35348 22160
rect 34848 22120 35348 22148
rect 34848 22108 34854 22120
rect 35342 22108 35348 22120
rect 35400 22108 35406 22160
rect 39301 22151 39359 22157
rect 39301 22117 39313 22151
rect 39347 22148 39359 22151
rect 40144 22148 40172 22176
rect 40589 22151 40647 22157
rect 40589 22148 40601 22151
rect 39347 22120 40601 22148
rect 39347 22117 39359 22120
rect 39301 22111 39359 22117
rect 40589 22117 40601 22120
rect 40635 22117 40647 22151
rect 40589 22111 40647 22117
rect 30558 22080 30564 22092
rect 23860 22052 24532 22080
rect 30519 22052 30564 22080
rect 10229 22015 10287 22021
rect 10100 21984 10145 22012
rect 10100 21972 10106 21984
rect 10229 21981 10241 22015
rect 10275 21981 10287 22015
rect 10229 21975 10287 21981
rect 10321 22015 10379 22021
rect 10321 21981 10333 22015
rect 10367 22012 10379 22015
rect 10778 22012 10784 22024
rect 10367 21984 10784 22012
rect 10367 21981 10379 21984
rect 10321 21975 10379 21981
rect 10778 21972 10784 21984
rect 10836 21972 10842 22024
rect 11054 22012 11060 22024
rect 11015 21984 11060 22012
rect 11054 21972 11060 21984
rect 11112 21972 11118 22024
rect 13170 21972 13176 22024
rect 13228 22012 13234 22024
rect 13449 22015 13507 22021
rect 13449 22012 13461 22015
rect 13228 21984 13461 22012
rect 13228 21972 13234 21984
rect 13449 21981 13461 21984
rect 13495 21981 13507 22015
rect 13449 21975 13507 21981
rect 13538 21972 13544 22024
rect 13596 22012 13602 22024
rect 14093 22015 14151 22021
rect 14093 22012 14105 22015
rect 13596 21984 14105 22012
rect 13596 21972 13602 21984
rect 14093 21981 14105 21984
rect 14139 21981 14151 22015
rect 14093 21975 14151 21981
rect 14461 22015 14519 22021
rect 14461 21981 14473 22015
rect 14507 22012 14519 22015
rect 16298 22012 16304 22024
rect 14507 21984 16304 22012
rect 14507 21981 14519 21984
rect 14461 21975 14519 21981
rect 16298 21972 16304 21984
rect 16356 21972 16362 22024
rect 19886 22012 19892 22024
rect 16408 21984 19892 22012
rect 2924 21916 3188 21944
rect 3988 21916 5304 21944
rect 9125 21947 9183 21953
rect 2924 21904 2930 21916
rect 2501 21879 2559 21885
rect 2501 21845 2513 21879
rect 2547 21876 2559 21879
rect 2682 21876 2688 21888
rect 2547 21848 2688 21876
rect 2547 21845 2559 21848
rect 2501 21839 2559 21845
rect 2682 21836 2688 21848
rect 2740 21836 2746 21888
rect 3142 21876 3148 21888
rect 3103 21848 3148 21876
rect 3142 21836 3148 21848
rect 3200 21876 3206 21888
rect 3988 21876 4016 21916
rect 9125 21913 9137 21947
rect 9171 21944 9183 21947
rect 9416 21944 9444 21972
rect 9171 21916 9444 21944
rect 9171 21913 9183 21916
rect 9125 21907 9183 21913
rect 15746 21904 15752 21956
rect 15804 21944 15810 21956
rect 16408 21953 16436 21984
rect 19886 21972 19892 21984
rect 19944 21972 19950 22024
rect 20073 22015 20131 22021
rect 20073 21981 20085 22015
rect 20119 22012 20131 22015
rect 20533 22015 20591 22021
rect 20533 22012 20545 22015
rect 20119 21984 20545 22012
rect 20119 21981 20131 21984
rect 20073 21975 20131 21981
rect 20533 21981 20545 21984
rect 20579 22012 20591 22015
rect 20622 22012 20628 22024
rect 20579 21984 20628 22012
rect 20579 21981 20591 21984
rect 20533 21975 20591 21981
rect 20622 21972 20628 21984
rect 20680 21972 20686 22024
rect 20714 21972 20720 22024
rect 20772 22012 20778 22024
rect 21177 22015 21235 22021
rect 20772 21984 20817 22012
rect 20772 21972 20778 21984
rect 21177 21981 21189 22015
rect 21223 21981 21235 22015
rect 21450 22012 21456 22024
rect 21411 21984 21456 22012
rect 21177 21975 21235 21981
rect 16393 21947 16451 21953
rect 16393 21944 16405 21947
rect 15804 21916 16405 21944
rect 15804 21904 15810 21916
rect 16393 21913 16405 21916
rect 16439 21913 16451 21947
rect 16393 21907 16451 21913
rect 16482 21904 16488 21956
rect 16540 21944 16546 21956
rect 16577 21947 16635 21953
rect 16577 21944 16589 21947
rect 16540 21916 16589 21944
rect 16540 21904 16546 21916
rect 16577 21913 16589 21916
rect 16623 21944 16635 21947
rect 16623 21916 20300 21944
rect 16623 21913 16635 21916
rect 16577 21907 16635 21913
rect 4154 21876 4160 21888
rect 3200 21848 4016 21876
rect 4115 21848 4160 21876
rect 3200 21836 3206 21848
rect 4154 21836 4160 21848
rect 4212 21836 4218 21888
rect 4525 21879 4583 21885
rect 4525 21845 4537 21879
rect 4571 21876 4583 21879
rect 5353 21879 5411 21885
rect 5353 21876 5365 21879
rect 4571 21848 5365 21876
rect 4571 21845 4583 21848
rect 4525 21839 4583 21845
rect 5353 21845 5365 21848
rect 5399 21876 5411 21879
rect 6730 21876 6736 21888
rect 5399 21848 6736 21876
rect 5399 21845 5411 21848
rect 5353 21839 5411 21845
rect 6730 21836 6736 21848
rect 6788 21836 6794 21888
rect 9306 21836 9312 21888
rect 9364 21885 9370 21888
rect 9364 21879 9383 21885
rect 9371 21845 9383 21879
rect 9364 21839 9383 21845
rect 9493 21879 9551 21885
rect 9493 21845 9505 21879
rect 9539 21876 9551 21879
rect 10042 21876 10048 21888
rect 9539 21848 10048 21876
rect 9539 21845 9551 21848
rect 9493 21839 9551 21845
rect 9364 21836 9370 21839
rect 10042 21836 10048 21848
rect 10100 21836 10106 21888
rect 10502 21876 10508 21888
rect 10463 21848 10508 21876
rect 10502 21836 10508 21848
rect 10560 21836 10566 21888
rect 11238 21876 11244 21888
rect 11199 21848 11244 21876
rect 11238 21836 11244 21848
rect 11296 21836 11302 21888
rect 13170 21836 13176 21888
rect 13228 21876 13234 21888
rect 13357 21879 13415 21885
rect 13357 21876 13369 21879
rect 13228 21848 13369 21876
rect 13228 21836 13234 21848
rect 13357 21845 13369 21848
rect 13403 21845 13415 21879
rect 13357 21839 13415 21845
rect 14461 21879 14519 21885
rect 14461 21845 14473 21879
rect 14507 21876 14519 21879
rect 15194 21876 15200 21888
rect 14507 21848 15200 21876
rect 14507 21845 14519 21848
rect 14461 21839 14519 21845
rect 15194 21836 15200 21848
rect 15252 21836 15258 21888
rect 19334 21836 19340 21888
rect 19392 21876 19398 21888
rect 20162 21876 20168 21888
rect 19392 21848 20168 21876
rect 19392 21836 19398 21848
rect 20162 21836 20168 21848
rect 20220 21836 20226 21888
rect 20272 21876 20300 21916
rect 21082 21876 21088 21888
rect 20272 21848 21088 21876
rect 21082 21836 21088 21848
rect 21140 21836 21146 21888
rect 21192 21876 21220 21975
rect 21450 21972 21456 21984
rect 21508 21972 21514 22024
rect 21542 21972 21548 22024
rect 21600 22012 21606 22024
rect 21600 21984 21645 22012
rect 21600 21972 21606 21984
rect 23658 21972 23664 22024
rect 23716 22012 23722 22024
rect 24394 22012 24400 22024
rect 23716 21984 24256 22012
rect 24355 21984 24400 22012
rect 23716 21972 23722 21984
rect 21358 21904 21364 21956
rect 21416 21944 21422 21956
rect 21726 21944 21732 21956
rect 21416 21916 21732 21944
rect 21416 21904 21422 21916
rect 21726 21904 21732 21916
rect 21784 21904 21790 21956
rect 23477 21947 23535 21953
rect 23477 21913 23489 21947
rect 23523 21944 23535 21947
rect 24118 21944 24124 21956
rect 23523 21916 24124 21944
rect 23523 21913 23535 21916
rect 23477 21907 23535 21913
rect 21634 21876 21640 21888
rect 21192 21848 21640 21876
rect 21634 21836 21640 21848
rect 21692 21836 21698 21888
rect 22094 21836 22100 21888
rect 22152 21876 22158 21888
rect 22925 21879 22983 21885
rect 22925 21876 22937 21879
rect 22152 21848 22937 21876
rect 22152 21836 22158 21848
rect 22925 21845 22937 21848
rect 22971 21876 22983 21879
rect 23492 21876 23520 21907
rect 24118 21904 24124 21916
rect 24176 21904 24182 21956
rect 24228 21944 24256 21984
rect 24394 21972 24400 21984
rect 24452 21972 24458 22024
rect 24504 22021 24532 22052
rect 30558 22040 30564 22052
rect 30616 22080 30622 22092
rect 30834 22080 30840 22092
rect 30616 22052 30840 22080
rect 30616 22040 30622 22052
rect 30834 22040 30840 22052
rect 30892 22040 30898 22092
rect 36814 22080 36820 22092
rect 36775 22052 36820 22080
rect 36814 22040 36820 22052
rect 36872 22040 36878 22092
rect 38194 22040 38200 22092
rect 38252 22080 38258 22092
rect 38841 22083 38899 22089
rect 38841 22080 38853 22083
rect 38252 22052 38853 22080
rect 38252 22040 38258 22052
rect 38841 22049 38853 22052
rect 38887 22049 38899 22083
rect 38841 22043 38899 22049
rect 40773 22083 40831 22089
rect 40773 22049 40785 22083
rect 40819 22080 40831 22083
rect 42536 22080 42564 22176
rect 56965 22151 57023 22157
rect 56965 22117 56977 22151
rect 57011 22148 57023 22151
rect 57011 22120 57045 22148
rect 57011 22117 57023 22120
rect 56965 22111 57023 22117
rect 56980 22080 57008 22111
rect 57054 22080 57060 22092
rect 40819 22052 42564 22080
rect 46492 22052 46888 22080
rect 56980 22052 57060 22080
rect 40819 22049 40831 22052
rect 40773 22043 40831 22049
rect 46492 22024 46520 22052
rect 24489 22015 24547 22021
rect 24489 21981 24501 22015
rect 24535 21981 24547 22015
rect 24489 21975 24547 21981
rect 24673 22015 24731 22021
rect 24673 21981 24685 22015
rect 24719 21981 24731 22015
rect 24673 21975 24731 21981
rect 24688 21944 24716 21975
rect 24762 21972 24768 22024
rect 24820 22012 24826 22024
rect 25685 22015 25743 22021
rect 24820 21984 24865 22012
rect 24820 21972 24826 21984
rect 25685 21981 25697 22015
rect 25731 21981 25743 22015
rect 25685 21975 25743 21981
rect 34149 22015 34207 22021
rect 34149 21981 34161 22015
rect 34195 22012 34207 22015
rect 34514 22012 34520 22024
rect 34195 21984 34520 22012
rect 34195 21981 34207 21984
rect 34149 21975 34207 21981
rect 25700 21944 25728 21975
rect 34514 21972 34520 21984
rect 34572 22012 34578 22024
rect 34701 22015 34759 22021
rect 34701 22012 34713 22015
rect 34572 21984 34713 22012
rect 34572 21972 34578 21984
rect 34701 21981 34713 21984
rect 34747 21981 34759 22015
rect 34701 21975 34759 21981
rect 36909 22015 36967 22021
rect 36909 21981 36921 22015
rect 36955 22012 36967 22015
rect 37274 22012 37280 22024
rect 36955 21984 37280 22012
rect 36955 21981 36967 21984
rect 36909 21975 36967 21981
rect 37274 21972 37280 21984
rect 37332 21972 37338 22024
rect 38930 22012 38936 22024
rect 38891 21984 38936 22012
rect 38930 21972 38936 21984
rect 38988 21972 38994 22024
rect 39022 21972 39028 22024
rect 39080 22012 39086 22024
rect 42797 22015 42855 22021
rect 42797 22012 42809 22015
rect 39080 21984 42809 22012
rect 39080 21972 39086 21984
rect 42797 21981 42809 21984
rect 42843 22012 42855 22015
rect 42886 22012 42892 22024
rect 42843 21984 42892 22012
rect 42843 21981 42855 21984
rect 42797 21975 42855 21981
rect 42886 21972 42892 21984
rect 42944 21972 42950 22024
rect 42978 21972 42984 22024
rect 43036 22012 43042 22024
rect 45646 22012 45652 22024
rect 43036 21984 43081 22012
rect 45607 21984 45652 22012
rect 43036 21972 43042 21984
rect 45646 21972 45652 21984
rect 45704 21972 45710 22024
rect 45925 22015 45983 22021
rect 45925 21981 45937 22015
rect 45971 22012 45983 22015
rect 46474 22012 46480 22024
rect 45971 21984 46480 22012
rect 45971 21981 45983 21984
rect 45925 21975 45983 21981
rect 46474 21972 46480 21984
rect 46532 21972 46538 22024
rect 46860 22021 46888 22052
rect 57054 22040 57060 22052
rect 57112 22040 57118 22092
rect 46569 22015 46627 22021
rect 46569 21981 46581 22015
rect 46615 22012 46627 22015
rect 46845 22015 46903 22021
rect 46615 21984 46796 22012
rect 46615 21981 46627 21984
rect 46569 21975 46627 21981
rect 26145 21947 26203 21953
rect 26145 21944 26157 21947
rect 24228 21916 26157 21944
rect 26145 21913 26157 21916
rect 26191 21913 26203 21947
rect 26145 21907 26203 21913
rect 26620 21916 29868 21944
rect 22971 21848 23520 21876
rect 22971 21845 22983 21848
rect 22925 21839 22983 21845
rect 23566 21836 23572 21888
rect 23624 21876 23630 21888
rect 23677 21879 23735 21885
rect 23677 21876 23689 21879
rect 23624 21848 23689 21876
rect 23624 21836 23630 21848
rect 23677 21845 23689 21848
rect 23723 21845 23735 21879
rect 23677 21839 23735 21845
rect 25314 21836 25320 21888
rect 25372 21876 25378 21888
rect 25501 21879 25559 21885
rect 25501 21876 25513 21879
rect 25372 21848 25513 21876
rect 25372 21836 25378 21848
rect 25501 21845 25513 21848
rect 25547 21876 25559 21879
rect 26620 21876 26648 21916
rect 29840 21888 29868 21916
rect 32674 21904 32680 21956
rect 32732 21944 32738 21956
rect 40310 21944 40316 21956
rect 32732 21916 40316 21944
rect 32732 21904 32738 21916
rect 40310 21904 40316 21916
rect 40368 21904 40374 21956
rect 45664 21944 45692 21972
rect 46661 21947 46719 21953
rect 46661 21944 46673 21947
rect 45664 21916 46673 21944
rect 46661 21913 46673 21916
rect 46707 21913 46719 21947
rect 46661 21907 46719 21913
rect 26786 21876 26792 21888
rect 25547 21848 26648 21876
rect 26747 21848 26792 21876
rect 25547 21845 25559 21848
rect 25501 21839 25559 21845
rect 26786 21836 26792 21848
rect 26844 21836 26850 21888
rect 29822 21836 29828 21888
rect 29880 21876 29886 21888
rect 33042 21876 33048 21888
rect 29880 21848 33048 21876
rect 29880 21836 29886 21848
rect 33042 21836 33048 21848
rect 33100 21836 33106 21888
rect 33318 21876 33324 21888
rect 33279 21848 33324 21876
rect 33318 21836 33324 21848
rect 33376 21836 33382 21888
rect 34698 21836 34704 21888
rect 34756 21876 34762 21888
rect 35437 21879 35495 21885
rect 35437 21876 35449 21879
rect 34756 21848 35449 21876
rect 34756 21836 34762 21848
rect 35437 21845 35449 21848
rect 35483 21845 35495 21879
rect 38194 21876 38200 21888
rect 38155 21848 38200 21876
rect 35437 21839 35495 21845
rect 38194 21836 38200 21848
rect 38252 21836 38258 21888
rect 45741 21879 45799 21885
rect 45741 21845 45753 21879
rect 45787 21876 45799 21879
rect 45830 21876 45836 21888
rect 45787 21848 45836 21876
rect 45787 21845 45799 21848
rect 45741 21839 45799 21845
rect 45830 21836 45836 21848
rect 45888 21876 45894 21888
rect 46768 21876 46796 21984
rect 46845 21981 46857 22015
rect 46891 21981 46903 22015
rect 46845 21975 46903 21981
rect 56689 22015 56747 22021
rect 56689 21981 56701 22015
rect 56735 21981 56747 22015
rect 56689 21975 56747 21981
rect 56965 22015 57023 22021
rect 56965 21981 56977 22015
rect 57011 22012 57023 22015
rect 57146 22012 57152 22024
rect 57011 21984 57152 22012
rect 57011 21981 57023 21984
rect 56965 21975 57023 21981
rect 56704 21944 56732 21975
rect 57146 21972 57152 21984
rect 57204 21972 57210 22024
rect 57974 21944 57980 21956
rect 56704 21916 57980 21944
rect 57974 21904 57980 21916
rect 58032 21904 58038 21956
rect 45888 21848 46796 21876
rect 45888 21836 45894 21848
rect 55674 21836 55680 21888
rect 55732 21876 55738 21888
rect 56781 21879 56839 21885
rect 56781 21876 56793 21879
rect 55732 21848 56793 21876
rect 55732 21836 55738 21848
rect 56781 21845 56793 21848
rect 56827 21845 56839 21879
rect 56781 21839 56839 21845
rect 1104 21786 58880 21808
rect 1104 21734 19574 21786
rect 19626 21734 19638 21786
rect 19690 21734 19702 21786
rect 19754 21734 19766 21786
rect 19818 21734 19830 21786
rect 19882 21734 50294 21786
rect 50346 21734 50358 21786
rect 50410 21734 50422 21786
rect 50474 21734 50486 21786
rect 50538 21734 50550 21786
rect 50602 21734 58880 21786
rect 1104 21712 58880 21734
rect 2225 21675 2283 21681
rect 2225 21641 2237 21675
rect 2271 21672 2283 21675
rect 2866 21672 2872 21684
rect 2271 21644 2872 21672
rect 2271 21641 2283 21644
rect 2225 21635 2283 21641
rect 2866 21632 2872 21644
rect 2924 21672 2930 21684
rect 2924 21644 3096 21672
rect 2924 21632 2930 21644
rect 2240 21576 2774 21604
rect 2240 21548 2268 21576
rect 1394 21536 1400 21548
rect 1355 21508 1400 21536
rect 1394 21496 1400 21508
rect 1452 21496 1458 21548
rect 2133 21539 2191 21545
rect 2133 21505 2145 21539
rect 2179 21536 2191 21539
rect 2222 21536 2228 21548
rect 2179 21508 2228 21536
rect 2179 21505 2191 21508
rect 2133 21499 2191 21505
rect 2222 21496 2228 21508
rect 2280 21496 2286 21548
rect 2746 21536 2774 21576
rect 2961 21539 3019 21545
rect 2961 21536 2973 21539
rect 2746 21508 2973 21536
rect 2961 21505 2973 21508
rect 3007 21505 3019 21539
rect 2961 21499 3019 21505
rect 2774 21428 2780 21480
rect 2832 21468 2838 21480
rect 2832 21440 2877 21468
rect 2832 21428 2838 21440
rect 3068 21400 3096 21644
rect 4614 21632 4620 21684
rect 4672 21672 4678 21684
rect 5166 21672 5172 21684
rect 4672 21644 5172 21672
rect 4672 21632 4678 21644
rect 5166 21632 5172 21644
rect 5224 21632 5230 21684
rect 9591 21675 9649 21681
rect 9591 21641 9603 21675
rect 9637 21672 9649 21675
rect 9950 21672 9956 21684
rect 9637 21644 9956 21672
rect 9637 21641 9649 21644
rect 9591 21635 9649 21641
rect 9950 21632 9956 21644
rect 10008 21632 10014 21684
rect 11514 21672 11520 21684
rect 10428 21644 11520 21672
rect 3145 21607 3203 21613
rect 3145 21573 3157 21607
rect 3191 21604 3203 21607
rect 5074 21604 5080 21616
rect 3191 21576 5080 21604
rect 3191 21573 3203 21576
rect 3145 21567 3203 21573
rect 5074 21564 5080 21576
rect 5132 21564 5138 21616
rect 9490 21604 9496 21616
rect 4154 21536 4160 21548
rect 4115 21508 4160 21536
rect 4154 21496 4160 21508
rect 4212 21496 4218 21548
rect 4614 21536 4620 21548
rect 4575 21508 4620 21536
rect 4614 21496 4620 21508
rect 4672 21496 4678 21548
rect 6730 21496 6736 21548
rect 6788 21536 6794 21548
rect 7101 21539 7159 21545
rect 7101 21536 7113 21539
rect 6788 21508 7113 21536
rect 6788 21496 6794 21508
rect 7101 21505 7113 21508
rect 7147 21505 7159 21539
rect 7101 21499 7159 21505
rect 7558 21496 7564 21548
rect 7616 21536 7622 21548
rect 7653 21539 7711 21545
rect 7653 21536 7665 21539
rect 7616 21508 7665 21536
rect 7616 21496 7622 21508
rect 7653 21505 7665 21508
rect 7699 21505 7711 21539
rect 7653 21499 7711 21505
rect 8588 21468 8616 21590
rect 9451 21576 9496 21604
rect 9490 21564 9496 21576
rect 9548 21564 9554 21616
rect 9674 21604 9680 21616
rect 9635 21576 9680 21604
rect 9674 21564 9680 21576
rect 9732 21604 9738 21616
rect 10428 21604 10456 21644
rect 11514 21632 11520 21644
rect 11572 21632 11578 21684
rect 13538 21672 13544 21684
rect 13499 21644 13544 21672
rect 13538 21632 13544 21644
rect 13596 21632 13602 21684
rect 15930 21632 15936 21684
rect 15988 21672 15994 21684
rect 16025 21675 16083 21681
rect 16025 21672 16037 21675
rect 15988 21644 16037 21672
rect 15988 21632 15994 21644
rect 16025 21641 16037 21644
rect 16071 21672 16083 21675
rect 16482 21672 16488 21684
rect 16071 21644 16488 21672
rect 16071 21641 16083 21644
rect 16025 21635 16083 21641
rect 16482 21632 16488 21644
rect 16540 21632 16546 21684
rect 19705 21675 19763 21681
rect 19705 21641 19717 21675
rect 19751 21672 19763 21675
rect 20070 21672 20076 21684
rect 19751 21644 20076 21672
rect 19751 21641 19763 21644
rect 19705 21635 19763 21641
rect 20070 21632 20076 21644
rect 20128 21632 20134 21684
rect 20530 21672 20536 21684
rect 20180 21644 20536 21672
rect 14182 21604 14188 21616
rect 9732 21576 10456 21604
rect 12820 21576 14188 21604
rect 9732 21564 9738 21576
rect 9766 21536 9772 21548
rect 9727 21508 9772 21536
rect 9766 21496 9772 21508
rect 9824 21496 9830 21548
rect 9858 21496 9864 21548
rect 9916 21536 9922 21548
rect 10321 21539 10379 21545
rect 10321 21536 10333 21539
rect 9916 21508 10333 21536
rect 9916 21496 9922 21508
rect 10321 21505 10333 21508
rect 10367 21505 10379 21539
rect 10321 21499 10379 21505
rect 10505 21539 10563 21545
rect 10505 21505 10517 21539
rect 10551 21536 10563 21539
rect 12820 21536 12848 21576
rect 14182 21564 14188 21576
rect 14240 21564 14246 21616
rect 17129 21607 17187 21613
rect 17129 21573 17141 21607
rect 17175 21604 17187 21607
rect 17586 21604 17592 21616
rect 17175 21576 17592 21604
rect 17175 21573 17187 21576
rect 17129 21567 17187 21573
rect 17586 21564 17592 21576
rect 17644 21564 17650 21616
rect 18690 21564 18696 21616
rect 18748 21604 18754 21616
rect 19429 21607 19487 21613
rect 18748 21576 19196 21604
rect 18748 21564 18754 21576
rect 10551 21508 12848 21536
rect 10551 21505 10563 21508
rect 10505 21499 10563 21505
rect 12894 21496 12900 21548
rect 12952 21536 12958 21548
rect 12989 21539 13047 21545
rect 12989 21536 13001 21539
rect 12952 21508 13001 21536
rect 12952 21496 12958 21508
rect 12989 21505 13001 21508
rect 13035 21505 13047 21539
rect 13170 21536 13176 21548
rect 13131 21508 13176 21536
rect 12989 21499 13047 21505
rect 13170 21496 13176 21508
rect 13228 21496 13234 21548
rect 13265 21539 13323 21545
rect 13265 21505 13277 21539
rect 13311 21505 13323 21539
rect 13265 21499 13323 21505
rect 11054 21468 11060 21480
rect 8588 21440 11060 21468
rect 11054 21428 11060 21440
rect 11112 21428 11118 21480
rect 11238 21428 11244 21480
rect 11296 21468 11302 21480
rect 13280 21468 13308 21499
rect 13354 21496 13360 21548
rect 13412 21536 13418 21548
rect 14369 21539 14427 21545
rect 13412 21508 13457 21536
rect 13412 21496 13418 21508
rect 14369 21505 14381 21539
rect 14415 21536 14427 21539
rect 14918 21536 14924 21548
rect 14415 21508 14924 21536
rect 14415 21505 14427 21508
rect 14369 21499 14427 21505
rect 14918 21496 14924 21508
rect 14976 21496 14982 21548
rect 19058 21536 19064 21548
rect 19019 21508 19064 21536
rect 19058 21496 19064 21508
rect 19116 21496 19122 21548
rect 19168 21545 19196 21576
rect 19429 21573 19441 21607
rect 19475 21604 19487 21607
rect 19978 21604 19984 21616
rect 19475 21576 19984 21604
rect 19475 21573 19487 21576
rect 19429 21567 19487 21573
rect 19978 21564 19984 21576
rect 20036 21604 20042 21616
rect 20180 21604 20208 21644
rect 20530 21632 20536 21644
rect 20588 21632 20594 21684
rect 20898 21632 20904 21684
rect 20956 21672 20962 21684
rect 21542 21672 21548 21684
rect 20956 21644 21548 21672
rect 20956 21632 20962 21644
rect 21542 21632 21548 21644
rect 21600 21632 21606 21684
rect 23106 21672 23112 21684
rect 23067 21644 23112 21672
rect 23106 21632 23112 21644
rect 23164 21632 23170 21684
rect 23658 21672 23664 21684
rect 23619 21644 23664 21672
rect 23658 21632 23664 21644
rect 23716 21632 23722 21684
rect 25590 21672 25596 21684
rect 24136 21644 25268 21672
rect 25551 21644 25596 21672
rect 20346 21604 20352 21616
rect 20036 21576 20208 21604
rect 20307 21576 20352 21604
rect 20036 21564 20042 21576
rect 20346 21564 20352 21576
rect 20404 21564 20410 21616
rect 21082 21564 21088 21616
rect 21140 21604 21146 21616
rect 23124 21604 23152 21632
rect 24136 21604 24164 21644
rect 21140 21576 23060 21604
rect 23124 21576 24164 21604
rect 21140 21564 21146 21576
rect 19610 21545 19616 21548
rect 19154 21539 19212 21545
rect 19154 21505 19166 21539
rect 19200 21505 19212 21539
rect 19154 21499 19212 21505
rect 19337 21539 19395 21545
rect 19337 21505 19349 21539
rect 19383 21505 19395 21539
rect 19337 21499 19395 21505
rect 19567 21539 19616 21545
rect 19567 21505 19579 21539
rect 19613 21505 19616 21539
rect 19567 21499 19616 21505
rect 11296 21440 12940 21468
rect 11296 21428 11302 21440
rect 8018 21400 8024 21412
rect 3068 21372 8024 21400
rect 8018 21360 8024 21372
rect 8076 21360 8082 21412
rect 1578 21332 1584 21344
rect 1539 21304 1584 21332
rect 1578 21292 1584 21304
rect 1636 21292 1642 21344
rect 5810 21332 5816 21344
rect 5771 21304 5816 21332
rect 5810 21292 5816 21304
rect 5868 21292 5874 21344
rect 12912 21332 12940 21440
rect 13004 21440 13308 21468
rect 13004 21412 13032 21440
rect 18046 21428 18052 21480
rect 18104 21468 18110 21480
rect 19352 21468 19380 21499
rect 19610 21496 19616 21499
rect 19668 21496 19674 21548
rect 22830 21536 22836 21548
rect 19725 21508 22836 21536
rect 18104 21440 19380 21468
rect 18104 21428 18110 21440
rect 12986 21360 12992 21412
rect 13044 21360 13050 21412
rect 19725 21400 19753 21508
rect 22830 21496 22836 21508
rect 22888 21496 22894 21548
rect 23032 21536 23060 21576
rect 24210 21564 24216 21616
rect 24268 21604 24274 21616
rect 24413 21607 24471 21613
rect 24413 21604 24425 21607
rect 24268 21576 24313 21604
rect 24268 21564 24274 21576
rect 24412 21573 24425 21604
rect 24459 21573 24471 21607
rect 25240 21604 25268 21644
rect 25590 21632 25596 21644
rect 25648 21632 25654 21684
rect 31570 21672 31576 21684
rect 31531 21644 31576 21672
rect 31570 21632 31576 21644
rect 31628 21632 31634 21684
rect 31662 21632 31668 21684
rect 31720 21672 31726 21684
rect 32674 21672 32680 21684
rect 31720 21644 32680 21672
rect 31720 21632 31726 21644
rect 32674 21632 32680 21644
rect 32732 21632 32738 21684
rect 32769 21675 32827 21681
rect 32769 21641 32781 21675
rect 32815 21672 32827 21675
rect 32950 21672 32956 21684
rect 32815 21644 32956 21672
rect 32815 21641 32827 21644
rect 32769 21635 32827 21641
rect 32950 21632 32956 21644
rect 33008 21632 33014 21684
rect 34425 21675 34483 21681
rect 34425 21641 34437 21675
rect 34471 21672 34483 21675
rect 34514 21672 34520 21684
rect 34471 21644 34520 21672
rect 34471 21641 34483 21644
rect 34425 21635 34483 21641
rect 34514 21632 34520 21644
rect 34572 21632 34578 21684
rect 34606 21632 34612 21684
rect 34664 21672 34670 21684
rect 39022 21672 39028 21684
rect 34664 21644 39028 21672
rect 34664 21632 34670 21644
rect 39022 21632 39028 21644
rect 39080 21632 39086 21684
rect 46385 21675 46443 21681
rect 46385 21641 46397 21675
rect 46431 21672 46443 21675
rect 49053 21675 49111 21681
rect 46431 21644 48452 21672
rect 46431 21641 46443 21644
rect 46385 21635 46443 21641
rect 26237 21607 26295 21613
rect 26237 21604 26249 21607
rect 25240 21576 26249 21604
rect 24412 21567 24471 21573
rect 26237 21573 26249 21576
rect 26283 21604 26295 21607
rect 26786 21604 26792 21616
rect 26283 21576 26792 21604
rect 26283 21573 26295 21576
rect 26237 21567 26295 21573
rect 24302 21536 24308 21548
rect 23032 21508 24308 21536
rect 24302 21496 24308 21508
rect 24360 21496 24366 21548
rect 24412 21468 24440 21567
rect 26786 21564 26792 21576
rect 26844 21564 26850 21616
rect 27982 21564 27988 21616
rect 28040 21604 28046 21616
rect 32968 21604 32996 21632
rect 28040 21576 32996 21604
rect 28040 21564 28046 21576
rect 25038 21536 25044 21548
rect 24999 21508 25044 21536
rect 25038 21496 25044 21508
rect 25096 21496 25102 21548
rect 25130 21496 25136 21548
rect 25188 21536 25194 21548
rect 25314 21536 25320 21548
rect 25188 21508 25233 21536
rect 25275 21508 25320 21536
rect 25188 21496 25194 21508
rect 25314 21496 25320 21508
rect 25372 21496 25378 21548
rect 25406 21496 25412 21548
rect 25464 21536 25470 21548
rect 25464 21508 25509 21536
rect 25464 21496 25470 21508
rect 26326 21496 26332 21548
rect 26384 21536 26390 21548
rect 27433 21539 27491 21545
rect 27433 21536 27445 21539
rect 26384 21508 27445 21536
rect 26384 21496 26390 21508
rect 27433 21505 27445 21508
rect 27479 21505 27491 21539
rect 27433 21499 27491 21505
rect 27617 21539 27675 21545
rect 27617 21505 27629 21539
rect 27663 21536 27675 21539
rect 27798 21536 27804 21548
rect 27663 21508 27804 21536
rect 27663 21505 27675 21508
rect 27617 21499 27675 21505
rect 27798 21496 27804 21508
rect 27856 21496 27862 21548
rect 30558 21536 30564 21548
rect 30519 21508 30564 21536
rect 30558 21496 30564 21508
rect 30616 21496 30622 21548
rect 30929 21539 30987 21545
rect 30929 21505 30941 21539
rect 30975 21536 30987 21539
rect 32968 21536 32996 21576
rect 35342 21564 35348 21616
rect 35400 21604 35406 21616
rect 45002 21604 45008 21616
rect 35400 21576 45008 21604
rect 35400 21564 35406 21576
rect 45002 21564 45008 21576
rect 45060 21564 45066 21616
rect 48424 21548 48452 21644
rect 49053 21641 49065 21675
rect 49099 21672 49111 21675
rect 49326 21672 49332 21684
rect 49099 21644 49332 21672
rect 49099 21641 49111 21644
rect 49053 21635 49111 21641
rect 49326 21632 49332 21644
rect 49384 21632 49390 21684
rect 52181 21675 52239 21681
rect 52181 21641 52193 21675
rect 52227 21672 52239 21675
rect 53006 21672 53012 21684
rect 52227 21644 53012 21672
rect 52227 21641 52239 21644
rect 52181 21635 52239 21641
rect 53006 21632 53012 21644
rect 53064 21632 53070 21684
rect 53282 21672 53288 21684
rect 53243 21644 53288 21672
rect 53282 21632 53288 21644
rect 53340 21632 53346 21684
rect 54389 21675 54447 21681
rect 54389 21641 54401 21675
rect 54435 21672 54447 21675
rect 54478 21672 54484 21684
rect 54435 21644 54484 21672
rect 54435 21641 54447 21644
rect 54389 21635 54447 21641
rect 54478 21632 54484 21644
rect 54536 21632 54542 21684
rect 56505 21675 56563 21681
rect 56505 21641 56517 21675
rect 56551 21672 56563 21675
rect 56686 21672 56692 21684
rect 56551 21644 56692 21672
rect 56551 21641 56563 21644
rect 56505 21635 56563 21641
rect 56686 21632 56692 21644
rect 56744 21632 56750 21684
rect 57057 21675 57115 21681
rect 57057 21641 57069 21675
rect 57103 21672 57115 21675
rect 57146 21672 57152 21684
rect 57103 21644 57152 21672
rect 57103 21641 57115 21644
rect 57057 21635 57115 21641
rect 57146 21632 57152 21644
rect 57204 21632 57210 21684
rect 57974 21672 57980 21684
rect 57935 21644 57980 21672
rect 57974 21632 57980 21644
rect 58032 21632 58038 21684
rect 49344 21604 49372 21632
rect 53300 21604 53328 21632
rect 53742 21604 53748 21616
rect 49344 21576 49924 21604
rect 33229 21539 33287 21545
rect 33229 21536 33241 21539
rect 30975 21508 31754 21536
rect 32968 21508 33241 21536
rect 30975 21505 30987 21508
rect 30929 21499 30987 21505
rect 25682 21468 25688 21480
rect 13096 21372 19753 21400
rect 19812 21440 25688 21468
rect 13096 21332 13124 21372
rect 12912 21304 13124 21332
rect 14185 21335 14243 21341
rect 14185 21301 14197 21335
rect 14231 21332 14243 21335
rect 16298 21332 16304 21344
rect 14231 21304 16304 21332
rect 14231 21301 14243 21304
rect 14185 21295 14243 21301
rect 16298 21292 16304 21304
rect 16356 21292 16362 21344
rect 17218 21332 17224 21344
rect 17179 21304 17224 21332
rect 17218 21292 17224 21304
rect 17276 21292 17282 21344
rect 18414 21292 18420 21344
rect 18472 21332 18478 21344
rect 18509 21335 18567 21341
rect 18509 21332 18521 21335
rect 18472 21304 18521 21332
rect 18472 21292 18478 21304
rect 18509 21301 18521 21304
rect 18555 21301 18567 21335
rect 18509 21295 18567 21301
rect 18598 21292 18604 21344
rect 18656 21332 18662 21344
rect 19812 21332 19840 21440
rect 25682 21428 25688 21440
rect 25740 21428 25746 21480
rect 31726 21468 31754 21508
rect 33229 21505 33241 21508
rect 33275 21505 33287 21539
rect 33229 21499 33287 21505
rect 34790 21496 34796 21548
rect 34848 21536 34854 21548
rect 35437 21539 35495 21545
rect 35437 21536 35449 21539
rect 34848 21508 35449 21536
rect 34848 21496 34854 21508
rect 35437 21505 35449 21508
rect 35483 21505 35495 21539
rect 35437 21499 35495 21505
rect 45646 21496 45652 21548
rect 45704 21536 45710 21548
rect 46385 21539 46443 21545
rect 46385 21536 46397 21539
rect 45704 21508 46397 21536
rect 45704 21496 45710 21508
rect 46385 21505 46397 21508
rect 46431 21505 46443 21539
rect 48406 21536 48412 21548
rect 48319 21508 48412 21536
rect 46385 21499 46443 21505
rect 48406 21496 48412 21508
rect 48464 21496 48470 21548
rect 49694 21536 49700 21548
rect 49655 21508 49700 21536
rect 49694 21496 49700 21508
rect 49752 21496 49758 21548
rect 49896 21545 49924 21576
rect 51736 21576 53052 21604
rect 53300 21576 53748 21604
rect 49881 21539 49939 21545
rect 49881 21505 49893 21539
rect 49927 21505 49939 21539
rect 49881 21499 49939 21505
rect 51736 21480 51764 21576
rect 53024 21545 53052 21576
rect 53742 21564 53748 21576
rect 53800 21604 53806 21616
rect 53800 21576 53880 21604
rect 53800 21564 53806 21576
rect 53852 21545 53880 21576
rect 56336 21576 57192 21604
rect 51997 21539 52055 21545
rect 51997 21505 52009 21539
rect 52043 21536 52055 21539
rect 52733 21539 52791 21545
rect 52733 21536 52745 21539
rect 52043 21508 52745 21536
rect 52043 21505 52055 21508
rect 51997 21499 52055 21505
rect 52733 21505 52745 21508
rect 52779 21505 52791 21539
rect 52733 21499 52791 21505
rect 53009 21539 53067 21545
rect 53009 21505 53021 21539
rect 53055 21536 53067 21539
rect 53837 21539 53895 21545
rect 53055 21508 53328 21536
rect 53055 21505 53067 21508
rect 53009 21499 53067 21505
rect 33321 21471 33379 21477
rect 33321 21468 33333 21471
rect 31726 21440 33333 21468
rect 33321 21437 33333 21440
rect 33367 21468 33379 21471
rect 37274 21468 37280 21480
rect 33367 21440 37280 21468
rect 33367 21437 33379 21440
rect 33321 21431 33379 21437
rect 37274 21428 37280 21440
rect 37332 21428 37338 21480
rect 45830 21468 45836 21480
rect 45791 21440 45836 21468
rect 45830 21428 45836 21440
rect 45888 21428 45894 21480
rect 46474 21468 46480 21480
rect 46435 21440 46480 21468
rect 46474 21428 46480 21440
rect 46532 21428 46538 21480
rect 48314 21468 48320 21480
rect 48275 21440 48320 21468
rect 48314 21428 48320 21440
rect 48372 21428 48378 21480
rect 51718 21468 51724 21480
rect 51679 21440 51724 21468
rect 51718 21428 51724 21440
rect 51776 21428 51782 21480
rect 20346 21360 20352 21412
rect 20404 21400 20410 21412
rect 21450 21400 21456 21412
rect 20404 21372 21456 21400
rect 20404 21360 20410 21372
rect 21450 21360 21456 21372
rect 21508 21360 21514 21412
rect 21818 21360 21824 21412
rect 21876 21400 21882 21412
rect 26510 21400 26516 21412
rect 21876 21372 26516 21400
rect 21876 21360 21882 21372
rect 26510 21360 26516 21372
rect 26568 21360 26574 21412
rect 27525 21403 27583 21409
rect 27525 21369 27537 21403
rect 27571 21400 27583 21403
rect 36814 21400 36820 21412
rect 27571 21372 36820 21400
rect 27571 21369 27583 21372
rect 27525 21363 27583 21369
rect 36814 21360 36820 21372
rect 36872 21360 36878 21412
rect 49234 21360 49240 21412
rect 49292 21400 49298 21412
rect 52012 21400 52040 21499
rect 53193 21471 53251 21477
rect 53193 21437 53205 21471
rect 53239 21437 53251 21471
rect 53300 21468 53328 21508
rect 53837 21505 53849 21539
rect 53883 21505 53895 21539
rect 53837 21499 53895 21505
rect 53929 21539 53987 21545
rect 53929 21505 53941 21539
rect 53975 21505 53987 21539
rect 54110 21536 54116 21548
rect 54071 21508 54116 21536
rect 53929 21499 53987 21505
rect 53944 21468 53972 21499
rect 54110 21496 54116 21508
rect 54168 21496 54174 21548
rect 54202 21496 54208 21548
rect 54260 21536 54266 21548
rect 56336 21545 56364 21576
rect 56321 21539 56379 21545
rect 54260 21508 54305 21536
rect 54260 21496 54266 21508
rect 56321 21505 56333 21539
rect 56367 21505 56379 21539
rect 56962 21536 56968 21548
rect 56923 21508 56968 21536
rect 56321 21499 56379 21505
rect 56962 21496 56968 21508
rect 57020 21496 57026 21548
rect 57164 21545 57192 21576
rect 57149 21539 57207 21545
rect 57149 21505 57161 21539
rect 57195 21536 57207 21539
rect 57330 21536 57336 21548
rect 57195 21508 57336 21536
rect 57195 21505 57207 21508
rect 57149 21499 57207 21505
rect 57330 21496 57336 21508
rect 57388 21536 57394 21548
rect 57885 21539 57943 21545
rect 57885 21536 57897 21539
rect 57388 21508 57897 21536
rect 57388 21496 57394 21508
rect 57885 21505 57897 21508
rect 57931 21505 57943 21539
rect 57885 21499 57943 21505
rect 53300 21440 53972 21468
rect 53193 21431 53251 21437
rect 49292 21372 52040 21400
rect 49292 21360 49298 21372
rect 18656 21304 19840 21332
rect 20441 21335 20499 21341
rect 18656 21292 18662 21304
rect 20441 21301 20453 21335
rect 20487 21332 20499 21335
rect 20622 21332 20628 21344
rect 20487 21304 20628 21332
rect 20487 21301 20499 21304
rect 20441 21295 20499 21301
rect 20622 21292 20628 21304
rect 20680 21292 20686 21344
rect 20714 21292 20720 21344
rect 20772 21332 20778 21344
rect 21085 21335 21143 21341
rect 21085 21332 21097 21335
rect 20772 21304 21097 21332
rect 20772 21292 20778 21304
rect 21085 21301 21097 21304
rect 21131 21332 21143 21335
rect 22738 21332 22744 21344
rect 21131 21304 22744 21332
rect 21131 21301 21143 21304
rect 21085 21295 21143 21301
rect 22738 21292 22744 21304
rect 22796 21332 22802 21344
rect 23750 21332 23756 21344
rect 22796 21304 23756 21332
rect 22796 21292 22802 21304
rect 23750 21292 23756 21304
rect 23808 21292 23814 21344
rect 24302 21292 24308 21344
rect 24360 21332 24366 21344
rect 24397 21335 24455 21341
rect 24397 21332 24409 21335
rect 24360 21304 24409 21332
rect 24360 21292 24366 21304
rect 24397 21301 24409 21304
rect 24443 21301 24455 21335
rect 24397 21295 24455 21301
rect 24581 21335 24639 21341
rect 24581 21301 24593 21335
rect 24627 21332 24639 21335
rect 25130 21332 25136 21344
rect 24627 21304 25136 21332
rect 24627 21301 24639 21304
rect 24581 21295 24639 21301
rect 25130 21292 25136 21304
rect 25188 21292 25194 21344
rect 25958 21292 25964 21344
rect 26016 21332 26022 21344
rect 26145 21335 26203 21341
rect 26145 21332 26157 21335
rect 26016 21304 26157 21332
rect 26016 21292 26022 21304
rect 26145 21301 26157 21304
rect 26191 21332 26203 21335
rect 29086 21332 29092 21344
rect 26191 21304 29092 21332
rect 26191 21301 26203 21304
rect 26145 21295 26203 21301
rect 29086 21292 29092 21304
rect 29144 21292 29150 21344
rect 30009 21335 30067 21341
rect 30009 21301 30021 21335
rect 30055 21332 30067 21335
rect 30374 21332 30380 21344
rect 30055 21304 30380 21332
rect 30055 21301 30067 21304
rect 30009 21295 30067 21301
rect 30374 21292 30380 21304
rect 30432 21292 30438 21344
rect 35621 21335 35679 21341
rect 35621 21301 35633 21335
rect 35667 21332 35679 21335
rect 36998 21332 37004 21344
rect 35667 21304 37004 21332
rect 35667 21301 35679 21304
rect 35621 21295 35679 21301
rect 36998 21292 37004 21304
rect 37056 21292 37062 21344
rect 43346 21332 43352 21344
rect 43307 21304 43352 21332
rect 43346 21292 43352 21304
rect 43404 21292 43410 21344
rect 49789 21335 49847 21341
rect 49789 21301 49801 21335
rect 49835 21332 49847 21335
rect 51074 21332 51080 21344
rect 49835 21304 51080 21332
rect 49835 21301 49847 21304
rect 49789 21295 49847 21301
rect 51074 21292 51080 21304
rect 51132 21292 51138 21344
rect 51810 21332 51816 21344
rect 51723 21304 51816 21332
rect 51810 21292 51816 21304
rect 51868 21332 51874 21344
rect 53208 21332 53236 21431
rect 55674 21428 55680 21480
rect 55732 21468 55738 21480
rect 56137 21471 56195 21477
rect 56137 21468 56149 21471
rect 55732 21440 56149 21468
rect 55732 21428 55738 21440
rect 56137 21437 56149 21440
rect 56183 21437 56195 21471
rect 56137 21431 56195 21437
rect 51868 21304 53236 21332
rect 51868 21292 51874 21304
rect 1104 21242 58880 21264
rect 1104 21190 4214 21242
rect 4266 21190 4278 21242
rect 4330 21190 4342 21242
rect 4394 21190 4406 21242
rect 4458 21190 4470 21242
rect 4522 21190 34934 21242
rect 34986 21190 34998 21242
rect 35050 21190 35062 21242
rect 35114 21190 35126 21242
rect 35178 21190 35190 21242
rect 35242 21190 58880 21242
rect 1104 21168 58880 21190
rect 1394 21128 1400 21140
rect 1355 21100 1400 21128
rect 1394 21088 1400 21100
rect 1452 21088 1458 21140
rect 3142 21088 3148 21140
rect 3200 21128 3206 21140
rect 4341 21131 4399 21137
rect 4341 21128 4353 21131
rect 3200 21100 4353 21128
rect 3200 21088 3206 21100
rect 4341 21097 4353 21100
rect 4387 21097 4399 21131
rect 9490 21128 9496 21140
rect 9451 21100 9496 21128
rect 4341 21091 4399 21097
rect 9490 21088 9496 21100
rect 9548 21088 9554 21140
rect 9766 21088 9772 21140
rect 9824 21128 9830 21140
rect 10137 21131 10195 21137
rect 10137 21128 10149 21131
rect 9824 21100 10149 21128
rect 9824 21088 9830 21100
rect 10137 21097 10149 21100
rect 10183 21097 10195 21131
rect 10137 21091 10195 21097
rect 13354 21088 13360 21140
rect 13412 21128 13418 21140
rect 14093 21131 14151 21137
rect 14093 21128 14105 21131
rect 13412 21100 14105 21128
rect 13412 21088 13418 21100
rect 14093 21097 14105 21100
rect 14139 21128 14151 21131
rect 14642 21128 14648 21140
rect 14139 21100 14648 21128
rect 14139 21097 14151 21100
rect 14093 21091 14151 21097
rect 14642 21088 14648 21100
rect 14700 21088 14706 21140
rect 14826 21088 14832 21140
rect 14884 21128 14890 21140
rect 14884 21100 19661 21128
rect 14884 21088 14890 21100
rect 5810 21020 5816 21072
rect 5868 21060 5874 21072
rect 14550 21060 14556 21072
rect 5868 21032 14556 21060
rect 5868 21020 5874 21032
rect 14550 21020 14556 21032
rect 14608 21020 14614 21072
rect 15381 21063 15439 21069
rect 15381 21029 15393 21063
rect 15427 21029 15439 21063
rect 15381 21023 15439 21029
rect 2869 20995 2927 21001
rect 2869 20961 2881 20995
rect 2915 20992 2927 20995
rect 4614 20992 4620 21004
rect 2915 20964 4620 20992
rect 2915 20961 2927 20964
rect 2869 20955 2927 20961
rect 2498 20924 2504 20936
rect 2459 20896 2504 20924
rect 2498 20884 2504 20896
rect 2556 20884 2562 20936
rect 2682 20924 2688 20936
rect 2643 20896 2688 20924
rect 2682 20884 2688 20896
rect 2740 20884 2746 20936
rect 4264 20933 4292 20964
rect 4614 20952 4620 20964
rect 4672 20952 4678 21004
rect 5074 20992 5080 21004
rect 4724 20964 5080 20992
rect 4249 20927 4307 20933
rect 4249 20893 4261 20927
rect 4295 20893 4307 20927
rect 4249 20887 4307 20893
rect 4433 20927 4491 20933
rect 4433 20893 4445 20927
rect 4479 20924 4491 20927
rect 4724 20924 4752 20964
rect 5074 20952 5080 20964
rect 5132 20952 5138 21004
rect 6730 20992 6736 21004
rect 6691 20964 6736 20992
rect 6730 20952 6736 20964
rect 6788 20952 6794 21004
rect 7101 20995 7159 21001
rect 7101 20961 7113 20995
rect 7147 20992 7159 20995
rect 7466 20992 7472 21004
rect 7147 20964 7472 20992
rect 7147 20961 7159 20964
rect 7101 20955 7159 20961
rect 7466 20952 7472 20964
rect 7524 20952 7530 21004
rect 13814 20952 13820 21004
rect 13872 20992 13878 21004
rect 13872 20964 15332 20992
rect 13872 20952 13878 20964
rect 4479 20896 4752 20924
rect 4801 20927 4859 20933
rect 4479 20893 4491 20896
rect 4433 20887 4491 20893
rect 4801 20893 4813 20927
rect 4847 20924 4859 20927
rect 4890 20924 4896 20936
rect 4847 20896 4896 20924
rect 4847 20893 4859 20896
rect 4801 20887 4859 20893
rect 4890 20884 4896 20896
rect 4948 20924 4954 20936
rect 6641 20927 6699 20933
rect 6641 20924 6653 20927
rect 4948 20896 6653 20924
rect 4948 20884 4954 20896
rect 6641 20893 6653 20896
rect 6687 20924 6699 20927
rect 7558 20924 7564 20936
rect 6687 20896 7564 20924
rect 6687 20893 6699 20896
rect 6641 20887 6699 20893
rect 7558 20884 7564 20896
rect 7616 20884 7622 20936
rect 8294 20884 8300 20936
rect 8352 20924 8358 20936
rect 9306 20924 9312 20936
rect 8352 20896 9312 20924
rect 8352 20884 8358 20896
rect 9306 20884 9312 20896
rect 9364 20924 9370 20936
rect 9953 20927 10011 20933
rect 9953 20924 9965 20927
rect 9364 20896 9965 20924
rect 9364 20884 9370 20896
rect 9953 20893 9965 20896
rect 9999 20893 10011 20927
rect 10778 20924 10784 20936
rect 10739 20896 10784 20924
rect 9953 20887 10011 20893
rect 10778 20884 10784 20896
rect 10836 20884 10842 20936
rect 13265 20927 13323 20933
rect 13265 20893 13277 20927
rect 13311 20924 13323 20927
rect 13722 20924 13728 20936
rect 13311 20896 13728 20924
rect 13311 20893 13323 20896
rect 13265 20887 13323 20893
rect 13722 20884 13728 20896
rect 13780 20924 13786 20936
rect 14826 20924 14832 20936
rect 13780 20896 14832 20924
rect 13780 20884 13786 20896
rect 14826 20884 14832 20896
rect 14884 20884 14890 20936
rect 14918 20884 14924 20936
rect 14976 20924 14982 20936
rect 15197 20927 15255 20933
rect 15197 20924 15209 20927
rect 14976 20896 15209 20924
rect 14976 20884 14982 20896
rect 15197 20893 15209 20896
rect 15243 20893 15255 20927
rect 15197 20887 15255 20893
rect 7834 20856 7840 20868
rect 4632 20828 7840 20856
rect 4632 20797 4660 20828
rect 7834 20816 7840 20828
rect 7892 20816 7898 20868
rect 8110 20816 8116 20868
rect 8168 20856 8174 20868
rect 10796 20856 10824 20884
rect 8168 20828 10824 20856
rect 8168 20816 8174 20828
rect 12986 20816 12992 20868
rect 13044 20856 13050 20868
rect 13081 20859 13139 20865
rect 13081 20856 13093 20859
rect 13044 20828 13093 20856
rect 13044 20816 13050 20828
rect 13081 20825 13093 20828
rect 13127 20825 13139 20859
rect 13081 20819 13139 20825
rect 13170 20816 13176 20868
rect 13228 20856 13234 20868
rect 15010 20856 15016 20868
rect 13228 20828 15016 20856
rect 13228 20816 13234 20828
rect 15010 20816 15016 20828
rect 15068 20816 15074 20868
rect 15105 20859 15163 20865
rect 15105 20825 15117 20859
rect 15151 20825 15163 20859
rect 15304 20856 15332 20964
rect 15396 20924 15424 21023
rect 16114 21020 16120 21072
rect 16172 21060 16178 21072
rect 17037 21063 17095 21069
rect 17037 21060 17049 21063
rect 16172 21032 17049 21060
rect 16172 21020 16178 21032
rect 17037 21029 17049 21032
rect 17083 21029 17095 21063
rect 17037 21023 17095 21029
rect 17218 21020 17224 21072
rect 17276 21060 17282 21072
rect 19518 21060 19524 21072
rect 17276 21032 19524 21060
rect 17276 21020 17282 21032
rect 19518 21020 19524 21032
rect 19576 21020 19582 21072
rect 17236 20992 17264 21020
rect 18046 20992 18052 21004
rect 16224 20964 17264 20992
rect 18007 20964 18052 20992
rect 16224 20933 16252 20964
rect 18046 20952 18052 20964
rect 18104 20952 18110 21004
rect 18598 20992 18604 21004
rect 18156 20964 18604 20992
rect 15841 20927 15899 20933
rect 15841 20924 15853 20927
rect 15396 20896 15853 20924
rect 15841 20893 15853 20896
rect 15887 20893 15899 20927
rect 15841 20887 15899 20893
rect 15934 20927 15992 20933
rect 15934 20893 15946 20927
rect 15980 20893 15992 20927
rect 15934 20887 15992 20893
rect 16209 20927 16267 20933
rect 16209 20893 16221 20927
rect 16255 20893 16267 20927
rect 16209 20887 16267 20893
rect 15948 20856 15976 20887
rect 16298 20884 16304 20936
rect 16356 20933 16362 20936
rect 16356 20924 16364 20933
rect 18156 20924 18184 20964
rect 18598 20952 18604 20964
rect 18656 20952 18662 21004
rect 19633 20992 19661 21100
rect 19794 21088 19800 21140
rect 19852 21128 19858 21140
rect 24762 21128 24768 21140
rect 19852 21100 24768 21128
rect 19852 21088 19858 21100
rect 24762 21088 24768 21100
rect 24820 21088 24826 21140
rect 25038 21088 25044 21140
rect 25096 21128 25102 21140
rect 25961 21131 26019 21137
rect 25961 21128 25973 21131
rect 25096 21100 25973 21128
rect 25096 21088 25102 21100
rect 25961 21097 25973 21100
rect 26007 21097 26019 21131
rect 25961 21091 26019 21097
rect 27801 21131 27859 21137
rect 27801 21097 27813 21131
rect 27847 21128 27859 21131
rect 30742 21128 30748 21140
rect 27847 21100 30748 21128
rect 27847 21097 27859 21100
rect 27801 21091 27859 21097
rect 30742 21088 30748 21100
rect 30800 21088 30806 21140
rect 31662 21128 31668 21140
rect 30944 21100 31668 21128
rect 22189 21063 22247 21069
rect 20640 21032 22140 21060
rect 20640 20992 20668 21032
rect 21358 20992 21364 21004
rect 19633 20964 20668 20992
rect 20732 20964 21364 20992
rect 16356 20896 16401 20924
rect 16500 20896 18184 20924
rect 16356 20887 16364 20896
rect 16356 20884 16362 20887
rect 16114 20856 16120 20868
rect 15304 20828 15976 20856
rect 16075 20828 16120 20856
rect 15105 20819 15163 20825
rect 4617 20791 4675 20797
rect 4617 20757 4629 20791
rect 4663 20757 4675 20791
rect 6454 20788 6460 20800
rect 6415 20760 6460 20788
rect 4617 20751 4675 20757
rect 6454 20748 6460 20760
rect 6512 20748 6518 20800
rect 10873 20791 10931 20797
rect 10873 20757 10885 20791
rect 10919 20788 10931 20791
rect 15120 20788 15148 20819
rect 16114 20816 16120 20828
rect 16172 20816 16178 20868
rect 16500 20856 16528 20896
rect 18322 20884 18328 20936
rect 18380 20924 18386 20936
rect 19426 20933 19432 20936
rect 18417 20927 18475 20933
rect 18417 20924 18429 20927
rect 18380 20896 18429 20924
rect 18380 20884 18386 20896
rect 18417 20893 18429 20896
rect 18463 20893 18475 20927
rect 18417 20887 18475 20893
rect 18509 20927 18567 20933
rect 18509 20893 18521 20927
rect 18555 20893 18567 20927
rect 19245 20927 19303 20933
rect 19245 20924 19257 20927
rect 18509 20887 18567 20893
rect 18708 20896 19257 20924
rect 18138 20856 18144 20868
rect 16224 20828 16528 20856
rect 18099 20828 18144 20856
rect 16224 20788 16252 20828
rect 18138 20816 18144 20828
rect 18196 20816 18202 20868
rect 16482 20788 16488 20800
rect 10919 20760 16252 20788
rect 16443 20760 16488 20788
rect 10919 20757 10931 20760
rect 10873 20751 10931 20757
rect 16482 20748 16488 20760
rect 16540 20748 16546 20800
rect 18414 20748 18420 20800
rect 18472 20788 18478 20800
rect 18524 20788 18552 20887
rect 18708 20797 18736 20896
rect 19245 20893 19257 20896
rect 19291 20893 19303 20927
rect 19245 20887 19303 20893
rect 19393 20927 19432 20933
rect 19393 20893 19405 20927
rect 19393 20887 19432 20893
rect 19426 20884 19432 20887
rect 19484 20884 19490 20936
rect 19710 20927 19768 20933
rect 19710 20893 19722 20927
rect 19756 20924 19768 20927
rect 19886 20924 19892 20936
rect 19756 20896 19892 20924
rect 19756 20893 19768 20896
rect 19710 20887 19768 20893
rect 19886 20884 19892 20896
rect 19944 20924 19950 20936
rect 20070 20924 20076 20936
rect 19944 20896 20076 20924
rect 19944 20884 19950 20896
rect 20070 20884 20076 20896
rect 20128 20884 20134 20936
rect 20346 20884 20352 20936
rect 20404 20924 20410 20936
rect 20732 20933 20760 20964
rect 21358 20952 21364 20964
rect 21416 20952 21422 21004
rect 20533 20927 20591 20933
rect 20533 20924 20545 20927
rect 20404 20896 20545 20924
rect 20404 20884 20410 20896
rect 20533 20893 20545 20896
rect 20579 20893 20591 20927
rect 20533 20887 20591 20893
rect 20717 20927 20775 20933
rect 20717 20893 20729 20927
rect 20763 20893 20775 20927
rect 20898 20924 20904 20936
rect 20859 20896 20904 20924
rect 20717 20887 20775 20893
rect 20898 20884 20904 20896
rect 20956 20884 20962 20936
rect 21545 20927 21603 20933
rect 21545 20924 21557 20927
rect 21100 20896 21557 20924
rect 19521 20859 19579 20865
rect 19521 20825 19533 20859
rect 19567 20825 19579 20859
rect 19521 20819 19579 20825
rect 19613 20859 19671 20865
rect 19613 20825 19625 20859
rect 19659 20856 19671 20859
rect 20438 20856 20444 20868
rect 19659 20828 20444 20856
rect 19659 20825 19671 20828
rect 19613 20819 19671 20825
rect 18472 20760 18552 20788
rect 18693 20791 18751 20797
rect 18472 20748 18478 20760
rect 18693 20757 18705 20791
rect 18739 20757 18751 20791
rect 18693 20751 18751 20757
rect 19426 20748 19432 20800
rect 19484 20788 19490 20800
rect 19536 20788 19564 20819
rect 20438 20816 20444 20828
rect 20496 20816 20502 20868
rect 20622 20816 20628 20868
rect 20680 20856 20686 20868
rect 20806 20856 20812 20868
rect 20680 20828 20812 20856
rect 20680 20816 20686 20828
rect 20806 20816 20812 20828
rect 20864 20816 20870 20868
rect 19484 20760 19564 20788
rect 19889 20791 19947 20797
rect 19484 20748 19490 20760
rect 19889 20757 19901 20791
rect 19935 20788 19947 20791
rect 20254 20788 20260 20800
rect 19935 20760 20260 20788
rect 19935 20757 19947 20760
rect 19889 20751 19947 20757
rect 20254 20748 20260 20760
rect 20312 20748 20318 20800
rect 21100 20797 21128 20896
rect 21545 20893 21557 20896
rect 21591 20893 21603 20927
rect 21545 20887 21603 20893
rect 21634 20884 21640 20936
rect 21692 20933 21698 20936
rect 21692 20927 21723 20933
rect 21711 20893 21723 20927
rect 21692 20887 21723 20893
rect 21692 20884 21698 20887
rect 21818 20884 21824 20936
rect 21876 20924 21882 20936
rect 22010 20927 22068 20933
rect 21876 20896 21921 20924
rect 21876 20884 21882 20896
rect 22010 20893 22022 20927
rect 22056 20893 22068 20927
rect 22112 20924 22140 21032
rect 22189 21029 22201 21063
rect 22235 21029 22247 21063
rect 22189 21023 22247 21029
rect 22204 20992 22232 21023
rect 22830 21020 22836 21072
rect 22888 21060 22894 21072
rect 23753 21063 23811 21069
rect 23753 21060 23765 21063
rect 22888 21032 23765 21060
rect 22888 21020 22894 21032
rect 23753 21029 23765 21032
rect 23799 21060 23811 21063
rect 24210 21060 24216 21072
rect 23799 21032 24216 21060
rect 23799 21029 23811 21032
rect 23753 21023 23811 21029
rect 24210 21020 24216 21032
rect 24268 21020 24274 21072
rect 27614 21020 27620 21072
rect 27672 21060 27678 21072
rect 28261 21063 28319 21069
rect 28261 21060 28273 21063
rect 27672 21032 28273 21060
rect 27672 21020 27678 21032
rect 28261 21029 28273 21032
rect 28307 21060 28319 21063
rect 28810 21060 28816 21072
rect 28307 21032 28816 21060
rect 28307 21029 28319 21032
rect 28261 21023 28319 21029
rect 28810 21020 28816 21032
rect 28868 21060 28874 21072
rect 28905 21063 28963 21069
rect 28905 21060 28917 21063
rect 28868 21032 28917 21060
rect 28868 21020 28874 21032
rect 28905 21029 28917 21032
rect 28951 21029 28963 21063
rect 28905 21023 28963 21029
rect 30101 21063 30159 21069
rect 30101 21029 30113 21063
rect 30147 21060 30159 21063
rect 30944 21060 30972 21100
rect 31662 21088 31668 21100
rect 31720 21088 31726 21140
rect 31754 21088 31760 21140
rect 31812 21128 31818 21140
rect 32769 21131 32827 21137
rect 32769 21128 32781 21131
rect 31812 21100 32781 21128
rect 31812 21088 31818 21100
rect 32769 21097 32781 21100
rect 32815 21097 32827 21131
rect 34606 21128 34612 21140
rect 32769 21091 32827 21097
rect 32876 21100 34612 21128
rect 30147 21032 30972 21060
rect 32033 21063 32091 21069
rect 30147 21029 30159 21032
rect 30101 21023 30159 21029
rect 32033 21029 32045 21063
rect 32079 21060 32091 21063
rect 32876 21060 32904 21100
rect 34606 21088 34612 21100
rect 34664 21088 34670 21140
rect 34977 21131 35035 21137
rect 34977 21097 34989 21131
rect 35023 21128 35035 21131
rect 35342 21128 35348 21140
rect 35023 21100 35348 21128
rect 35023 21097 35035 21100
rect 34977 21091 35035 21097
rect 35342 21088 35348 21100
rect 35400 21088 35406 21140
rect 42978 21088 42984 21140
rect 43036 21088 43042 21140
rect 45465 21131 45523 21137
rect 45465 21097 45477 21131
rect 45511 21128 45523 21131
rect 45646 21128 45652 21140
rect 45511 21100 45652 21128
rect 45511 21097 45523 21100
rect 45465 21091 45523 21097
rect 45646 21088 45652 21100
rect 45704 21088 45710 21140
rect 48406 21128 48412 21140
rect 48367 21100 48412 21128
rect 48406 21088 48412 21100
rect 48464 21088 48470 21140
rect 49605 21131 49663 21137
rect 49605 21097 49617 21131
rect 49651 21128 49663 21131
rect 49694 21128 49700 21140
rect 49651 21100 49700 21128
rect 49651 21097 49663 21100
rect 49605 21091 49663 21097
rect 49694 21088 49700 21100
rect 49752 21088 49758 21140
rect 51718 21088 51724 21140
rect 51776 21128 51782 21140
rect 51776 21100 52408 21128
rect 51776 21088 51782 21100
rect 32079 21032 32904 21060
rect 32953 21063 33011 21069
rect 32079 21029 32091 21032
rect 32033 21023 32091 21029
rect 32953 21029 32965 21063
rect 32999 21060 33011 21063
rect 42996 21060 43024 21088
rect 45278 21060 45284 21072
rect 32999 21032 45284 21060
rect 32999 21029 33011 21032
rect 32953 21023 33011 21029
rect 45278 21020 45284 21032
rect 45336 21020 45342 21072
rect 52380 21069 52408 21100
rect 53742 21088 53748 21140
rect 53800 21128 53806 21140
rect 53929 21131 53987 21137
rect 53929 21128 53941 21131
rect 53800 21100 53941 21128
rect 53800 21088 53806 21100
rect 53929 21097 53941 21100
rect 53975 21097 53987 21131
rect 53929 21091 53987 21097
rect 52365 21063 52423 21069
rect 52365 21029 52377 21063
rect 52411 21029 52423 21063
rect 52365 21023 52423 21029
rect 51724 21004 51776 21010
rect 36909 20995 36967 21001
rect 36909 20992 36921 20995
rect 22204 20964 36921 20992
rect 36909 20961 36921 20964
rect 36955 20961 36967 20995
rect 36909 20955 36967 20961
rect 42981 20995 43039 21001
rect 42981 20961 42993 20995
rect 43027 20992 43039 20995
rect 46474 20992 46480 21004
rect 43027 20964 46480 20992
rect 43027 20961 43039 20964
rect 42981 20955 43039 20961
rect 46474 20952 46480 20964
rect 46532 20952 46538 21004
rect 48777 20995 48835 21001
rect 48148 20964 48728 20992
rect 23566 20924 23572 20936
rect 22112 20896 23572 20924
rect 22010 20887 22068 20893
rect 21913 20859 21971 20865
rect 21913 20856 21925 20859
rect 21744 20828 21925 20856
rect 21744 20800 21772 20828
rect 21913 20825 21925 20828
rect 21959 20825 21971 20859
rect 22025 20856 22053 20887
rect 23566 20884 23572 20896
rect 23624 20924 23630 20936
rect 24397 20927 24455 20933
rect 24397 20924 24409 20927
rect 23624 20896 24409 20924
rect 23624 20884 23630 20896
rect 24397 20893 24409 20896
rect 24443 20893 24455 20927
rect 24670 20924 24676 20936
rect 24583 20896 24676 20924
rect 24397 20887 24455 20893
rect 24670 20884 24676 20896
rect 24728 20924 24734 20936
rect 25406 20924 25412 20936
rect 24728 20896 25412 20924
rect 24728 20884 24734 20896
rect 25406 20884 25412 20896
rect 25464 20884 25470 20936
rect 25682 20924 25688 20936
rect 25643 20896 25688 20924
rect 25682 20884 25688 20896
rect 25740 20924 25746 20936
rect 25740 20896 26372 20924
rect 25740 20884 25746 20896
rect 22370 20856 22376 20868
rect 22025 20828 22376 20856
rect 21913 20819 21971 20825
rect 22370 20816 22376 20828
rect 22428 20816 22434 20868
rect 25958 20856 25964 20868
rect 25919 20828 25964 20856
rect 25958 20816 25964 20828
rect 26016 20816 26022 20868
rect 26344 20856 26372 20896
rect 26510 20884 26516 20936
rect 26568 20924 26574 20936
rect 26605 20927 26663 20933
rect 26605 20924 26617 20927
rect 26568 20896 26617 20924
rect 26568 20884 26574 20896
rect 26605 20893 26617 20896
rect 26651 20893 26663 20927
rect 26605 20887 26663 20893
rect 27249 20927 27307 20933
rect 27249 20893 27261 20927
rect 27295 20893 27307 20927
rect 27522 20924 27528 20936
rect 27483 20896 27528 20924
rect 27249 20887 27307 20893
rect 27264 20856 27292 20887
rect 27522 20884 27528 20896
rect 27580 20884 27586 20936
rect 27617 20927 27675 20933
rect 27617 20893 27629 20927
rect 27663 20924 27675 20927
rect 28074 20924 28080 20936
rect 27663 20896 28080 20924
rect 27663 20893 27675 20896
rect 27617 20887 27675 20893
rect 26344 20828 27292 20856
rect 27338 20816 27344 20868
rect 27396 20856 27402 20868
rect 27433 20859 27491 20865
rect 27433 20856 27445 20859
rect 27396 20828 27445 20856
rect 27396 20816 27402 20828
rect 27433 20825 27445 20828
rect 27479 20825 27491 20859
rect 27433 20819 27491 20825
rect 21085 20791 21143 20797
rect 21085 20757 21097 20791
rect 21131 20757 21143 20791
rect 21085 20751 21143 20757
rect 21726 20748 21732 20800
rect 21784 20748 21790 20800
rect 25314 20748 25320 20800
rect 25372 20788 25378 20800
rect 25777 20791 25835 20797
rect 25777 20788 25789 20791
rect 25372 20760 25789 20788
rect 25372 20748 25378 20760
rect 25777 20757 25789 20760
rect 25823 20788 25835 20791
rect 26234 20788 26240 20800
rect 25823 20760 26240 20788
rect 25823 20757 25835 20760
rect 25777 20751 25835 20757
rect 26234 20748 26240 20760
rect 26292 20748 26298 20800
rect 26697 20791 26755 20797
rect 26697 20757 26709 20791
rect 26743 20788 26755 20791
rect 27632 20788 27660 20887
rect 28074 20884 28080 20896
rect 28132 20884 28138 20936
rect 29546 20924 29552 20936
rect 29507 20896 29552 20924
rect 29546 20884 29552 20896
rect 29604 20884 29610 20936
rect 29638 20884 29644 20936
rect 29696 20924 29702 20936
rect 29822 20924 29828 20936
rect 29696 20896 29741 20924
rect 29783 20896 29828 20924
rect 29696 20884 29702 20896
rect 29822 20884 29828 20896
rect 29880 20884 29886 20936
rect 29917 20927 29975 20933
rect 29917 20893 29929 20927
rect 29963 20893 29975 20927
rect 29917 20887 29975 20893
rect 28810 20816 28816 20868
rect 28868 20856 28874 20868
rect 29932 20856 29960 20887
rect 30374 20884 30380 20936
rect 30432 20924 30438 20936
rect 30745 20927 30803 20933
rect 30745 20924 30757 20927
rect 30432 20896 30757 20924
rect 30432 20884 30438 20896
rect 30745 20893 30757 20896
rect 30791 20893 30803 20927
rect 30745 20887 30803 20893
rect 30834 20884 30840 20936
rect 30892 20924 30898 20936
rect 31573 20927 31631 20933
rect 30892 20896 30937 20924
rect 30892 20884 30898 20896
rect 31573 20893 31585 20927
rect 31619 20893 31631 20927
rect 31573 20887 31631 20893
rect 28868 20828 29960 20856
rect 31588 20856 31616 20887
rect 31754 20884 31760 20936
rect 31812 20924 31818 20936
rect 32125 20927 32183 20933
rect 31812 20896 31857 20924
rect 31812 20884 31818 20896
rect 32125 20893 32137 20927
rect 32171 20924 32183 20927
rect 32171 20896 32628 20924
rect 32171 20893 32183 20896
rect 32125 20887 32183 20893
rect 32600 20865 32628 20896
rect 34790 20884 34796 20936
rect 34848 20924 34854 20936
rect 34977 20927 35035 20933
rect 34977 20924 34989 20927
rect 34848 20896 34989 20924
rect 34848 20884 34854 20896
rect 34977 20893 34989 20896
rect 35023 20893 35035 20927
rect 36998 20924 37004 20936
rect 36959 20896 37004 20924
rect 34977 20887 35035 20893
rect 36998 20884 37004 20896
rect 37056 20884 37062 20936
rect 40218 20884 40224 20936
rect 40276 20924 40282 20936
rect 40313 20927 40371 20933
rect 40313 20924 40325 20927
rect 40276 20896 40325 20924
rect 40276 20884 40282 20896
rect 40313 20893 40325 20896
rect 40359 20893 40371 20927
rect 41966 20924 41972 20936
rect 41927 20896 41972 20924
rect 40313 20887 40371 20893
rect 41966 20884 41972 20896
rect 42024 20884 42030 20936
rect 42150 20924 42156 20936
rect 42111 20896 42156 20924
rect 42150 20884 42156 20896
rect 42208 20884 42214 20936
rect 43438 20924 43444 20936
rect 43399 20896 43444 20924
rect 43438 20884 43444 20896
rect 43496 20884 43502 20936
rect 43622 20924 43628 20936
rect 43583 20896 43628 20924
rect 43622 20884 43628 20896
rect 43680 20884 43686 20936
rect 43901 20927 43959 20933
rect 43901 20893 43913 20927
rect 43947 20924 43959 20927
rect 45002 20924 45008 20936
rect 43947 20896 44772 20924
rect 44963 20896 45008 20924
rect 43947 20893 43959 20896
rect 43901 20887 43959 20893
rect 32585 20859 32643 20865
rect 31588 20828 32260 20856
rect 28868 20816 28874 20828
rect 26743 20760 27660 20788
rect 31113 20791 31171 20797
rect 26743 20757 26755 20760
rect 26697 20751 26755 20757
rect 31113 20757 31125 20791
rect 31159 20788 31171 20791
rect 31726 20788 31754 20828
rect 31159 20760 31754 20788
rect 32232 20788 32260 20828
rect 32585 20825 32597 20859
rect 32631 20856 32643 20859
rect 32674 20856 32680 20868
rect 32631 20828 32680 20856
rect 32631 20825 32643 20828
rect 32585 20819 32643 20825
rect 32674 20816 32680 20828
rect 32732 20816 32738 20868
rect 34514 20816 34520 20868
rect 34572 20856 34578 20868
rect 34701 20859 34759 20865
rect 34701 20856 34713 20859
rect 34572 20828 34713 20856
rect 34572 20816 34578 20828
rect 34701 20825 34713 20828
rect 34747 20825 34759 20859
rect 34882 20856 34888 20868
rect 34843 20828 34888 20856
rect 34701 20819 34759 20825
rect 34882 20816 34888 20828
rect 34940 20816 34946 20868
rect 40494 20856 40500 20868
rect 40455 20828 40500 20856
rect 40494 20816 40500 20828
rect 40552 20816 40558 20868
rect 43990 20856 43996 20868
rect 43951 20828 43996 20856
rect 43990 20816 43996 20828
rect 44048 20816 44054 20868
rect 44744 20856 44772 20896
rect 45002 20884 45008 20896
rect 45060 20884 45066 20936
rect 45278 20924 45284 20936
rect 45239 20896 45284 20924
rect 45278 20884 45284 20896
rect 45336 20884 45342 20936
rect 48148 20924 48176 20964
rect 48314 20924 48320 20936
rect 45526 20896 48176 20924
rect 48275 20896 48320 20924
rect 45526 20856 45554 20896
rect 48314 20884 48320 20896
rect 48372 20884 48378 20936
rect 48700 20924 48728 20964
rect 48777 20961 48789 20995
rect 48823 20992 48835 20995
rect 51074 20992 51080 21004
rect 48823 20964 50568 20992
rect 51035 20964 51080 20992
rect 48823 20961 48835 20964
rect 48777 20955 48835 20961
rect 49234 20924 49240 20936
rect 48700 20896 49240 20924
rect 49234 20884 49240 20896
rect 49292 20884 49298 20936
rect 49421 20927 49479 20933
rect 49421 20893 49433 20927
rect 49467 20893 49479 20927
rect 50540 20924 50568 20964
rect 51074 20952 51080 20964
rect 51132 20952 51138 21004
rect 51724 20946 51776 20952
rect 51350 20924 51356 20936
rect 50540 20896 51356 20924
rect 49421 20887 49479 20893
rect 44744 20828 45554 20856
rect 47486 20816 47492 20868
rect 47544 20856 47550 20868
rect 49436 20856 49464 20887
rect 51350 20884 51356 20896
rect 51408 20884 51414 20936
rect 51994 20924 52000 20936
rect 51955 20896 52000 20924
rect 51994 20884 52000 20896
rect 52052 20884 52058 20936
rect 52380 20924 52408 21023
rect 56318 21020 56324 21072
rect 56376 21020 56382 21072
rect 56686 21020 56692 21072
rect 56744 21020 56750 21072
rect 54110 20992 54116 21004
rect 54023 20964 54116 20992
rect 54110 20952 54116 20964
rect 54168 20992 54174 21004
rect 54386 20992 54392 21004
rect 54168 20964 54392 20992
rect 54168 20952 54174 20964
rect 54386 20952 54392 20964
rect 54444 20952 54450 21004
rect 56336 20992 56364 21020
rect 56704 20992 56732 21020
rect 56336 20964 56548 20992
rect 56704 20964 56916 20992
rect 53837 20927 53895 20933
rect 53837 20924 53849 20927
rect 52380 20896 53849 20924
rect 53837 20893 53849 20896
rect 53883 20893 53895 20927
rect 53837 20887 53895 20893
rect 54202 20884 54208 20936
rect 54260 20924 54266 20936
rect 55674 20924 55680 20936
rect 54260 20896 54305 20924
rect 55186 20896 55680 20924
rect 54260 20884 54266 20896
rect 47544 20828 49464 20856
rect 54297 20859 54355 20865
rect 47544 20816 47550 20828
rect 54297 20825 54309 20859
rect 54343 20856 54355 20859
rect 55186 20856 55214 20896
rect 55674 20884 55680 20896
rect 55732 20884 55738 20936
rect 56226 20884 56232 20936
rect 56284 20924 56290 20936
rect 56520 20933 56548 20964
rect 56367 20927 56425 20933
rect 56367 20924 56379 20927
rect 56284 20896 56379 20924
rect 56284 20884 56290 20896
rect 56367 20893 56379 20896
rect 56413 20893 56425 20927
rect 56367 20887 56425 20893
rect 56505 20927 56563 20933
rect 56505 20893 56517 20927
rect 56551 20893 56563 20927
rect 56778 20924 56784 20936
rect 56739 20896 56784 20924
rect 56505 20887 56563 20893
rect 56778 20884 56784 20896
rect 56836 20884 56842 20936
rect 56888 20933 56916 20964
rect 57698 20952 57704 21004
rect 57756 20992 57762 21004
rect 57885 20995 57943 21001
rect 57885 20992 57897 20995
rect 57756 20964 57897 20992
rect 57756 20952 57762 20964
rect 57885 20961 57897 20964
rect 57931 20961 57943 20995
rect 57885 20955 57943 20961
rect 56873 20927 56931 20933
rect 56873 20893 56885 20927
rect 56919 20893 56931 20927
rect 58158 20924 58164 20936
rect 58119 20896 58164 20924
rect 56873 20887 56931 20893
rect 58158 20884 58164 20896
rect 58216 20884 58222 20936
rect 55490 20856 55496 20868
rect 54343 20828 55214 20856
rect 55403 20828 55496 20856
rect 54343 20825 54355 20828
rect 54297 20819 54355 20825
rect 55490 20816 55496 20828
rect 55548 20856 55554 20868
rect 56594 20856 56600 20868
rect 55548 20828 56364 20856
rect 56555 20828 56600 20856
rect 55548 20816 55554 20828
rect 32769 20791 32827 20797
rect 32769 20788 32781 20791
rect 32232 20760 32781 20788
rect 31159 20757 31171 20760
rect 31113 20751 31171 20757
rect 32769 20757 32781 20760
rect 32815 20757 32827 20791
rect 37366 20788 37372 20800
rect 37327 20760 37372 20788
rect 32769 20751 32827 20757
rect 37366 20748 37372 20760
rect 37424 20748 37430 20800
rect 45094 20788 45100 20800
rect 45055 20760 45100 20788
rect 45094 20748 45100 20760
rect 45152 20748 45158 20800
rect 56226 20788 56232 20800
rect 56187 20760 56232 20788
rect 56226 20748 56232 20760
rect 56284 20748 56290 20800
rect 56336 20788 56364 20828
rect 56594 20816 56600 20828
rect 56652 20816 56658 20868
rect 56686 20816 56692 20868
rect 56744 20856 56750 20868
rect 56962 20856 56968 20868
rect 56744 20828 56968 20856
rect 56744 20816 56750 20828
rect 56962 20816 56968 20828
rect 57020 20816 57026 20868
rect 56704 20788 56732 20816
rect 56336 20760 56732 20788
rect 1104 20698 58880 20720
rect 1104 20646 19574 20698
rect 19626 20646 19638 20698
rect 19690 20646 19702 20698
rect 19754 20646 19766 20698
rect 19818 20646 19830 20698
rect 19882 20646 50294 20698
rect 50346 20646 50358 20698
rect 50410 20646 50422 20698
rect 50474 20646 50486 20698
rect 50538 20646 50550 20698
rect 50602 20646 58880 20698
rect 1104 20624 58880 20646
rect 3053 20587 3111 20593
rect 3053 20584 3065 20587
rect 2746 20556 3065 20584
rect 1486 20476 1492 20528
rect 1544 20516 1550 20528
rect 2222 20516 2228 20528
rect 1544 20488 2228 20516
rect 1544 20476 1550 20488
rect 2222 20476 2228 20488
rect 2280 20516 2286 20528
rect 2317 20519 2375 20525
rect 2317 20516 2329 20519
rect 2280 20488 2329 20516
rect 2280 20476 2286 20488
rect 2317 20485 2329 20488
rect 2363 20485 2375 20519
rect 2746 20516 2774 20556
rect 3053 20553 3065 20556
rect 3099 20584 3111 20587
rect 5258 20584 5264 20596
rect 3099 20556 5264 20584
rect 3099 20553 3111 20556
rect 3053 20547 3111 20553
rect 5258 20544 5264 20556
rect 5316 20544 5322 20596
rect 7466 20544 7472 20596
rect 7524 20584 7530 20596
rect 7929 20587 7987 20593
rect 7929 20584 7941 20587
rect 7524 20556 7941 20584
rect 7524 20544 7530 20556
rect 7929 20553 7941 20556
rect 7975 20584 7987 20587
rect 8202 20584 8208 20596
rect 7975 20556 8208 20584
rect 7975 20553 7987 20556
rect 7929 20547 7987 20553
rect 8202 20544 8208 20556
rect 8260 20544 8266 20596
rect 14642 20584 14648 20596
rect 14603 20556 14648 20584
rect 14642 20544 14648 20556
rect 14700 20544 14706 20596
rect 18049 20587 18107 20593
rect 18049 20553 18061 20587
rect 18095 20584 18107 20587
rect 18230 20584 18236 20596
rect 18095 20556 18236 20584
rect 18095 20553 18107 20556
rect 18049 20547 18107 20553
rect 18230 20544 18236 20556
rect 18288 20544 18294 20596
rect 18601 20587 18659 20593
rect 18601 20553 18613 20587
rect 18647 20584 18659 20587
rect 19058 20584 19064 20596
rect 18647 20556 19064 20584
rect 18647 20553 18659 20556
rect 18601 20547 18659 20553
rect 19058 20544 19064 20556
rect 19116 20544 19122 20596
rect 19150 20544 19156 20596
rect 19208 20584 19214 20596
rect 21726 20584 21732 20596
rect 19208 20556 21732 20584
rect 19208 20544 19214 20556
rect 21726 20544 21732 20556
rect 21784 20584 21790 20596
rect 21821 20587 21879 20593
rect 21821 20584 21833 20587
rect 21784 20556 21833 20584
rect 21784 20544 21790 20556
rect 21821 20553 21833 20556
rect 21867 20553 21879 20587
rect 21821 20547 21879 20553
rect 21910 20544 21916 20596
rect 21968 20584 21974 20596
rect 22370 20584 22376 20596
rect 21968 20556 22376 20584
rect 21968 20544 21974 20556
rect 22370 20544 22376 20556
rect 22428 20544 22434 20596
rect 24121 20587 24179 20593
rect 24121 20553 24133 20587
rect 24167 20584 24179 20587
rect 24302 20584 24308 20596
rect 24167 20556 24308 20584
rect 24167 20553 24179 20556
rect 24121 20547 24179 20553
rect 24302 20544 24308 20556
rect 24360 20544 24366 20596
rect 26510 20544 26516 20596
rect 26568 20584 26574 20596
rect 26973 20587 27031 20593
rect 26973 20584 26985 20587
rect 26568 20556 26985 20584
rect 26568 20544 26574 20556
rect 26973 20553 26985 20556
rect 27019 20553 27031 20587
rect 26973 20547 27031 20553
rect 29181 20587 29239 20593
rect 29181 20553 29193 20587
rect 29227 20584 29239 20587
rect 29638 20584 29644 20596
rect 29227 20556 29644 20584
rect 29227 20553 29239 20556
rect 29181 20547 29239 20553
rect 29638 20544 29644 20556
rect 29696 20544 29702 20596
rect 31205 20587 31263 20593
rect 31205 20553 31217 20587
rect 31251 20584 31263 20587
rect 31754 20584 31760 20596
rect 31251 20556 31760 20584
rect 31251 20553 31263 20556
rect 31205 20547 31263 20553
rect 31754 20544 31760 20556
rect 31812 20544 31818 20596
rect 33965 20587 34023 20593
rect 33965 20553 33977 20587
rect 34011 20584 34023 20587
rect 34517 20587 34575 20593
rect 34517 20584 34529 20587
rect 34011 20556 34529 20584
rect 34011 20553 34023 20556
rect 33965 20547 34023 20553
rect 34517 20553 34529 20556
rect 34563 20584 34575 20587
rect 34882 20584 34888 20596
rect 34563 20556 34888 20584
rect 34563 20553 34575 20556
rect 34517 20547 34575 20553
rect 34882 20544 34888 20556
rect 34940 20544 34946 20596
rect 40865 20587 40923 20593
rect 40865 20553 40877 20587
rect 40911 20584 40923 20587
rect 41966 20584 41972 20596
rect 40911 20556 41972 20584
rect 40911 20553 40923 20556
rect 40865 20547 40923 20553
rect 41966 20544 41972 20556
rect 42024 20544 42030 20596
rect 43717 20587 43775 20593
rect 43717 20553 43729 20587
rect 43763 20584 43775 20587
rect 47486 20584 47492 20596
rect 43763 20556 47492 20584
rect 43763 20553 43775 20556
rect 43717 20547 43775 20553
rect 47486 20544 47492 20556
rect 47544 20544 47550 20596
rect 51810 20584 51816 20596
rect 51771 20556 51816 20584
rect 51810 20544 51816 20556
rect 51868 20544 51874 20596
rect 57054 20544 57060 20596
rect 57112 20584 57118 20596
rect 57149 20587 57207 20593
rect 57149 20584 57161 20587
rect 57112 20556 57161 20584
rect 57112 20544 57118 20556
rect 57149 20553 57161 20556
rect 57195 20553 57207 20587
rect 57149 20547 57207 20553
rect 10410 20516 10416 20528
rect 2317 20479 2375 20485
rect 2424 20488 2774 20516
rect 10371 20488 10416 20516
rect 2130 20448 2136 20460
rect 2043 20420 2136 20448
rect 2130 20408 2136 20420
rect 2188 20448 2194 20460
rect 2424 20448 2452 20488
rect 10410 20476 10416 20488
rect 10468 20476 10474 20528
rect 13449 20519 13507 20525
rect 13449 20485 13461 20519
rect 13495 20516 13507 20519
rect 13814 20516 13820 20528
rect 13495 20488 13820 20516
rect 13495 20485 13507 20488
rect 13449 20479 13507 20485
rect 13814 20476 13820 20488
rect 13872 20476 13878 20528
rect 2188 20420 2452 20448
rect 2188 20408 2194 20420
rect 2498 20408 2504 20460
rect 2556 20448 2562 20460
rect 4065 20451 4123 20457
rect 4065 20448 4077 20451
rect 2556 20420 4077 20448
rect 2556 20408 2562 20420
rect 4065 20417 4077 20420
rect 4111 20417 4123 20451
rect 4065 20411 4123 20417
rect 4249 20451 4307 20457
rect 4249 20417 4261 20451
rect 4295 20448 4307 20451
rect 6454 20448 6460 20460
rect 4295 20420 6460 20448
rect 4295 20417 4307 20420
rect 4249 20411 4307 20417
rect 6454 20408 6460 20420
rect 6512 20408 6518 20460
rect 7834 20448 7840 20460
rect 7795 20420 7840 20448
rect 7834 20408 7840 20420
rect 7892 20408 7898 20460
rect 8018 20408 8024 20460
rect 8076 20448 8082 20460
rect 8113 20451 8171 20457
rect 8113 20448 8125 20451
rect 8076 20420 8125 20448
rect 8076 20408 8082 20420
rect 8113 20417 8125 20420
rect 8159 20417 8171 20451
rect 8113 20411 8171 20417
rect 9490 20408 9496 20460
rect 9548 20448 9554 20460
rect 9677 20451 9735 20457
rect 9677 20448 9689 20451
rect 9548 20420 9689 20448
rect 9548 20408 9554 20420
rect 9677 20417 9689 20420
rect 9723 20417 9735 20451
rect 9950 20448 9956 20460
rect 9911 20420 9956 20448
rect 9677 20411 9735 20417
rect 9950 20408 9956 20420
rect 10008 20448 10014 20460
rect 10318 20448 10324 20460
rect 10008 20420 10324 20448
rect 10008 20408 10014 20420
rect 10318 20408 10324 20420
rect 10376 20408 10382 20460
rect 12618 20408 12624 20460
rect 12676 20448 12682 20460
rect 13265 20451 13323 20457
rect 13265 20448 13277 20451
rect 12676 20420 13277 20448
rect 12676 20408 12682 20420
rect 13265 20417 13277 20420
rect 13311 20417 13323 20451
rect 13265 20411 13323 20417
rect 13354 20408 13360 20460
rect 13412 20448 13418 20460
rect 13567 20451 13625 20457
rect 13567 20448 13579 20451
rect 13412 20420 13457 20448
rect 13412 20408 13418 20420
rect 13556 20417 13579 20448
rect 13613 20417 13625 20451
rect 13556 20411 13625 20417
rect 3970 20380 3976 20392
rect 3931 20352 3976 20380
rect 3970 20340 3976 20352
rect 4028 20340 4034 20392
rect 4157 20383 4215 20389
rect 4157 20349 4169 20383
rect 4203 20349 4215 20383
rect 4157 20343 4215 20349
rect 4062 20272 4068 20324
rect 4120 20312 4126 20324
rect 4172 20312 4200 20343
rect 8113 20315 8171 20321
rect 4120 20284 4200 20312
rect 4356 20284 8064 20312
rect 4120 20272 4126 20284
rect 1946 20204 1952 20256
rect 2004 20244 2010 20256
rect 4356 20244 4384 20284
rect 2004 20216 4384 20244
rect 4433 20247 4491 20253
rect 2004 20204 2010 20216
rect 4433 20213 4445 20247
rect 4479 20244 4491 20247
rect 4890 20244 4896 20256
rect 4479 20216 4896 20244
rect 4479 20213 4491 20216
rect 4433 20207 4491 20213
rect 4890 20204 4896 20216
rect 4948 20204 4954 20256
rect 8036 20244 8064 20284
rect 8113 20281 8125 20315
rect 8159 20312 8171 20315
rect 9674 20312 9680 20324
rect 8159 20284 9680 20312
rect 8159 20281 8171 20284
rect 8113 20275 8171 20281
rect 9674 20272 9680 20284
rect 9732 20312 9738 20324
rect 9769 20315 9827 20321
rect 9769 20312 9781 20315
rect 9732 20284 9781 20312
rect 9732 20272 9738 20284
rect 9769 20281 9781 20284
rect 9815 20281 9827 20315
rect 13078 20312 13084 20324
rect 13039 20284 13084 20312
rect 9769 20275 9827 20281
rect 13078 20272 13084 20284
rect 13136 20272 13142 20324
rect 13556 20256 13584 20411
rect 13722 20408 13728 20460
rect 13780 20448 13786 20460
rect 18248 20448 18276 20544
rect 18322 20476 18328 20528
rect 18380 20516 18386 20528
rect 18380 20488 18644 20516
rect 18380 20476 18386 20488
rect 18616 20460 18644 20488
rect 24210 20476 24216 20528
rect 24268 20516 24274 20528
rect 25314 20516 25320 20528
rect 24268 20488 25320 20516
rect 24268 20476 24274 20488
rect 25314 20476 25320 20488
rect 25372 20476 25378 20528
rect 25682 20476 25688 20528
rect 25740 20516 25746 20528
rect 26053 20519 26111 20525
rect 26053 20516 26065 20519
rect 25740 20488 26065 20516
rect 25740 20476 25746 20488
rect 26053 20485 26065 20488
rect 26099 20485 26111 20519
rect 26053 20479 26111 20485
rect 27338 20476 27344 20528
rect 27396 20516 27402 20528
rect 27709 20519 27767 20525
rect 27709 20516 27721 20519
rect 27396 20488 27721 20516
rect 27396 20476 27402 20488
rect 27709 20485 27721 20488
rect 27755 20485 27767 20519
rect 27709 20479 27767 20485
rect 28813 20519 28871 20525
rect 28813 20485 28825 20519
rect 28859 20516 28871 20519
rect 28859 20488 28948 20516
rect 28859 20485 28871 20488
rect 28813 20479 28871 20485
rect 18509 20451 18567 20457
rect 18509 20448 18521 20451
rect 13780 20420 13825 20448
rect 18248 20420 18521 20448
rect 13780 20408 13786 20420
rect 18509 20417 18521 20420
rect 18555 20417 18567 20451
rect 18509 20411 18567 20417
rect 18598 20408 18604 20460
rect 18656 20448 18662 20460
rect 18693 20451 18751 20457
rect 18693 20448 18705 20451
rect 18656 20420 18705 20448
rect 18656 20408 18662 20420
rect 18693 20417 18705 20420
rect 18739 20417 18751 20451
rect 18693 20411 18751 20417
rect 19521 20451 19579 20457
rect 19521 20417 19533 20451
rect 19567 20448 19579 20451
rect 19978 20448 19984 20460
rect 19567 20420 19984 20448
rect 19567 20417 19579 20420
rect 19521 20411 19579 20417
rect 19978 20408 19984 20420
rect 20036 20408 20042 20460
rect 20257 20451 20315 20457
rect 20257 20417 20269 20451
rect 20303 20448 20315 20451
rect 20438 20448 20444 20460
rect 20303 20420 20444 20448
rect 20303 20417 20315 20420
rect 20257 20411 20315 20417
rect 20438 20408 20444 20420
rect 20496 20408 20502 20460
rect 18414 20380 18420 20392
rect 13648 20352 18420 20380
rect 13648 20324 13676 20352
rect 18414 20340 18420 20352
rect 18472 20340 18478 20392
rect 28920 20380 28948 20488
rect 28994 20476 29000 20528
rect 29052 20525 29058 20528
rect 29052 20519 29071 20525
rect 29059 20516 29071 20519
rect 32953 20519 33011 20525
rect 32953 20516 32965 20519
rect 29059 20488 29960 20516
rect 29059 20485 29071 20488
rect 29052 20479 29071 20485
rect 29052 20476 29058 20479
rect 29638 20448 29644 20460
rect 29599 20420 29644 20448
rect 29638 20408 29644 20420
rect 29696 20408 29702 20460
rect 29932 20457 29960 20488
rect 31726 20488 32965 20516
rect 29825 20451 29883 20457
rect 29825 20417 29837 20451
rect 29871 20417 29883 20451
rect 29825 20411 29883 20417
rect 29917 20451 29975 20457
rect 29917 20417 29929 20451
rect 29963 20448 29975 20451
rect 30098 20448 30104 20460
rect 29963 20420 30104 20448
rect 29963 20417 29975 20420
rect 29917 20411 29975 20417
rect 29840 20380 29868 20411
rect 30098 20408 30104 20420
rect 30156 20408 30162 20460
rect 30742 20408 30748 20460
rect 30800 20448 30806 20460
rect 30929 20451 30987 20457
rect 30929 20448 30941 20451
rect 30800 20420 30941 20448
rect 30800 20408 30806 20420
rect 30929 20417 30941 20420
rect 30975 20417 30987 20451
rect 30929 20411 30987 20417
rect 30374 20380 30380 20392
rect 28920 20352 29960 20380
rect 30335 20352 30380 20380
rect 13630 20272 13636 20324
rect 13688 20272 13694 20324
rect 15194 20272 15200 20324
rect 15252 20312 15258 20324
rect 18138 20312 18144 20324
rect 15252 20284 18144 20312
rect 15252 20272 15258 20284
rect 18138 20272 18144 20284
rect 18196 20312 18202 20324
rect 19150 20312 19156 20324
rect 18196 20284 19156 20312
rect 18196 20272 18202 20284
rect 19150 20272 19156 20284
rect 19208 20312 19214 20324
rect 19337 20315 19395 20321
rect 19337 20312 19349 20315
rect 19208 20284 19349 20312
rect 19208 20272 19214 20284
rect 19337 20281 19349 20284
rect 19383 20281 19395 20315
rect 19337 20275 19395 20281
rect 29546 20272 29552 20324
rect 29604 20312 29610 20324
rect 29641 20315 29699 20321
rect 29641 20312 29653 20315
rect 29604 20284 29653 20312
rect 29604 20272 29610 20284
rect 29641 20281 29653 20284
rect 29687 20281 29699 20315
rect 29932 20312 29960 20352
rect 30374 20340 30380 20352
rect 30432 20340 30438 20392
rect 30834 20340 30840 20392
rect 30892 20380 30898 20392
rect 31205 20383 31263 20389
rect 31205 20380 31217 20383
rect 30892 20352 31217 20380
rect 30892 20340 30898 20352
rect 31205 20349 31217 20352
rect 31251 20380 31263 20383
rect 31726 20380 31754 20488
rect 32953 20485 32965 20488
rect 32999 20485 33011 20519
rect 32953 20479 33011 20485
rect 31251 20352 31754 20380
rect 32968 20380 32996 20479
rect 33410 20476 33416 20528
rect 33468 20516 33474 20528
rect 33597 20519 33655 20525
rect 33597 20516 33609 20519
rect 33468 20488 33609 20516
rect 33468 20476 33474 20488
rect 33597 20485 33609 20488
rect 33643 20485 33655 20519
rect 33597 20479 33655 20485
rect 39209 20519 39267 20525
rect 39209 20485 39221 20519
rect 39255 20516 39267 20519
rect 42150 20516 42156 20528
rect 39255 20488 42156 20516
rect 39255 20485 39267 20488
rect 39209 20479 39267 20485
rect 42150 20476 42156 20488
rect 42208 20516 42214 20528
rect 42429 20519 42487 20525
rect 42429 20516 42441 20519
rect 42208 20488 42441 20516
rect 42208 20476 42214 20488
rect 42429 20485 42441 20488
rect 42475 20485 42487 20519
rect 44913 20519 44971 20525
rect 42429 20479 42487 20485
rect 43180 20488 44312 20516
rect 33502 20448 33508 20460
rect 33463 20420 33508 20448
rect 33502 20408 33508 20420
rect 33560 20408 33566 20460
rect 33781 20451 33839 20457
rect 33781 20417 33793 20451
rect 33827 20417 33839 20451
rect 33781 20411 33839 20417
rect 34425 20451 34483 20457
rect 34425 20417 34437 20451
rect 34471 20448 34483 20451
rect 34514 20448 34520 20460
rect 34471 20420 34520 20448
rect 34471 20417 34483 20420
rect 34425 20411 34483 20417
rect 33796 20380 33824 20411
rect 34514 20408 34520 20420
rect 34572 20408 34578 20460
rect 34698 20448 34704 20460
rect 34659 20420 34704 20448
rect 34698 20408 34704 20420
rect 34756 20408 34762 20460
rect 37366 20408 37372 20460
rect 37424 20448 37430 20460
rect 38286 20448 38292 20460
rect 37424 20420 38292 20448
rect 37424 20408 37430 20420
rect 38286 20408 38292 20420
rect 38344 20448 38350 20460
rect 38381 20451 38439 20457
rect 38381 20448 38393 20451
rect 38344 20420 38393 20448
rect 38344 20408 38350 20420
rect 38381 20417 38393 20420
rect 38427 20417 38439 20451
rect 40494 20448 40500 20460
rect 40455 20420 40500 20448
rect 38381 20411 38439 20417
rect 40494 20408 40500 20420
rect 40552 20408 40558 20460
rect 43180 20448 43208 20488
rect 43346 20448 43352 20460
rect 41892 20420 43208 20448
rect 43307 20420 43352 20448
rect 34790 20380 34796 20392
rect 32968 20352 34796 20380
rect 31251 20349 31263 20352
rect 31205 20343 31263 20349
rect 34790 20340 34796 20352
rect 34848 20340 34854 20392
rect 38470 20380 38476 20392
rect 38431 20352 38476 20380
rect 38470 20340 38476 20352
rect 38528 20340 38534 20392
rect 39758 20340 39764 20392
rect 39816 20380 39822 20392
rect 40405 20383 40463 20389
rect 40405 20380 40417 20383
rect 39816 20352 40417 20380
rect 39816 20340 39822 20352
rect 40405 20349 40417 20352
rect 40451 20349 40463 20383
rect 40405 20343 40463 20349
rect 31754 20312 31760 20324
rect 29932 20284 31760 20312
rect 29641 20275 29699 20281
rect 31754 20272 31760 20284
rect 31812 20272 31818 20324
rect 34885 20315 34943 20321
rect 34885 20281 34897 20315
rect 34931 20312 34943 20315
rect 41892 20312 41920 20420
rect 43346 20408 43352 20420
rect 43404 20448 43410 20460
rect 43990 20448 43996 20460
rect 43404 20420 43996 20448
rect 43404 20408 43410 20420
rect 43990 20408 43996 20420
rect 44048 20448 44054 20460
rect 44177 20451 44235 20457
rect 44177 20448 44189 20451
rect 44048 20420 44189 20448
rect 44048 20408 44054 20420
rect 44177 20417 44189 20420
rect 44223 20417 44235 20451
rect 44284 20448 44312 20488
rect 44913 20485 44925 20519
rect 44959 20516 44971 20519
rect 45002 20516 45008 20528
rect 44959 20488 45008 20516
rect 44959 20485 44971 20488
rect 44913 20479 44971 20485
rect 45002 20476 45008 20488
rect 45060 20476 45066 20528
rect 57238 20516 57244 20528
rect 57199 20488 57244 20516
rect 57238 20476 57244 20488
rect 57296 20476 57302 20528
rect 58158 20516 58164 20528
rect 58119 20488 58164 20516
rect 58158 20476 58164 20488
rect 58216 20476 58222 20528
rect 45094 20448 45100 20460
rect 44284 20420 45100 20448
rect 44177 20411 44235 20417
rect 45094 20408 45100 20420
rect 45152 20408 45158 20460
rect 45189 20451 45247 20457
rect 45189 20417 45201 20451
rect 45235 20448 45247 20451
rect 45278 20448 45284 20460
rect 45235 20420 45284 20448
rect 45235 20417 45247 20420
rect 45189 20411 45247 20417
rect 45278 20408 45284 20420
rect 45336 20408 45342 20460
rect 51074 20408 51080 20460
rect 51132 20448 51138 20460
rect 51169 20451 51227 20457
rect 51169 20448 51181 20451
rect 51132 20420 51181 20448
rect 51132 20408 51138 20420
rect 51169 20417 51181 20420
rect 51215 20417 51227 20451
rect 51350 20448 51356 20460
rect 51311 20420 51356 20448
rect 51169 20411 51227 20417
rect 51350 20408 51356 20420
rect 51408 20408 51414 20460
rect 51445 20451 51503 20457
rect 51445 20417 51457 20451
rect 51491 20417 51503 20451
rect 51445 20411 51503 20417
rect 51537 20451 51595 20457
rect 51537 20417 51549 20451
rect 51583 20448 51595 20451
rect 51718 20448 51724 20460
rect 51583 20420 51724 20448
rect 51583 20417 51595 20420
rect 51537 20411 51595 20417
rect 43438 20380 43444 20392
rect 43399 20352 43444 20380
rect 43438 20340 43444 20352
rect 43496 20340 43502 20392
rect 51460 20380 51488 20411
rect 51718 20408 51724 20420
rect 51776 20408 51782 20460
rect 56962 20448 56968 20460
rect 56923 20420 56968 20448
rect 56962 20408 56968 20420
rect 57020 20408 57026 20460
rect 51994 20380 52000 20392
rect 51460 20352 52000 20380
rect 51994 20340 52000 20352
rect 52052 20340 52058 20392
rect 34931 20284 41920 20312
rect 34931 20281 34943 20284
rect 34885 20275 34943 20281
rect 41966 20272 41972 20324
rect 42024 20312 42030 20324
rect 42705 20315 42763 20321
rect 42705 20312 42717 20315
rect 42024 20284 42717 20312
rect 42024 20272 42030 20284
rect 42705 20281 42717 20284
rect 42751 20281 42763 20315
rect 42705 20275 42763 20281
rect 45189 20315 45247 20321
rect 45189 20281 45201 20315
rect 45235 20312 45247 20315
rect 45830 20312 45836 20324
rect 45235 20284 45836 20312
rect 45235 20281 45247 20284
rect 45189 20275 45247 20281
rect 45830 20272 45836 20284
rect 45888 20272 45894 20324
rect 11146 20244 11152 20256
rect 8036 20216 11152 20244
rect 11146 20204 11152 20216
rect 11204 20204 11210 20256
rect 13538 20204 13544 20256
rect 13596 20244 13602 20256
rect 15746 20244 15752 20256
rect 13596 20216 15752 20244
rect 13596 20204 13602 20216
rect 15746 20204 15752 20216
rect 15804 20204 15810 20256
rect 18322 20204 18328 20256
rect 18380 20244 18386 20256
rect 20073 20247 20131 20253
rect 20073 20244 20085 20247
rect 18380 20216 20085 20244
rect 18380 20204 18386 20216
rect 20073 20213 20085 20216
rect 20119 20213 20131 20247
rect 25958 20244 25964 20256
rect 25919 20216 25964 20244
rect 20073 20207 20131 20213
rect 25958 20204 25964 20216
rect 26016 20204 26022 20256
rect 26050 20204 26056 20256
rect 26108 20244 26114 20256
rect 27706 20244 27712 20256
rect 26108 20216 27712 20244
rect 26108 20204 26114 20216
rect 27706 20204 27712 20216
rect 27764 20204 27770 20256
rect 27801 20247 27859 20253
rect 27801 20213 27813 20247
rect 27847 20244 27859 20247
rect 28258 20244 28264 20256
rect 27847 20216 28264 20244
rect 27847 20213 27859 20216
rect 27801 20207 27859 20213
rect 28258 20204 28264 20216
rect 28316 20204 28322 20256
rect 28997 20247 29055 20253
rect 28997 20213 29009 20247
rect 29043 20244 29055 20247
rect 29086 20244 29092 20256
rect 29043 20216 29092 20244
rect 29043 20213 29055 20216
rect 28997 20207 29055 20213
rect 29086 20204 29092 20216
rect 29144 20244 29150 20256
rect 29730 20244 29736 20256
rect 29144 20216 29736 20244
rect 29144 20204 29150 20216
rect 29730 20204 29736 20216
rect 29788 20204 29794 20256
rect 30374 20204 30380 20256
rect 30432 20244 30438 20256
rect 31021 20247 31079 20253
rect 31021 20244 31033 20247
rect 30432 20216 31033 20244
rect 30432 20204 30438 20216
rect 31021 20213 31033 20216
rect 31067 20213 31079 20247
rect 39758 20244 39764 20256
rect 39719 20216 39764 20244
rect 31021 20207 31079 20213
rect 39758 20204 39764 20216
rect 39816 20204 39822 20256
rect 42889 20247 42947 20253
rect 42889 20213 42901 20247
rect 42935 20244 42947 20247
rect 43533 20247 43591 20253
rect 43533 20244 43545 20247
rect 42935 20216 43545 20244
rect 42935 20213 42947 20216
rect 42889 20207 42947 20213
rect 43533 20213 43545 20216
rect 43579 20244 43591 20247
rect 43622 20244 43628 20256
rect 43579 20216 43628 20244
rect 43579 20213 43591 20216
rect 43533 20207 43591 20213
rect 43622 20204 43628 20216
rect 43680 20204 43686 20256
rect 54018 20204 54024 20256
rect 54076 20244 54082 20256
rect 56781 20247 56839 20253
rect 56781 20244 56793 20247
rect 54076 20216 56793 20244
rect 54076 20204 54082 20216
rect 56781 20213 56793 20216
rect 56827 20213 56839 20247
rect 56781 20207 56839 20213
rect 1104 20154 58880 20176
rect 1104 20102 4214 20154
rect 4266 20102 4278 20154
rect 4330 20102 4342 20154
rect 4394 20102 4406 20154
rect 4458 20102 4470 20154
rect 4522 20102 34934 20154
rect 34986 20102 34998 20154
rect 35050 20102 35062 20154
rect 35114 20102 35126 20154
rect 35178 20102 35190 20154
rect 35242 20102 58880 20154
rect 1104 20080 58880 20102
rect 3970 20000 3976 20052
rect 4028 20040 4034 20052
rect 4709 20043 4767 20049
rect 4709 20040 4721 20043
rect 4028 20012 4721 20040
rect 4028 20000 4034 20012
rect 4709 20009 4721 20012
rect 4755 20040 4767 20043
rect 5353 20043 5411 20049
rect 5353 20040 5365 20043
rect 4755 20012 5365 20040
rect 4755 20009 4767 20012
rect 4709 20003 4767 20009
rect 5353 20009 5365 20012
rect 5399 20009 5411 20043
rect 5353 20003 5411 20009
rect 5442 20000 5448 20052
rect 5500 20040 5506 20052
rect 8202 20040 8208 20052
rect 5500 20012 6040 20040
rect 8163 20012 8208 20040
rect 5500 20000 5506 20012
rect 3068 19944 5948 19972
rect 2866 19768 2872 19780
rect 2827 19740 2872 19768
rect 2866 19728 2872 19740
rect 2924 19728 2930 19780
rect 3068 19777 3096 19944
rect 5258 19864 5264 19916
rect 5316 19904 5322 19916
rect 5721 19907 5779 19913
rect 5721 19904 5733 19907
rect 5316 19876 5733 19904
rect 5316 19864 5322 19876
rect 5721 19873 5733 19876
rect 5767 19873 5779 19907
rect 5721 19867 5779 19873
rect 3237 19839 3295 19845
rect 3237 19805 3249 19839
rect 3283 19836 3295 19839
rect 4062 19836 4068 19848
rect 3283 19808 4068 19836
rect 3283 19805 3295 19808
rect 3237 19799 3295 19805
rect 4062 19796 4068 19808
rect 4120 19836 4126 19848
rect 4433 19839 4491 19845
rect 4433 19836 4445 19839
rect 4120 19808 4445 19836
rect 4120 19796 4126 19808
rect 4433 19805 4445 19808
rect 4479 19805 4491 19839
rect 4433 19799 4491 19805
rect 5534 19796 5540 19848
rect 5592 19836 5598 19848
rect 5920 19836 5948 19944
rect 6012 19904 6040 20012
rect 8202 20000 8208 20012
rect 8260 20000 8266 20052
rect 12986 20040 12992 20052
rect 8312 20012 12992 20040
rect 6914 19932 6920 19984
rect 6972 19972 6978 19984
rect 7193 19975 7251 19981
rect 7193 19972 7205 19975
rect 6972 19944 7205 19972
rect 6972 19932 6978 19944
rect 7193 19941 7205 19944
rect 7239 19972 7251 19975
rect 8110 19972 8116 19984
rect 7239 19944 8116 19972
rect 7239 19941 7251 19944
rect 7193 19935 7251 19941
rect 8110 19932 8116 19944
rect 8168 19932 8174 19984
rect 8312 19904 8340 20012
rect 12986 20000 12992 20012
rect 13044 20000 13050 20052
rect 13538 20040 13544 20052
rect 13499 20012 13544 20040
rect 13538 20000 13544 20012
rect 13596 20000 13602 20052
rect 14642 20000 14648 20052
rect 14700 20040 14706 20052
rect 15381 20043 15439 20049
rect 15381 20040 15393 20043
rect 14700 20012 15393 20040
rect 14700 20000 14706 20012
rect 15381 20009 15393 20012
rect 15427 20040 15439 20043
rect 16758 20040 16764 20052
rect 15427 20012 16764 20040
rect 15427 20009 15439 20012
rect 15381 20003 15439 20009
rect 16758 20000 16764 20012
rect 16816 20040 16822 20052
rect 26050 20040 26056 20052
rect 16816 20012 26056 20040
rect 16816 20000 16822 20012
rect 26050 20000 26056 20012
rect 26108 20000 26114 20052
rect 26510 20000 26516 20052
rect 26568 20040 26574 20052
rect 26605 20043 26663 20049
rect 26605 20040 26617 20043
rect 26568 20012 26617 20040
rect 26568 20000 26574 20012
rect 26605 20009 26617 20012
rect 26651 20009 26663 20043
rect 34149 20043 34207 20049
rect 26605 20003 26663 20009
rect 26804 20012 34100 20040
rect 11425 19975 11483 19981
rect 11425 19941 11437 19975
rect 11471 19972 11483 19975
rect 16301 19975 16359 19981
rect 16301 19972 16313 19975
rect 11471 19944 16313 19972
rect 11471 19941 11483 19944
rect 11425 19935 11483 19941
rect 16301 19941 16313 19944
rect 16347 19941 16359 19975
rect 20070 19972 20076 19984
rect 16301 19935 16359 19941
rect 19352 19944 20076 19972
rect 11146 19904 11152 19916
rect 6012 19876 8340 19904
rect 11107 19876 11152 19904
rect 7098 19836 7104 19848
rect 5592 19808 5637 19836
rect 5920 19808 7104 19836
rect 5592 19796 5598 19808
rect 7098 19796 7104 19808
rect 7156 19796 7162 19848
rect 7392 19845 7420 19876
rect 11146 19864 11152 19876
rect 11204 19864 11210 19916
rect 11974 19904 11980 19916
rect 11935 19876 11980 19904
rect 11974 19864 11980 19876
rect 12032 19864 12038 19916
rect 14108 19876 14872 19904
rect 7377 19839 7435 19845
rect 7377 19805 7389 19839
rect 7423 19805 7435 19839
rect 7377 19799 7435 19805
rect 7834 19796 7840 19848
rect 7892 19836 7898 19848
rect 9674 19836 9680 19848
rect 7892 19808 8156 19836
rect 9635 19808 9680 19836
rect 7892 19796 7898 19808
rect 3053 19771 3111 19777
rect 3053 19737 3065 19771
rect 3099 19737 3111 19771
rect 8018 19768 8024 19780
rect 3053 19731 3111 19737
rect 6104 19740 8024 19768
rect 4893 19703 4951 19709
rect 4893 19669 4905 19703
rect 4939 19700 4951 19703
rect 6104 19700 6132 19740
rect 8018 19728 8024 19740
rect 8076 19728 8082 19780
rect 8128 19768 8156 19808
rect 9674 19796 9680 19808
rect 9732 19796 9738 19848
rect 11057 19839 11115 19845
rect 11057 19805 11069 19839
rect 11103 19836 11115 19839
rect 11992 19836 12020 19864
rect 14108 19845 14136 19876
rect 11103 19808 12020 19836
rect 14093 19839 14151 19845
rect 11103 19805 11115 19808
rect 11057 19799 11115 19805
rect 14093 19805 14105 19839
rect 14139 19805 14151 19839
rect 14093 19799 14151 19805
rect 14277 19839 14335 19845
rect 14277 19805 14289 19839
rect 14323 19805 14335 19839
rect 14277 19799 14335 19805
rect 8221 19771 8279 19777
rect 8221 19768 8233 19771
rect 8128 19740 8233 19768
rect 8221 19737 8233 19740
rect 8267 19737 8279 19771
rect 9490 19768 9496 19780
rect 9403 19740 9496 19768
rect 8221 19731 8279 19737
rect 9490 19728 9496 19740
rect 9548 19728 9554 19780
rect 10045 19771 10103 19777
rect 10045 19737 10057 19771
rect 10091 19768 10103 19771
rect 10226 19768 10232 19780
rect 10091 19740 10232 19768
rect 10091 19737 10103 19740
rect 10045 19731 10103 19737
rect 10226 19728 10232 19740
rect 10284 19728 10290 19780
rect 13630 19728 13636 19780
rect 13688 19768 13694 19780
rect 14292 19768 14320 19799
rect 13688 19740 14320 19768
rect 13688 19728 13694 19740
rect 6270 19700 6276 19712
rect 4939 19672 6132 19700
rect 6231 19672 6276 19700
rect 4939 19669 4951 19672
rect 4893 19663 4951 19669
rect 6270 19660 6276 19672
rect 6328 19660 6334 19712
rect 7561 19703 7619 19709
rect 7561 19669 7573 19703
rect 7607 19700 7619 19703
rect 7834 19700 7840 19712
rect 7607 19672 7840 19700
rect 7607 19669 7619 19672
rect 7561 19663 7619 19669
rect 7834 19660 7840 19672
rect 7892 19660 7898 19712
rect 8389 19703 8447 19709
rect 8389 19669 8401 19703
rect 8435 19700 8447 19703
rect 9508 19700 9536 19728
rect 14182 19700 14188 19712
rect 8435 19672 9536 19700
rect 14143 19672 14188 19700
rect 8435 19669 8447 19672
rect 8389 19663 8447 19669
rect 14182 19660 14188 19672
rect 14240 19660 14246 19712
rect 14844 19709 14872 19876
rect 16316 19836 16344 19935
rect 19352 19913 19380 19944
rect 20070 19932 20076 19944
rect 20128 19932 20134 19984
rect 16485 19907 16543 19913
rect 16485 19873 16497 19907
rect 16531 19904 16543 19907
rect 19337 19907 19395 19913
rect 19337 19904 19349 19907
rect 16531 19876 19349 19904
rect 16531 19873 16543 19876
rect 16485 19867 16543 19873
rect 19337 19873 19349 19876
rect 19383 19873 19395 19907
rect 19337 19867 19395 19873
rect 19978 19864 19984 19916
rect 20036 19904 20042 19916
rect 26804 19904 26832 20012
rect 27433 19975 27491 19981
rect 27433 19941 27445 19975
rect 27479 19972 27491 19975
rect 34072 19972 34100 20012
rect 34149 20009 34161 20043
rect 34195 20040 34207 20043
rect 34514 20040 34520 20052
rect 34195 20012 34520 20040
rect 34195 20009 34207 20012
rect 34149 20003 34207 20009
rect 34514 20000 34520 20012
rect 34572 20000 34578 20052
rect 42794 20000 42800 20052
rect 42852 20040 42858 20052
rect 43165 20043 43223 20049
rect 43165 20040 43177 20043
rect 42852 20012 43177 20040
rect 42852 20000 42858 20012
rect 43165 20009 43177 20012
rect 43211 20009 43223 20043
rect 43165 20003 43223 20009
rect 53929 20043 53987 20049
rect 53929 20009 53941 20043
rect 53975 20040 53987 20043
rect 54202 20040 54208 20052
rect 53975 20012 54208 20040
rect 53975 20009 53987 20012
rect 53929 20003 53987 20009
rect 54202 20000 54208 20012
rect 54260 20000 54266 20052
rect 54386 20040 54392 20052
rect 54347 20012 54392 20040
rect 54386 20000 54392 20012
rect 54444 20000 54450 20052
rect 39758 19972 39764 19984
rect 27479 19944 31754 19972
rect 34072 19944 39764 19972
rect 27479 19941 27491 19944
rect 27433 19935 27491 19941
rect 28994 19904 29000 19916
rect 20036 19876 26832 19904
rect 28184 19876 29000 19904
rect 20036 19864 20042 19876
rect 17037 19839 17095 19845
rect 17037 19836 17049 19839
rect 16316 19808 17049 19836
rect 17037 19805 17049 19808
rect 17083 19805 17095 19839
rect 17037 19799 17095 19805
rect 18690 19796 18696 19848
rect 18748 19836 18754 19848
rect 19613 19839 19671 19845
rect 19613 19836 19625 19839
rect 18748 19808 19625 19836
rect 18748 19796 18754 19808
rect 16022 19768 16028 19780
rect 15983 19740 16028 19768
rect 16022 19728 16028 19740
rect 16080 19728 16086 19780
rect 17221 19771 17279 19777
rect 17221 19737 17233 19771
rect 17267 19768 17279 19771
rect 17770 19768 17776 19780
rect 17267 19740 17776 19768
rect 17267 19737 17279 19740
rect 17221 19731 17279 19737
rect 17770 19728 17776 19740
rect 17828 19728 17834 19780
rect 14829 19703 14887 19709
rect 14829 19669 14841 19703
rect 14875 19700 14887 19703
rect 18230 19700 18236 19712
rect 14875 19672 18236 19700
rect 14875 19669 14887 19672
rect 14829 19663 14887 19669
rect 18230 19660 18236 19672
rect 18288 19660 18294 19712
rect 19168 19700 19196 19808
rect 19613 19805 19625 19808
rect 19659 19805 19671 19839
rect 26326 19836 26332 19848
rect 19613 19799 19671 19805
rect 19720 19808 26332 19836
rect 19242 19728 19248 19780
rect 19300 19768 19306 19780
rect 19720 19768 19748 19808
rect 26326 19796 26332 19808
rect 26384 19796 26390 19848
rect 26510 19796 26516 19848
rect 26568 19836 26574 19848
rect 27154 19836 27160 19848
rect 26568 19808 27160 19836
rect 26568 19796 26574 19808
rect 27154 19796 27160 19808
rect 27212 19796 27218 19848
rect 28074 19836 28080 19848
rect 28035 19808 28080 19836
rect 28074 19796 28080 19808
rect 28132 19796 28138 19848
rect 28184 19780 28212 19876
rect 28994 19864 29000 19876
rect 29052 19864 29058 19916
rect 30834 19904 30840 19916
rect 30795 19876 30840 19904
rect 30834 19864 30840 19876
rect 30892 19864 30898 19916
rect 31726 19904 31754 19944
rect 39758 19932 39764 19944
rect 39816 19932 39822 19984
rect 33502 19904 33508 19916
rect 31726 19876 33508 19904
rect 33502 19864 33508 19876
rect 33560 19904 33566 19916
rect 38286 19904 38292 19916
rect 33560 19876 33916 19904
rect 38247 19876 38292 19904
rect 33560 19864 33566 19876
rect 28258 19796 28264 19848
rect 28316 19836 28322 19848
rect 28445 19839 28503 19845
rect 28316 19808 28361 19836
rect 28316 19796 28322 19808
rect 28445 19805 28457 19839
rect 28491 19836 28503 19839
rect 28810 19836 28816 19848
rect 28491 19808 28816 19836
rect 28491 19805 28503 19808
rect 28445 19799 28503 19805
rect 28810 19796 28816 19808
rect 28868 19836 28874 19848
rect 33888 19845 33916 19876
rect 38286 19864 38292 19876
rect 38344 19864 38350 19916
rect 38657 19907 38715 19913
rect 38657 19873 38669 19907
rect 38703 19904 38715 19907
rect 43438 19904 43444 19916
rect 38703 19876 43444 19904
rect 38703 19873 38715 19876
rect 38657 19867 38715 19873
rect 43438 19864 43444 19876
rect 43496 19864 43502 19916
rect 46753 19907 46811 19913
rect 46753 19873 46765 19907
rect 46799 19904 46811 19907
rect 46934 19904 46940 19916
rect 46799 19876 46940 19904
rect 46799 19873 46811 19876
rect 46753 19867 46811 19873
rect 46934 19864 46940 19876
rect 46992 19864 46998 19916
rect 47581 19907 47639 19913
rect 47581 19873 47593 19907
rect 47627 19904 47639 19907
rect 48314 19904 48320 19916
rect 47627 19876 48320 19904
rect 47627 19873 47639 19876
rect 47581 19867 47639 19873
rect 48314 19864 48320 19876
rect 48372 19864 48378 19916
rect 48958 19864 48964 19916
rect 49016 19904 49022 19916
rect 56781 19907 56839 19913
rect 49016 19876 53788 19904
rect 49016 19864 49022 19876
rect 28905 19839 28963 19845
rect 28905 19836 28917 19839
rect 28868 19808 28917 19836
rect 28868 19796 28874 19808
rect 28905 19805 28917 19808
rect 28951 19805 28963 19839
rect 28905 19799 28963 19805
rect 33873 19839 33931 19845
rect 33873 19805 33885 19839
rect 33919 19805 33931 19839
rect 33873 19799 33931 19805
rect 34149 19839 34207 19845
rect 34149 19805 34161 19839
rect 34195 19805 34207 19839
rect 34149 19799 34207 19805
rect 19300 19740 19748 19768
rect 19300 19728 19306 19740
rect 20898 19728 20904 19780
rect 20956 19768 20962 19780
rect 23293 19771 23351 19777
rect 23293 19768 23305 19771
rect 20956 19740 23305 19768
rect 20956 19728 20962 19740
rect 23293 19737 23305 19740
rect 23339 19737 23351 19771
rect 23293 19731 23351 19737
rect 25958 19728 25964 19780
rect 26016 19768 26022 19780
rect 27249 19771 27307 19777
rect 27249 19768 27261 19771
rect 26016 19740 27261 19768
rect 26016 19728 26022 19740
rect 27249 19737 27261 19740
rect 27295 19737 27307 19771
rect 27249 19731 27307 19737
rect 27433 19771 27491 19777
rect 27433 19737 27445 19771
rect 27479 19737 27491 19771
rect 28166 19768 28172 19780
rect 28127 19740 28172 19768
rect 27433 19731 27491 19737
rect 20070 19700 20076 19712
rect 19168 19672 20076 19700
rect 20070 19660 20076 19672
rect 20128 19660 20134 19712
rect 20990 19660 20996 19712
rect 21048 19700 21054 19712
rect 21637 19703 21695 19709
rect 21637 19700 21649 19703
rect 21048 19672 21649 19700
rect 21048 19660 21054 19672
rect 21637 19669 21649 19672
rect 21683 19700 21695 19703
rect 22186 19700 22192 19712
rect 21683 19672 22192 19700
rect 21683 19669 21695 19672
rect 21637 19663 21695 19669
rect 22186 19660 22192 19672
rect 22244 19660 22250 19712
rect 23198 19700 23204 19712
rect 23159 19672 23204 19700
rect 23198 19660 23204 19672
rect 23256 19660 23262 19712
rect 27448 19700 27476 19731
rect 28166 19728 28172 19740
rect 28224 19728 28230 19780
rect 27893 19703 27951 19709
rect 27893 19700 27905 19703
rect 27448 19672 27905 19700
rect 27893 19669 27905 19672
rect 27939 19669 27951 19703
rect 28276 19700 28304 19796
rect 29638 19728 29644 19780
rect 29696 19768 29702 19780
rect 31846 19768 31852 19780
rect 29696 19740 31852 19768
rect 29696 19728 29702 19740
rect 31846 19728 31852 19740
rect 31904 19768 31910 19780
rect 32217 19771 32275 19777
rect 32217 19768 32229 19771
rect 31904 19740 32229 19768
rect 31904 19728 31910 19740
rect 32217 19737 32229 19740
rect 32263 19737 32275 19771
rect 32217 19731 32275 19737
rect 32401 19771 32459 19777
rect 32401 19737 32413 19771
rect 32447 19768 32459 19771
rect 32858 19768 32864 19780
rect 32447 19740 32864 19768
rect 32447 19737 32459 19740
rect 32401 19731 32459 19737
rect 32858 19728 32864 19740
rect 32916 19728 32922 19780
rect 33410 19728 33416 19780
rect 33468 19768 33474 19780
rect 34057 19771 34115 19777
rect 34057 19768 34069 19771
rect 33468 19740 34069 19768
rect 33468 19728 33474 19740
rect 34057 19737 34069 19740
rect 34103 19737 34115 19771
rect 34164 19768 34192 19799
rect 34790 19796 34796 19848
rect 34848 19836 34854 19848
rect 34977 19839 35035 19845
rect 34977 19836 34989 19839
rect 34848 19808 34989 19836
rect 34848 19796 34854 19808
rect 34977 19805 34989 19808
rect 35023 19805 35035 19839
rect 35986 19836 35992 19848
rect 35947 19808 35992 19836
rect 34977 19799 35035 19805
rect 35986 19796 35992 19808
rect 36044 19796 36050 19848
rect 36170 19836 36176 19848
rect 36131 19808 36176 19836
rect 36170 19796 36176 19808
rect 36228 19796 36234 19848
rect 37001 19839 37059 19845
rect 37001 19805 37013 19839
rect 37047 19836 37059 19839
rect 38470 19836 38476 19848
rect 37047 19808 38476 19836
rect 37047 19805 37059 19808
rect 37001 19799 37059 19805
rect 38470 19796 38476 19808
rect 38528 19796 38534 19848
rect 44174 19796 44180 19848
rect 44232 19836 44238 19848
rect 47762 19836 47768 19848
rect 44232 19808 45554 19836
rect 47242 19822 47768 19836
rect 44232 19796 44238 19808
rect 34164 19740 34836 19768
rect 34057 19731 34115 19737
rect 29914 19700 29920 19712
rect 28276 19672 29920 19700
rect 27893 19663 27951 19669
rect 29914 19660 29920 19672
rect 29972 19660 29978 19712
rect 34808 19709 34836 19740
rect 42702 19728 42708 19780
rect 42760 19768 42766 19780
rect 42981 19771 43039 19777
rect 42981 19768 42993 19771
rect 42760 19740 42993 19768
rect 42760 19728 42766 19740
rect 42981 19737 42993 19740
rect 43027 19737 43039 19771
rect 45526 19768 45554 19808
rect 47228 19808 47768 19822
rect 47228 19768 47256 19808
rect 47762 19796 47768 19808
rect 47820 19796 47826 19848
rect 49878 19796 49884 19848
rect 49936 19836 49942 19848
rect 50157 19839 50215 19845
rect 50157 19836 50169 19839
rect 49936 19808 50169 19836
rect 49936 19796 49942 19808
rect 50157 19805 50169 19808
rect 50203 19805 50215 19839
rect 50157 19799 50215 19805
rect 50525 19839 50583 19845
rect 50525 19805 50537 19839
rect 50571 19836 50583 19839
rect 50614 19836 50620 19848
rect 50571 19808 50620 19836
rect 50571 19805 50583 19808
rect 50525 19799 50583 19805
rect 45526 19740 47256 19768
rect 50172 19768 50200 19799
rect 50614 19796 50620 19808
rect 50672 19796 50678 19848
rect 50706 19796 50712 19848
rect 50764 19836 50770 19848
rect 53466 19836 53472 19848
rect 50764 19808 50809 19836
rect 53427 19808 53472 19836
rect 50764 19796 50770 19808
rect 53466 19796 53472 19808
rect 53524 19796 53530 19848
rect 53760 19845 53788 19876
rect 56781 19873 56793 19907
rect 56827 19904 56839 19907
rect 57330 19904 57336 19916
rect 56827 19876 57336 19904
rect 56827 19873 56839 19876
rect 56781 19867 56839 19873
rect 57330 19864 57336 19876
rect 57388 19864 57394 19916
rect 53745 19839 53803 19845
rect 53745 19805 53757 19839
rect 53791 19836 53803 19839
rect 53926 19836 53932 19848
rect 53791 19808 53932 19836
rect 53791 19805 53803 19808
rect 53745 19799 53803 19805
rect 53926 19796 53932 19808
rect 53984 19836 53990 19848
rect 54389 19839 54447 19845
rect 54389 19836 54401 19839
rect 53984 19808 54401 19836
rect 53984 19796 53990 19808
rect 54389 19805 54401 19808
rect 54435 19805 54447 19839
rect 56686 19836 56692 19848
rect 56647 19808 56692 19836
rect 54389 19799 54447 19805
rect 56686 19796 56692 19808
rect 56744 19796 56750 19848
rect 56870 19836 56876 19848
rect 56831 19808 56876 19836
rect 56870 19796 56876 19808
rect 56928 19796 56934 19848
rect 56965 19839 57023 19845
rect 56965 19805 56977 19839
rect 57011 19836 57023 19839
rect 57146 19836 57152 19848
rect 57011 19808 57152 19836
rect 57011 19805 57023 19808
rect 56965 19799 57023 19805
rect 57146 19796 57152 19808
rect 57204 19796 57210 19848
rect 50982 19768 50988 19780
rect 50172 19740 50988 19768
rect 42981 19731 43039 19737
rect 50982 19728 50988 19740
rect 51040 19728 51046 19780
rect 54481 19771 54539 19777
rect 54481 19737 54493 19771
rect 54527 19737 54539 19771
rect 54662 19768 54668 19780
rect 54623 19740 54668 19768
rect 54481 19731 54539 19737
rect 34793 19703 34851 19709
rect 34793 19669 34805 19703
rect 34839 19700 34851 19703
rect 38838 19700 38844 19712
rect 34839 19672 38844 19700
rect 34839 19669 34851 19672
rect 34793 19663 34851 19669
rect 38838 19660 38844 19672
rect 38896 19660 38902 19712
rect 41782 19660 41788 19712
rect 41840 19700 41846 19712
rect 42429 19703 42487 19709
rect 42429 19700 42441 19703
rect 41840 19672 42441 19700
rect 41840 19660 41846 19672
rect 42429 19669 42441 19672
rect 42475 19700 42487 19703
rect 43181 19703 43239 19709
rect 43181 19700 43193 19703
rect 42475 19672 43193 19700
rect 42475 19669 42487 19672
rect 42429 19663 42487 19669
rect 43181 19669 43193 19672
rect 43227 19669 43239 19703
rect 43181 19663 43239 19669
rect 43349 19703 43407 19709
rect 43349 19669 43361 19703
rect 43395 19700 43407 19703
rect 48774 19700 48780 19712
rect 43395 19672 48780 19700
rect 43395 19669 43407 19672
rect 43349 19663 43407 19669
rect 48774 19660 48780 19672
rect 48832 19660 48838 19712
rect 50525 19703 50583 19709
rect 50525 19669 50537 19703
rect 50571 19700 50583 19703
rect 51994 19700 52000 19712
rect 50571 19672 52000 19700
rect 50571 19669 50583 19672
rect 50525 19663 50583 19669
rect 51994 19660 52000 19672
rect 52052 19660 52058 19712
rect 53558 19700 53564 19712
rect 53519 19672 53564 19700
rect 53558 19660 53564 19672
rect 53616 19700 53622 19712
rect 54496 19700 54524 19731
rect 54662 19728 54668 19740
rect 54720 19728 54726 19780
rect 56502 19700 56508 19712
rect 53616 19672 54524 19700
rect 56463 19672 56508 19700
rect 53616 19660 53622 19672
rect 56502 19660 56508 19672
rect 56560 19660 56566 19712
rect 1104 19610 58880 19632
rect 1104 19558 19574 19610
rect 19626 19558 19638 19610
rect 19690 19558 19702 19610
rect 19754 19558 19766 19610
rect 19818 19558 19830 19610
rect 19882 19558 50294 19610
rect 50346 19558 50358 19610
rect 50410 19558 50422 19610
rect 50474 19558 50486 19610
rect 50538 19558 50550 19610
rect 50602 19558 58880 19610
rect 1104 19536 58880 19558
rect 2866 19456 2872 19508
rect 2924 19496 2930 19508
rect 4985 19499 5043 19505
rect 4985 19496 4997 19499
rect 2924 19468 4997 19496
rect 2924 19456 2930 19468
rect 1394 19320 1400 19372
rect 1452 19360 1458 19372
rect 3344 19369 3372 19468
rect 4985 19465 4997 19468
rect 5031 19496 5043 19499
rect 5442 19496 5448 19508
rect 5031 19468 5448 19496
rect 5031 19465 5043 19468
rect 4985 19459 5043 19465
rect 5442 19456 5448 19468
rect 5500 19456 5506 19508
rect 13357 19499 13415 19505
rect 13357 19465 13369 19499
rect 13403 19496 13415 19499
rect 14366 19496 14372 19508
rect 13403 19468 14372 19496
rect 13403 19465 13415 19468
rect 13357 19459 13415 19465
rect 14366 19456 14372 19468
rect 14424 19456 14430 19508
rect 17773 19499 17831 19505
rect 17773 19465 17785 19499
rect 17819 19496 17831 19499
rect 18598 19496 18604 19508
rect 17819 19468 18604 19496
rect 17819 19465 17831 19468
rect 17773 19459 17831 19465
rect 18598 19456 18604 19468
rect 18656 19456 18662 19508
rect 18785 19499 18843 19505
rect 18785 19465 18797 19499
rect 18831 19465 18843 19499
rect 18785 19459 18843 19465
rect 7742 19428 7748 19440
rect 7208 19400 7748 19428
rect 7208 19372 7236 19400
rect 7742 19388 7748 19400
rect 7800 19388 7806 19440
rect 9950 19388 9956 19440
rect 10008 19428 10014 19440
rect 12529 19431 12587 19437
rect 12529 19428 12541 19431
rect 10008 19400 12541 19428
rect 10008 19388 10014 19400
rect 12529 19397 12541 19400
rect 12575 19397 12587 19431
rect 12529 19391 12587 19397
rect 14182 19388 14188 19440
rect 14240 19428 14246 19440
rect 15930 19428 15936 19440
rect 14240 19400 15148 19428
rect 15891 19400 15936 19428
rect 14240 19388 14246 19400
rect 1489 19363 1547 19369
rect 1489 19360 1501 19363
rect 1452 19332 1501 19360
rect 1452 19320 1458 19332
rect 1489 19329 1501 19332
rect 1535 19329 1547 19363
rect 1489 19323 1547 19329
rect 3329 19363 3387 19369
rect 3329 19329 3341 19363
rect 3375 19329 3387 19363
rect 3329 19323 3387 19329
rect 3697 19363 3755 19369
rect 3697 19329 3709 19363
rect 3743 19329 3755 19363
rect 3697 19323 3755 19329
rect 5077 19363 5135 19369
rect 5077 19329 5089 19363
rect 5123 19360 5135 19363
rect 5534 19360 5540 19372
rect 5123 19332 5540 19360
rect 5123 19329 5135 19332
rect 5077 19323 5135 19329
rect 3712 19292 3740 19323
rect 5534 19320 5540 19332
rect 5592 19360 5598 19372
rect 5721 19363 5779 19369
rect 5721 19360 5733 19363
rect 5592 19332 5733 19360
rect 5592 19320 5598 19332
rect 5721 19329 5733 19332
rect 5767 19360 5779 19363
rect 6270 19360 6276 19372
rect 5767 19332 6276 19360
rect 5767 19329 5779 19332
rect 5721 19323 5779 19329
rect 6270 19320 6276 19332
rect 6328 19320 6334 19372
rect 7190 19360 7196 19372
rect 7103 19332 7196 19360
rect 7190 19320 7196 19332
rect 7248 19320 7254 19372
rect 7466 19360 7472 19372
rect 7427 19332 7472 19360
rect 7466 19320 7472 19332
rect 7524 19320 7530 19372
rect 7929 19363 7987 19369
rect 7929 19329 7941 19363
rect 7975 19360 7987 19363
rect 8018 19360 8024 19372
rect 7975 19332 8024 19360
rect 7975 19329 7987 19332
rect 7929 19323 7987 19329
rect 8018 19320 8024 19332
rect 8076 19320 8082 19372
rect 13630 19360 13636 19372
rect 13591 19332 13636 19360
rect 13630 19320 13636 19332
rect 13688 19320 13694 19372
rect 13909 19363 13967 19369
rect 13909 19329 13921 19363
rect 13955 19360 13967 19363
rect 14642 19360 14648 19372
rect 13955 19332 14648 19360
rect 13955 19329 13967 19332
rect 13909 19323 13967 19329
rect 14642 19320 14648 19332
rect 14700 19320 14706 19372
rect 14826 19360 14832 19372
rect 14787 19332 14832 19360
rect 14826 19320 14832 19332
rect 14884 19320 14890 19372
rect 15120 19369 15148 19400
rect 15930 19388 15936 19400
rect 15988 19388 15994 19440
rect 18046 19388 18052 19440
rect 18104 19428 18110 19440
rect 18506 19428 18512 19440
rect 18104 19400 18368 19428
rect 18467 19400 18512 19428
rect 18104 19388 18110 19400
rect 15105 19363 15163 19369
rect 15105 19329 15117 19363
rect 15151 19329 15163 19363
rect 15105 19323 15163 19329
rect 15194 19320 15200 19372
rect 15252 19360 15258 19372
rect 15473 19363 15531 19369
rect 15252 19332 15297 19360
rect 15252 19320 15258 19332
rect 15473 19329 15485 19363
rect 15519 19329 15531 19363
rect 15473 19323 15531 19329
rect 3970 19292 3976 19304
rect 3712 19264 3976 19292
rect 3970 19252 3976 19264
rect 4028 19292 4034 19304
rect 6914 19292 6920 19304
rect 4028 19264 6920 19292
rect 4028 19252 4034 19264
rect 6914 19252 6920 19264
rect 6972 19252 6978 19304
rect 7742 19292 7748 19304
rect 7703 19264 7748 19292
rect 7742 19252 7748 19264
rect 7800 19252 7806 19304
rect 10781 19295 10839 19301
rect 10781 19261 10793 19295
rect 10827 19292 10839 19295
rect 11146 19292 11152 19304
rect 10827 19264 11152 19292
rect 10827 19261 10839 19264
rect 10781 19255 10839 19261
rect 11146 19252 11152 19264
rect 11204 19252 11210 19304
rect 13538 19292 13544 19304
rect 13499 19264 13544 19292
rect 13538 19252 13544 19264
rect 13596 19252 13602 19304
rect 14001 19295 14059 19301
rect 14001 19261 14013 19295
rect 14047 19292 14059 19295
rect 14734 19292 14740 19304
rect 14047 19264 14740 19292
rect 14047 19261 14059 19264
rect 14001 19255 14059 19261
rect 14734 19252 14740 19264
rect 14792 19252 14798 19304
rect 15488 19292 15516 19323
rect 16022 19320 16028 19372
rect 16080 19360 16086 19372
rect 17589 19363 17647 19369
rect 17589 19360 17601 19363
rect 16080 19332 17601 19360
rect 16080 19320 16086 19332
rect 17589 19329 17601 19332
rect 17635 19329 17647 19363
rect 17770 19360 17776 19372
rect 17731 19332 17776 19360
rect 17589 19323 17647 19329
rect 17770 19320 17776 19332
rect 17828 19320 17834 19372
rect 18230 19360 18236 19372
rect 18191 19332 18236 19360
rect 18230 19320 18236 19332
rect 18288 19320 18294 19372
rect 18340 19360 18368 19400
rect 18506 19388 18512 19400
rect 18564 19388 18570 19440
rect 18417 19363 18475 19369
rect 18417 19360 18429 19363
rect 18340 19332 18429 19360
rect 18417 19329 18429 19332
rect 18463 19329 18475 19363
rect 18417 19323 18475 19329
rect 18601 19363 18659 19369
rect 18601 19329 18613 19363
rect 18647 19360 18659 19363
rect 18690 19360 18696 19372
rect 18647 19332 18696 19360
rect 18647 19329 18659 19332
rect 18601 19323 18659 19329
rect 18690 19320 18696 19332
rect 18748 19320 18754 19372
rect 18800 19360 18828 19459
rect 18874 19456 18880 19508
rect 18932 19496 18938 19508
rect 19889 19499 19947 19505
rect 18932 19468 19656 19496
rect 18932 19456 18938 19468
rect 19150 19388 19156 19440
rect 19208 19428 19214 19440
rect 19208 19400 19380 19428
rect 19208 19388 19214 19400
rect 19352 19369 19380 19400
rect 19245 19363 19303 19369
rect 19245 19360 19257 19363
rect 18800 19332 19257 19360
rect 19245 19329 19257 19332
rect 19291 19329 19303 19363
rect 19245 19323 19303 19329
rect 19338 19363 19396 19369
rect 19338 19329 19350 19363
rect 19384 19329 19396 19363
rect 19518 19360 19524 19372
rect 19479 19332 19524 19360
rect 19338 19323 19396 19329
rect 19518 19320 19524 19332
rect 19576 19320 19582 19372
rect 19628 19369 19656 19468
rect 19889 19465 19901 19499
rect 19935 19496 19947 19499
rect 19978 19496 19984 19508
rect 19935 19468 19984 19496
rect 19935 19465 19947 19468
rect 19889 19459 19947 19465
rect 19978 19456 19984 19468
rect 20036 19456 20042 19508
rect 22370 19496 22376 19508
rect 21836 19468 22376 19496
rect 21450 19388 21456 19440
rect 21508 19428 21514 19440
rect 21508 19400 21772 19428
rect 21508 19388 21514 19400
rect 19613 19363 19671 19369
rect 19613 19329 19625 19363
rect 19659 19329 19671 19363
rect 19613 19323 19671 19329
rect 16206 19292 16212 19304
rect 15488 19264 16212 19292
rect 16206 19252 16212 19264
rect 16264 19252 16270 19304
rect 16758 19292 16764 19304
rect 16719 19264 16764 19292
rect 16758 19252 16764 19264
rect 16816 19252 16822 19304
rect 19628 19292 19656 19323
rect 19702 19320 19708 19372
rect 19760 19369 19766 19372
rect 19760 19360 19768 19369
rect 21085 19363 21143 19369
rect 19760 19332 19805 19360
rect 19760 19323 19768 19332
rect 21085 19329 21097 19363
rect 21131 19329 21143 19363
rect 21085 19323 21143 19329
rect 19760 19320 19766 19323
rect 19978 19292 19984 19304
rect 19628 19264 19984 19292
rect 19978 19252 19984 19264
rect 20036 19292 20042 19304
rect 20441 19295 20499 19301
rect 20441 19292 20453 19295
rect 20036 19264 20453 19292
rect 20036 19252 20042 19264
rect 20441 19261 20453 19264
rect 20487 19261 20499 19295
rect 20441 19255 20499 19261
rect 21100 19292 21128 19323
rect 21450 19292 21456 19304
rect 21100 19264 21456 19292
rect 7650 19184 7656 19236
rect 7708 19224 7714 19236
rect 7837 19227 7895 19233
rect 7837 19224 7849 19227
rect 7708 19196 7849 19224
rect 7708 19184 7714 19196
rect 7837 19193 7849 19196
rect 7883 19193 7895 19227
rect 7837 19187 7895 19193
rect 10502 19184 10508 19236
rect 10560 19224 10566 19236
rect 10560 19196 16160 19224
rect 10560 19184 10566 19196
rect 16132 19168 16160 19196
rect 16390 19184 16396 19236
rect 16448 19224 16454 19236
rect 21100 19224 21128 19264
rect 21450 19252 21456 19264
rect 21508 19252 21514 19304
rect 21744 19292 21772 19400
rect 21836 19369 21864 19468
rect 22370 19456 22376 19468
rect 22428 19456 22434 19508
rect 22465 19499 22523 19505
rect 22465 19465 22477 19499
rect 22511 19496 22523 19499
rect 23382 19496 23388 19508
rect 22511 19468 23388 19496
rect 22511 19465 22523 19468
rect 22465 19459 22523 19465
rect 23382 19456 23388 19468
rect 23440 19456 23446 19508
rect 24029 19499 24087 19505
rect 24029 19465 24041 19499
rect 24075 19465 24087 19499
rect 24946 19496 24952 19508
rect 24029 19459 24087 19465
rect 24228 19468 24952 19496
rect 22094 19428 22100 19440
rect 22055 19400 22100 19428
rect 22094 19388 22100 19400
rect 22152 19428 22158 19440
rect 22738 19428 22744 19440
rect 22152 19400 22744 19428
rect 22152 19388 22158 19400
rect 22738 19388 22744 19400
rect 22796 19388 22802 19440
rect 21827 19363 21885 19369
rect 21827 19329 21839 19363
rect 21873 19329 21885 19363
rect 21827 19323 21885 19329
rect 21914 19363 21972 19369
rect 21914 19329 21926 19363
rect 21960 19360 21972 19363
rect 22186 19360 22192 19372
rect 21960 19332 21993 19360
rect 22147 19332 22192 19360
rect 21960 19329 21972 19332
rect 21914 19323 21972 19329
rect 21928 19292 21956 19323
rect 22186 19320 22192 19332
rect 22244 19320 22250 19372
rect 22286 19363 22344 19369
rect 22286 19329 22298 19363
rect 22332 19329 22344 19363
rect 22286 19323 22344 19329
rect 21744 19264 21956 19292
rect 16448 19196 21128 19224
rect 16448 19184 16454 19196
rect 21910 19184 21916 19236
rect 21968 19224 21974 19236
rect 22296 19224 22324 19323
rect 23014 19320 23020 19372
rect 23072 19360 23078 19372
rect 23201 19363 23259 19369
rect 23201 19360 23213 19363
rect 23072 19332 23213 19360
rect 23072 19320 23078 19332
rect 23201 19329 23213 19332
rect 23247 19329 23259 19363
rect 23201 19323 23259 19329
rect 23290 19320 23296 19372
rect 23348 19360 23354 19372
rect 23474 19360 23480 19372
rect 23348 19332 23393 19360
rect 23435 19332 23480 19360
rect 23348 19320 23354 19332
rect 23474 19320 23480 19332
rect 23532 19320 23538 19372
rect 23569 19363 23627 19369
rect 23569 19329 23581 19363
rect 23615 19360 23627 19363
rect 24044 19360 24072 19459
rect 24228 19369 24256 19468
rect 24946 19456 24952 19468
rect 25004 19456 25010 19508
rect 28074 19456 28080 19508
rect 28132 19496 28138 19508
rect 29730 19496 29736 19508
rect 28132 19468 29736 19496
rect 28132 19456 28138 19468
rect 29730 19456 29736 19468
rect 29788 19456 29794 19508
rect 32674 19496 32680 19508
rect 32635 19468 32680 19496
rect 32674 19456 32680 19468
rect 32732 19456 32738 19508
rect 34790 19456 34796 19508
rect 34848 19496 34854 19508
rect 35069 19499 35127 19505
rect 35069 19496 35081 19499
rect 34848 19468 35081 19496
rect 34848 19456 34854 19468
rect 35069 19465 35081 19468
rect 35115 19465 35127 19499
rect 44174 19496 44180 19508
rect 44135 19468 44180 19496
rect 35069 19459 35127 19465
rect 44174 19456 44180 19468
rect 44232 19456 44238 19508
rect 50614 19456 50620 19508
rect 50672 19496 50678 19508
rect 50801 19499 50859 19505
rect 50801 19496 50813 19499
rect 50672 19468 50813 19496
rect 50672 19456 50678 19468
rect 50801 19465 50813 19468
rect 50847 19465 50859 19499
rect 50801 19459 50859 19465
rect 24305 19431 24363 19437
rect 24305 19397 24317 19431
rect 24351 19428 24363 19431
rect 24670 19428 24676 19440
rect 24351 19400 24676 19428
rect 24351 19397 24363 19400
rect 24305 19391 24363 19397
rect 24670 19388 24676 19400
rect 24728 19388 24734 19440
rect 28994 19388 29000 19440
rect 29052 19428 29058 19440
rect 35986 19428 35992 19440
rect 29052 19400 35992 19428
rect 29052 19388 29058 19400
rect 35986 19388 35992 19400
rect 36044 19388 36050 19440
rect 43257 19431 43315 19437
rect 43257 19397 43269 19431
rect 43303 19428 43315 19431
rect 47949 19431 48007 19437
rect 43303 19400 47900 19428
rect 43303 19397 43315 19400
rect 43257 19391 43315 19397
rect 23615 19332 24072 19360
rect 24213 19363 24271 19369
rect 23615 19329 23627 19332
rect 23569 19323 23627 19329
rect 24213 19329 24225 19363
rect 24259 19329 24271 19363
rect 24213 19323 24271 19329
rect 24397 19363 24455 19369
rect 24397 19329 24409 19363
rect 24443 19360 24455 19363
rect 24486 19360 24492 19372
rect 24443 19332 24492 19360
rect 24443 19329 24455 19332
rect 24397 19323 24455 19329
rect 24486 19320 24492 19332
rect 24544 19320 24550 19372
rect 24581 19363 24639 19369
rect 24581 19329 24593 19363
rect 24627 19360 24639 19363
rect 24762 19360 24768 19372
rect 24627 19332 24768 19360
rect 24627 19329 24639 19332
rect 24581 19323 24639 19329
rect 24762 19320 24768 19332
rect 24820 19320 24826 19372
rect 28261 19363 28319 19369
rect 28261 19329 28273 19363
rect 28307 19360 28319 19363
rect 31389 19363 31447 19369
rect 31389 19360 31401 19363
rect 28307 19332 31401 19360
rect 28307 19329 28319 19332
rect 28261 19323 28319 19329
rect 31389 19329 31401 19332
rect 31435 19360 31447 19363
rect 31754 19360 31760 19372
rect 31435 19332 31760 19360
rect 31435 19329 31447 19332
rect 31389 19323 31447 19329
rect 31754 19320 31760 19332
rect 31812 19360 31818 19372
rect 32401 19363 32459 19369
rect 31812 19332 32352 19360
rect 31812 19320 31818 19332
rect 32324 19304 32352 19332
rect 32401 19329 32413 19363
rect 32447 19360 32459 19363
rect 34330 19360 34336 19372
rect 32447 19332 32628 19360
rect 34291 19332 34336 19360
rect 32447 19329 32459 19332
rect 32401 19323 32459 19329
rect 23106 19252 23112 19304
rect 23164 19292 23170 19304
rect 24302 19292 24308 19304
rect 23164 19264 24308 19292
rect 23164 19252 23170 19264
rect 24302 19252 24308 19264
rect 24360 19252 24366 19304
rect 26234 19252 26240 19304
rect 26292 19292 26298 19304
rect 27433 19295 27491 19301
rect 27433 19292 27445 19295
rect 26292 19264 27445 19292
rect 26292 19252 26298 19264
rect 27433 19261 27445 19264
rect 27479 19292 27491 19295
rect 27985 19295 28043 19301
rect 27985 19292 27997 19295
rect 27479 19264 27997 19292
rect 27479 19261 27491 19264
rect 27433 19255 27491 19261
rect 27985 19261 27997 19264
rect 28031 19261 28043 19295
rect 27985 19255 28043 19261
rect 31018 19252 31024 19304
rect 31076 19292 31082 19304
rect 32217 19295 32275 19301
rect 32217 19292 32229 19295
rect 31076 19264 32229 19292
rect 31076 19252 31082 19264
rect 32217 19261 32229 19264
rect 32263 19261 32275 19295
rect 32217 19255 32275 19261
rect 32306 19252 32312 19304
rect 32364 19292 32370 19304
rect 32493 19295 32551 19301
rect 32364 19264 32409 19292
rect 32364 19252 32370 19264
rect 32493 19261 32505 19295
rect 32539 19261 32551 19295
rect 32493 19255 32551 19261
rect 21968 19196 22324 19224
rect 23017 19227 23075 19233
rect 21968 19184 21974 19196
rect 23017 19193 23029 19227
rect 23063 19224 23075 19227
rect 28994 19224 29000 19236
rect 23063 19196 29000 19224
rect 23063 19193 23075 19196
rect 23017 19187 23075 19193
rect 28994 19184 29000 19196
rect 29052 19184 29058 19236
rect 31386 19184 31392 19236
rect 31444 19224 31450 19236
rect 32508 19224 32536 19255
rect 31444 19196 32536 19224
rect 31444 19184 31450 19196
rect 1765 19159 1823 19165
rect 1765 19125 1777 19159
rect 1811 19156 1823 19159
rect 2682 19156 2688 19168
rect 1811 19128 2688 19156
rect 1811 19125 1823 19128
rect 1765 19119 1823 19125
rect 2682 19116 2688 19128
rect 2740 19116 2746 19168
rect 4062 19156 4068 19168
rect 4023 19128 4068 19156
rect 4062 19116 4068 19128
rect 4120 19116 4126 19168
rect 12805 19159 12863 19165
rect 12805 19125 12817 19159
rect 12851 19156 12863 19159
rect 12986 19156 12992 19168
rect 12851 19128 12992 19156
rect 12851 19125 12863 19128
rect 12805 19119 12863 19125
rect 12986 19116 12992 19128
rect 13044 19116 13050 19168
rect 16114 19116 16120 19168
rect 16172 19156 16178 19168
rect 16482 19156 16488 19168
rect 16172 19128 16488 19156
rect 16172 19116 16178 19128
rect 16482 19116 16488 19128
rect 16540 19156 16546 19168
rect 18138 19156 18144 19168
rect 16540 19128 18144 19156
rect 16540 19116 16546 19128
rect 18138 19116 18144 19128
rect 18196 19116 18202 19168
rect 21177 19159 21235 19165
rect 21177 19125 21189 19159
rect 21223 19156 21235 19159
rect 23382 19156 23388 19168
rect 21223 19128 23388 19156
rect 21223 19125 21235 19128
rect 21177 19119 21235 19125
rect 23382 19116 23388 19128
rect 23440 19116 23446 19168
rect 29454 19116 29460 19168
rect 29512 19156 29518 19168
rect 31478 19156 31484 19168
rect 29512 19128 31484 19156
rect 29512 19116 29518 19128
rect 31478 19116 31484 19128
rect 31536 19116 31542 19168
rect 31754 19116 31760 19168
rect 31812 19156 31818 19168
rect 32600 19156 32628 19332
rect 34330 19320 34336 19332
rect 34388 19320 34394 19372
rect 36170 19360 36176 19372
rect 34532 19332 36176 19360
rect 34532 19233 34560 19332
rect 36170 19320 36176 19332
rect 36228 19320 36234 19372
rect 36998 19320 37004 19372
rect 37056 19360 37062 19372
rect 37182 19360 37188 19372
rect 37056 19332 37188 19360
rect 37056 19320 37062 19332
rect 37182 19320 37188 19332
rect 37240 19360 37246 19372
rect 38105 19363 38163 19369
rect 38105 19360 38117 19363
rect 37240 19332 38117 19360
rect 37240 19320 37246 19332
rect 38105 19329 38117 19332
rect 38151 19329 38163 19363
rect 38105 19323 38163 19329
rect 42702 19320 42708 19372
rect 42760 19360 42766 19372
rect 42981 19363 43039 19369
rect 42981 19360 42993 19363
rect 42760 19332 42993 19360
rect 42760 19320 42766 19332
rect 42981 19329 42993 19332
rect 43027 19329 43039 19363
rect 43809 19363 43867 19369
rect 43809 19360 43821 19363
rect 42981 19323 43039 19329
rect 43088 19332 43821 19360
rect 38010 19292 38016 19304
rect 37971 19264 38016 19292
rect 38010 19252 38016 19264
rect 38068 19252 38074 19304
rect 42794 19292 42800 19304
rect 42755 19264 42800 19292
rect 42794 19252 42800 19264
rect 42852 19292 42858 19304
rect 43088 19292 43116 19332
rect 43809 19329 43821 19332
rect 43855 19329 43867 19363
rect 43990 19360 43996 19372
rect 43951 19332 43996 19360
rect 43809 19323 43867 19329
rect 43990 19320 43996 19332
rect 44048 19320 44054 19372
rect 45557 19363 45615 19369
rect 45557 19329 45569 19363
rect 45603 19329 45615 19363
rect 45557 19323 45615 19329
rect 42852 19264 43116 19292
rect 43349 19295 43407 19301
rect 42852 19252 42858 19264
rect 43349 19261 43361 19295
rect 43395 19261 43407 19295
rect 43349 19255 43407 19261
rect 34517 19227 34575 19233
rect 34517 19193 34529 19227
rect 34563 19193 34575 19227
rect 43364 19224 43392 19255
rect 45094 19252 45100 19304
rect 45152 19292 45158 19304
rect 45572 19292 45600 19323
rect 46014 19320 46020 19372
rect 46072 19320 46078 19372
rect 46569 19363 46627 19369
rect 46569 19329 46581 19363
rect 46615 19360 46627 19363
rect 46934 19360 46940 19372
rect 46615 19332 46940 19360
rect 46615 19329 46627 19332
rect 46569 19323 46627 19329
rect 46934 19320 46940 19332
rect 46992 19360 46998 19372
rect 47581 19363 47639 19369
rect 47581 19360 47593 19363
rect 46992 19332 47593 19360
rect 46992 19320 46998 19332
rect 47581 19329 47593 19332
rect 47627 19329 47639 19363
rect 47762 19360 47768 19372
rect 47723 19332 47768 19360
rect 47581 19323 47639 19329
rect 47762 19320 47768 19332
rect 47820 19320 47826 19372
rect 47872 19360 47900 19400
rect 47949 19397 47961 19431
rect 47995 19428 48007 19431
rect 50816 19428 50844 19459
rect 50982 19456 50988 19508
rect 51040 19496 51046 19508
rect 51537 19499 51595 19505
rect 51537 19496 51549 19499
rect 51040 19468 51549 19496
rect 51040 19456 51046 19468
rect 51537 19465 51549 19468
rect 51583 19465 51595 19499
rect 51537 19459 51595 19465
rect 56226 19456 56232 19508
rect 56284 19496 56290 19508
rect 57238 19496 57244 19508
rect 56284 19468 57244 19496
rect 56284 19456 56290 19468
rect 57238 19456 57244 19468
rect 57296 19456 57302 19508
rect 51353 19431 51411 19437
rect 51353 19428 51365 19431
rect 47995 19400 49464 19428
rect 47995 19397 48007 19400
rect 47949 19391 48007 19397
rect 48774 19360 48780 19372
rect 47872 19332 48636 19360
rect 48735 19332 48780 19360
rect 45152 19264 45600 19292
rect 48608 19292 48636 19332
rect 48774 19320 48780 19332
rect 48832 19320 48838 19372
rect 48958 19360 48964 19372
rect 48884 19332 48964 19360
rect 48884 19292 48912 19332
rect 48958 19320 48964 19332
rect 49016 19360 49022 19372
rect 49436 19369 49464 19400
rect 50172 19400 50568 19428
rect 50816 19400 51365 19428
rect 50172 19372 50200 19400
rect 49421 19363 49479 19369
rect 49016 19332 49109 19360
rect 49016 19320 49022 19332
rect 49421 19329 49433 19363
rect 49467 19329 49479 19363
rect 49421 19323 49479 19329
rect 48608 19264 48912 19292
rect 49436 19292 49464 19323
rect 49510 19320 49516 19372
rect 49568 19360 49574 19372
rect 49694 19360 49700 19372
rect 49568 19332 49613 19360
rect 49655 19332 49700 19360
rect 49568 19320 49574 19332
rect 49694 19320 49700 19332
rect 49752 19320 49758 19372
rect 49789 19363 49847 19369
rect 49789 19329 49801 19363
rect 49835 19360 49847 19363
rect 50154 19360 50160 19372
rect 49835 19332 50160 19360
rect 49835 19329 49847 19332
rect 49789 19323 49847 19329
rect 50154 19320 50160 19332
rect 50212 19320 50218 19372
rect 50430 19360 50436 19372
rect 50391 19332 50436 19360
rect 50430 19320 50436 19332
rect 50488 19320 50494 19372
rect 50540 19360 50568 19400
rect 51353 19397 51365 19400
rect 51399 19397 51411 19431
rect 51353 19391 51411 19397
rect 56594 19388 56600 19440
rect 56652 19428 56658 19440
rect 56965 19431 57023 19437
rect 56965 19428 56977 19431
rect 56652 19400 56977 19428
rect 56652 19388 56658 19400
rect 56965 19397 56977 19400
rect 57011 19397 57023 19431
rect 56965 19391 57023 19397
rect 50801 19363 50859 19369
rect 50801 19360 50813 19363
rect 50540 19332 50813 19360
rect 50801 19329 50813 19332
rect 50847 19329 50859 19363
rect 50801 19323 50859 19329
rect 53466 19320 53472 19372
rect 53524 19360 53530 19372
rect 54021 19363 54079 19369
rect 54021 19360 54033 19363
rect 53524 19332 54033 19360
rect 53524 19320 53530 19332
rect 54021 19329 54033 19332
rect 54067 19360 54079 19363
rect 54662 19360 54668 19372
rect 54067 19332 54668 19360
rect 54067 19329 54079 19332
rect 54021 19323 54079 19329
rect 54662 19320 54668 19332
rect 54720 19320 54726 19372
rect 56781 19363 56839 19369
rect 56781 19329 56793 19363
rect 56827 19360 56839 19363
rect 56870 19360 56876 19372
rect 56827 19332 56876 19360
rect 56827 19329 56839 19332
rect 56781 19323 56839 19329
rect 56870 19320 56876 19332
rect 56928 19360 56934 19372
rect 57882 19360 57888 19372
rect 56928 19332 57888 19360
rect 56928 19320 56934 19332
rect 57882 19320 57888 19332
rect 57940 19320 57946 19372
rect 49602 19292 49608 19304
rect 49436 19264 49608 19292
rect 45152 19252 45158 19264
rect 49602 19252 49608 19264
rect 49660 19292 49666 19304
rect 50525 19295 50583 19301
rect 50525 19292 50537 19295
rect 49660 19264 50537 19292
rect 49660 19252 49666 19264
rect 50525 19261 50537 19264
rect 50571 19261 50583 19295
rect 50525 19255 50583 19261
rect 50614 19252 50620 19304
rect 50672 19292 50678 19304
rect 50709 19295 50767 19301
rect 50709 19292 50721 19295
rect 50672 19264 50721 19292
rect 50672 19252 50678 19264
rect 50709 19261 50721 19264
rect 50755 19261 50767 19295
rect 50709 19255 50767 19261
rect 52730 19252 52736 19304
rect 52788 19292 52794 19304
rect 53558 19292 53564 19304
rect 52788 19264 53564 19292
rect 52788 19252 52794 19264
rect 53558 19252 53564 19264
rect 53616 19252 53622 19304
rect 53926 19292 53932 19304
rect 53887 19264 53932 19292
rect 53926 19252 53932 19264
rect 53984 19252 53990 19304
rect 34517 19187 34575 19193
rect 41800 19196 43392 19224
rect 48777 19227 48835 19233
rect 41800 19168 41828 19196
rect 48777 19193 48789 19227
rect 48823 19224 48835 19227
rect 49878 19224 49884 19236
rect 48823 19196 49884 19224
rect 48823 19193 48835 19196
rect 48777 19187 48835 19193
rect 49878 19184 49884 19196
rect 49936 19184 49942 19236
rect 49973 19227 50031 19233
rect 49973 19193 49985 19227
rect 50019 19224 50031 19227
rect 50019 19196 50752 19224
rect 50019 19193 50031 19196
rect 49973 19187 50031 19193
rect 50724 19168 50752 19196
rect 31812 19128 32628 19156
rect 38381 19159 38439 19165
rect 31812 19116 31818 19128
rect 38381 19125 38393 19159
rect 38427 19156 38439 19159
rect 40310 19156 40316 19168
rect 38427 19128 40316 19156
rect 38427 19125 38439 19128
rect 38381 19119 38439 19125
rect 40310 19116 40316 19128
rect 40368 19116 40374 19168
rect 41782 19156 41788 19168
rect 41743 19128 41788 19156
rect 41782 19116 41788 19128
rect 41840 19116 41846 19168
rect 50706 19116 50712 19168
rect 50764 19156 50770 19168
rect 51537 19159 51595 19165
rect 51537 19156 51549 19159
rect 50764 19128 51549 19156
rect 50764 19116 50770 19128
rect 51537 19125 51549 19128
rect 51583 19125 51595 19159
rect 51718 19156 51724 19168
rect 51679 19128 51724 19156
rect 51537 19119 51595 19125
rect 51718 19116 51724 19128
rect 51776 19116 51782 19168
rect 54205 19159 54263 19165
rect 54205 19125 54217 19159
rect 54251 19156 54263 19159
rect 56594 19156 56600 19168
rect 54251 19128 56600 19156
rect 54251 19125 54263 19128
rect 54205 19119 54263 19125
rect 56594 19116 56600 19128
rect 56652 19116 56658 19168
rect 57146 19156 57152 19168
rect 57059 19128 57152 19156
rect 57146 19116 57152 19128
rect 57204 19156 57210 19168
rect 57698 19156 57704 19168
rect 57204 19128 57704 19156
rect 57204 19116 57210 19128
rect 57698 19116 57704 19128
rect 57756 19116 57762 19168
rect 1104 19066 58880 19088
rect 1104 19014 4214 19066
rect 4266 19014 4278 19066
rect 4330 19014 4342 19066
rect 4394 19014 4406 19066
rect 4458 19014 4470 19066
rect 4522 19014 34934 19066
rect 34986 19014 34998 19066
rect 35050 19014 35062 19066
rect 35114 19014 35126 19066
rect 35178 19014 35190 19066
rect 35242 19014 58880 19066
rect 1104 18992 58880 19014
rect 1394 18952 1400 18964
rect 1355 18924 1400 18952
rect 1394 18912 1400 18924
rect 1452 18912 1458 18964
rect 4062 18912 4068 18964
rect 4120 18952 4126 18964
rect 7469 18955 7527 18961
rect 7469 18952 7481 18955
rect 4120 18924 7481 18952
rect 4120 18912 4126 18924
rect 7469 18921 7481 18924
rect 7515 18952 7527 18955
rect 7742 18952 7748 18964
rect 7515 18924 7748 18952
rect 7515 18921 7527 18924
rect 7469 18915 7527 18921
rect 7742 18912 7748 18924
rect 7800 18912 7806 18964
rect 10229 18955 10287 18961
rect 10229 18921 10241 18955
rect 10275 18952 10287 18955
rect 11054 18952 11060 18964
rect 10275 18924 11060 18952
rect 10275 18921 10287 18924
rect 10229 18915 10287 18921
rect 11054 18912 11060 18924
rect 11112 18912 11118 18964
rect 11149 18955 11207 18961
rect 11149 18921 11161 18955
rect 11195 18952 11207 18955
rect 17862 18952 17868 18964
rect 11195 18924 17868 18952
rect 11195 18921 11207 18924
rect 11149 18915 11207 18921
rect 5721 18887 5779 18893
rect 5721 18853 5733 18887
rect 5767 18884 5779 18887
rect 10502 18884 10508 18896
rect 5767 18856 10508 18884
rect 5767 18853 5779 18856
rect 5721 18847 5779 18853
rect 10502 18844 10508 18856
rect 10560 18844 10566 18896
rect 17420 18893 17448 18924
rect 17862 18912 17868 18924
rect 17920 18912 17926 18964
rect 18046 18952 18052 18964
rect 18007 18924 18052 18952
rect 18046 18912 18052 18924
rect 18104 18912 18110 18964
rect 19613 18955 19671 18961
rect 19613 18921 19625 18955
rect 19659 18952 19671 18955
rect 19702 18952 19708 18964
rect 19659 18924 19708 18952
rect 19659 18921 19671 18924
rect 19613 18915 19671 18921
rect 19702 18912 19708 18924
rect 19760 18952 19766 18964
rect 20622 18952 20628 18964
rect 19760 18924 20628 18952
rect 19760 18912 19766 18924
rect 20622 18912 20628 18924
rect 20680 18912 20686 18964
rect 22189 18955 22247 18961
rect 22189 18921 22201 18955
rect 22235 18952 22247 18955
rect 22370 18952 22376 18964
rect 22235 18924 22376 18952
rect 22235 18921 22247 18924
rect 22189 18915 22247 18921
rect 22370 18912 22376 18924
rect 22428 18912 22434 18964
rect 23474 18912 23480 18964
rect 23532 18952 23538 18964
rect 24397 18955 24455 18961
rect 24397 18952 24409 18955
rect 23532 18924 24409 18952
rect 23532 18912 23538 18924
rect 24397 18921 24409 18924
rect 24443 18921 24455 18955
rect 24397 18915 24455 18921
rect 27154 18912 27160 18964
rect 27212 18952 27218 18964
rect 28994 18952 29000 18964
rect 27212 18924 29000 18952
rect 27212 18912 27218 18924
rect 28994 18912 29000 18924
rect 29052 18952 29058 18964
rect 30650 18952 30656 18964
rect 29052 18924 30656 18952
rect 29052 18912 29058 18924
rect 30650 18912 30656 18924
rect 30708 18912 30714 18964
rect 31018 18952 31024 18964
rect 30979 18924 31024 18952
rect 31018 18912 31024 18924
rect 31076 18912 31082 18964
rect 32858 18952 32864 18964
rect 32819 18924 32864 18952
rect 32858 18912 32864 18924
rect 32916 18912 32922 18964
rect 34149 18955 34207 18961
rect 34149 18921 34161 18955
rect 34195 18952 34207 18955
rect 34698 18952 34704 18964
rect 34195 18924 34704 18952
rect 34195 18921 34207 18924
rect 34149 18915 34207 18921
rect 34698 18912 34704 18924
rect 34756 18912 34762 18964
rect 42705 18955 42763 18961
rect 42705 18921 42717 18955
rect 42751 18952 42763 18955
rect 43990 18952 43996 18964
rect 42751 18924 43996 18952
rect 42751 18921 42763 18924
rect 42705 18915 42763 18921
rect 43990 18912 43996 18924
rect 44048 18912 44054 18964
rect 46017 18955 46075 18961
rect 46017 18921 46029 18955
rect 46063 18952 46075 18955
rect 49510 18952 49516 18964
rect 46063 18924 49516 18952
rect 46063 18921 46075 18924
rect 46017 18915 46075 18921
rect 49510 18912 49516 18924
rect 49568 18952 49574 18964
rect 50430 18952 50436 18964
rect 49568 18924 50436 18952
rect 49568 18912 49574 18924
rect 50430 18912 50436 18924
rect 50488 18912 50494 18964
rect 51718 18912 51724 18964
rect 51776 18952 51782 18964
rect 52365 18955 52423 18961
rect 52365 18952 52377 18955
rect 51776 18924 52377 18952
rect 51776 18912 51782 18924
rect 52365 18921 52377 18924
rect 52411 18952 52423 18955
rect 53190 18952 53196 18964
rect 52411 18924 53196 18952
rect 52411 18921 52423 18924
rect 52365 18915 52423 18921
rect 53190 18912 53196 18924
rect 53248 18912 53254 18964
rect 53466 18912 53472 18964
rect 53524 18952 53530 18964
rect 53745 18955 53803 18961
rect 53745 18952 53757 18955
rect 53524 18924 53757 18952
rect 53524 18912 53530 18924
rect 53745 18921 53757 18924
rect 53791 18921 53803 18955
rect 53745 18915 53803 18921
rect 17405 18887 17463 18893
rect 10796 18856 16344 18884
rect 7466 18816 7472 18828
rect 7392 18788 7472 18816
rect 1578 18708 1584 18760
rect 1636 18748 1642 18760
rect 2317 18751 2375 18757
rect 2317 18748 2329 18751
rect 1636 18720 2329 18748
rect 1636 18708 1642 18720
rect 2317 18717 2329 18720
rect 2363 18717 2375 18751
rect 2317 18711 2375 18717
rect 4062 18708 4068 18760
rect 4120 18748 4126 18760
rect 4249 18751 4307 18757
rect 4249 18748 4261 18751
rect 4120 18720 4261 18748
rect 4120 18708 4126 18720
rect 4249 18717 4261 18720
rect 4295 18717 4307 18751
rect 4890 18748 4896 18760
rect 4851 18720 4896 18748
rect 4249 18711 4307 18717
rect 4890 18708 4896 18720
rect 4948 18708 4954 18760
rect 7190 18748 7196 18760
rect 7151 18720 7196 18748
rect 7190 18708 7196 18720
rect 7248 18708 7254 18760
rect 7392 18757 7420 18788
rect 7466 18776 7472 18788
rect 7524 18776 7530 18828
rect 7653 18819 7711 18825
rect 7653 18785 7665 18819
rect 7699 18816 7711 18819
rect 8018 18816 8024 18828
rect 7699 18788 8024 18816
rect 7699 18785 7711 18788
rect 7653 18779 7711 18785
rect 8018 18776 8024 18788
rect 8076 18776 8082 18828
rect 7377 18751 7435 18757
rect 7377 18717 7389 18751
rect 7423 18717 7435 18751
rect 7558 18748 7564 18760
rect 7519 18720 7564 18748
rect 7377 18711 7435 18717
rect 7558 18708 7564 18720
rect 7616 18708 7622 18760
rect 2501 18683 2559 18689
rect 2501 18649 2513 18683
rect 2547 18680 2559 18683
rect 4982 18680 4988 18692
rect 2547 18652 4988 18680
rect 2547 18649 2559 18652
rect 2501 18643 2559 18649
rect 4982 18640 4988 18652
rect 5040 18640 5046 18692
rect 6270 18640 6276 18692
rect 6328 18680 6334 18692
rect 10796 18680 10824 18856
rect 10965 18819 11023 18825
rect 10965 18785 10977 18819
rect 11011 18816 11023 18819
rect 11701 18819 11759 18825
rect 11701 18816 11713 18819
rect 11011 18788 11713 18816
rect 11011 18785 11023 18788
rect 10965 18779 11023 18785
rect 11701 18785 11713 18788
rect 11747 18816 11759 18819
rect 13538 18816 13544 18828
rect 11747 18788 12434 18816
rect 13499 18788 13544 18816
rect 11747 18785 11759 18788
rect 11701 18779 11759 18785
rect 10873 18751 10931 18757
rect 10873 18717 10885 18751
rect 10919 18748 10931 18751
rect 11054 18748 11060 18760
rect 10919 18720 11060 18748
rect 10919 18717 10931 18720
rect 10873 18711 10931 18717
rect 11054 18708 11060 18720
rect 11112 18708 11118 18760
rect 6328 18652 10824 18680
rect 6328 18640 6334 18652
rect 7929 18615 7987 18621
rect 7929 18581 7941 18615
rect 7975 18612 7987 18615
rect 8662 18612 8668 18624
rect 7975 18584 8668 18612
rect 7975 18581 7987 18584
rect 7929 18575 7987 18581
rect 8662 18572 8668 18584
rect 8720 18572 8726 18624
rect 12406 18612 12434 18788
rect 13538 18776 13544 18788
rect 13596 18776 13602 18828
rect 15194 18816 15200 18828
rect 15155 18788 15200 18816
rect 15194 18776 15200 18788
rect 15252 18776 15258 18828
rect 14366 18748 14372 18760
rect 14327 18720 14372 18748
rect 14366 18708 14372 18720
rect 14424 18708 14430 18760
rect 14918 18748 14924 18760
rect 14879 18720 14924 18748
rect 14918 18708 14924 18720
rect 14976 18708 14982 18760
rect 15286 18748 15292 18760
rect 15247 18720 15292 18748
rect 15286 18708 15292 18720
rect 15344 18708 15350 18760
rect 15841 18751 15899 18757
rect 15841 18717 15853 18751
rect 15887 18717 15899 18751
rect 16206 18748 16212 18760
rect 16119 18720 16212 18748
rect 15841 18711 15899 18717
rect 14734 18640 14740 18692
rect 14792 18680 14798 18692
rect 15856 18680 15884 18711
rect 16206 18708 16212 18720
rect 16264 18708 16270 18760
rect 16316 18748 16344 18856
rect 17405 18853 17417 18887
rect 17451 18853 17463 18887
rect 17405 18847 17463 18853
rect 20165 18887 20223 18893
rect 20165 18853 20177 18887
rect 20211 18884 20223 18887
rect 20714 18884 20720 18896
rect 20211 18856 20720 18884
rect 20211 18853 20223 18856
rect 20165 18847 20223 18853
rect 20714 18844 20720 18856
rect 20772 18884 20778 18896
rect 21266 18884 21272 18896
rect 20772 18856 21272 18884
rect 20772 18844 20778 18856
rect 21266 18844 21272 18856
rect 21324 18844 21330 18896
rect 27614 18884 27620 18896
rect 21376 18856 26556 18884
rect 27575 18856 27620 18884
rect 21376 18816 21404 18856
rect 17604 18788 21404 18816
rect 17604 18748 17632 18788
rect 21450 18776 21456 18828
rect 21508 18816 21514 18828
rect 21508 18788 21864 18816
rect 21508 18776 21514 18788
rect 16316 18720 17632 18748
rect 17862 18708 17868 18760
rect 17920 18748 17926 18760
rect 18049 18751 18107 18757
rect 18049 18748 18061 18751
rect 17920 18720 18061 18748
rect 17920 18708 17926 18720
rect 18049 18717 18061 18720
rect 18095 18717 18107 18751
rect 18049 18711 18107 18717
rect 18233 18751 18291 18757
rect 18233 18717 18245 18751
rect 18279 18748 18291 18751
rect 19242 18748 19248 18760
rect 18279 18720 19248 18748
rect 18279 18717 18291 18720
rect 18233 18711 18291 18717
rect 16114 18680 16120 18692
rect 14792 18652 16120 18680
rect 14792 18640 14798 18652
rect 16114 18640 16120 18652
rect 16172 18640 16178 18692
rect 16224 18680 16252 18708
rect 16942 18680 16948 18692
rect 16224 18652 16948 18680
rect 16942 18640 16948 18652
rect 17000 18640 17006 18692
rect 17129 18683 17187 18689
rect 17129 18649 17141 18683
rect 17175 18680 17187 18683
rect 17770 18680 17776 18692
rect 17175 18652 17776 18680
rect 17175 18649 17187 18652
rect 17129 18643 17187 18649
rect 17770 18640 17776 18652
rect 17828 18680 17834 18692
rect 18248 18680 18276 18711
rect 19242 18708 19248 18720
rect 19300 18708 19306 18760
rect 19429 18751 19487 18757
rect 19429 18717 19441 18751
rect 19475 18717 19487 18751
rect 19429 18711 19487 18717
rect 17828 18652 18276 18680
rect 17828 18640 17834 18652
rect 18874 18640 18880 18692
rect 18932 18680 18938 18692
rect 19444 18680 19472 18711
rect 20806 18708 20812 18760
rect 20864 18748 20870 18760
rect 21637 18751 21695 18757
rect 21637 18748 21649 18751
rect 20864 18720 21649 18748
rect 20864 18708 20870 18720
rect 21637 18717 21649 18720
rect 21683 18748 21695 18751
rect 21726 18748 21732 18760
rect 21683 18720 21732 18748
rect 21683 18717 21695 18720
rect 21637 18711 21695 18717
rect 21726 18708 21732 18720
rect 21784 18708 21790 18760
rect 21836 18748 21864 18788
rect 22094 18776 22100 18828
rect 22152 18816 22158 18828
rect 22152 18788 24624 18816
rect 22152 18776 22158 18788
rect 21913 18751 21971 18757
rect 21913 18748 21925 18751
rect 21836 18720 21925 18748
rect 21913 18717 21925 18720
rect 21959 18717 21971 18751
rect 21913 18711 21971 18717
rect 22005 18751 22063 18757
rect 22005 18717 22017 18751
rect 22051 18748 22063 18751
rect 23198 18748 23204 18760
rect 22051 18720 23204 18748
rect 22051 18717 22063 18720
rect 22005 18711 22063 18717
rect 23198 18708 23204 18720
rect 23256 18708 23262 18760
rect 24596 18757 24624 18788
rect 24397 18751 24455 18757
rect 24397 18717 24409 18751
rect 24443 18717 24455 18751
rect 24397 18711 24455 18717
rect 24581 18751 24639 18757
rect 24581 18717 24593 18751
rect 24627 18748 24639 18751
rect 25041 18751 25099 18757
rect 25041 18748 25053 18751
rect 24627 18720 25053 18748
rect 24627 18717 24639 18720
rect 24581 18711 24639 18717
rect 25041 18717 25053 18720
rect 25087 18717 25099 18751
rect 25682 18748 25688 18760
rect 25643 18720 25688 18748
rect 25041 18711 25099 18717
rect 18932 18652 19472 18680
rect 18932 18640 18938 18652
rect 21358 18640 21364 18692
rect 21416 18680 21422 18692
rect 21818 18680 21824 18692
rect 21416 18652 21824 18680
rect 21416 18640 21422 18652
rect 21818 18640 21824 18652
rect 21876 18640 21882 18692
rect 24210 18680 24216 18692
rect 22066 18652 24216 18680
rect 12802 18612 12808 18624
rect 12406 18584 12808 18612
rect 12802 18572 12808 18584
rect 12860 18572 12866 18624
rect 17589 18615 17647 18621
rect 17589 18581 17601 18615
rect 17635 18612 17647 18615
rect 17954 18612 17960 18624
rect 17635 18584 17960 18612
rect 17635 18581 17647 18584
rect 17589 18575 17647 18581
rect 17954 18572 17960 18584
rect 18012 18572 18018 18624
rect 18138 18572 18144 18624
rect 18196 18612 18202 18624
rect 22066 18612 22094 18652
rect 24210 18640 24216 18652
rect 24268 18640 24274 18692
rect 18196 18584 22094 18612
rect 23845 18615 23903 18621
rect 18196 18572 18202 18584
rect 23845 18581 23857 18615
rect 23891 18612 23903 18615
rect 24412 18612 24440 18711
rect 24486 18612 24492 18624
rect 23891 18584 24492 18612
rect 23891 18581 23903 18584
rect 23845 18575 23903 18581
rect 24486 18572 24492 18584
rect 24544 18572 24550 18624
rect 25056 18612 25084 18711
rect 25682 18708 25688 18720
rect 25740 18708 25746 18760
rect 26053 18751 26111 18757
rect 26053 18717 26065 18751
rect 26099 18748 26111 18751
rect 26418 18748 26424 18760
rect 26099 18720 26424 18748
rect 26099 18717 26111 18720
rect 26053 18711 26111 18717
rect 26418 18708 26424 18720
rect 26476 18708 26482 18760
rect 26528 18748 26556 18856
rect 27614 18844 27620 18856
rect 27672 18844 27678 18896
rect 27706 18844 27712 18896
rect 27764 18884 27770 18896
rect 31202 18884 31208 18896
rect 27764 18856 31208 18884
rect 27764 18844 27770 18856
rect 31202 18844 31208 18856
rect 31260 18844 31266 18896
rect 31478 18844 31484 18896
rect 31536 18884 31542 18896
rect 34514 18884 34520 18896
rect 31536 18856 34520 18884
rect 31536 18844 31542 18856
rect 34514 18844 34520 18856
rect 34572 18844 34578 18896
rect 35986 18844 35992 18896
rect 36044 18884 36050 18896
rect 36265 18887 36323 18893
rect 36265 18884 36277 18887
rect 36044 18856 36277 18884
rect 36044 18844 36050 18856
rect 36265 18853 36277 18856
rect 36311 18853 36323 18887
rect 36265 18847 36323 18853
rect 41785 18887 41843 18893
rect 41785 18853 41797 18887
rect 41831 18884 41843 18887
rect 42794 18884 42800 18896
rect 41831 18856 42800 18884
rect 41831 18853 41843 18856
rect 41785 18847 41843 18853
rect 42794 18844 42800 18856
rect 42852 18844 42858 18896
rect 50448 18884 50476 18912
rect 50448 18856 50568 18884
rect 27798 18776 27804 18828
rect 27856 18816 27862 18828
rect 40310 18816 40316 18828
rect 27856 18788 38516 18816
rect 40271 18788 40316 18816
rect 27856 18776 27862 18788
rect 27706 18748 27712 18760
rect 26528 18720 27712 18748
rect 27706 18708 27712 18720
rect 27764 18708 27770 18760
rect 28077 18751 28135 18757
rect 28077 18717 28089 18751
rect 28123 18748 28135 18751
rect 29178 18748 29184 18760
rect 28123 18720 29184 18748
rect 28123 18717 28135 18720
rect 28077 18711 28135 18717
rect 29178 18708 29184 18720
rect 29236 18708 29242 18760
rect 29730 18748 29736 18760
rect 29643 18720 29736 18748
rect 29730 18708 29736 18720
rect 29788 18708 29794 18760
rect 29914 18748 29920 18760
rect 29875 18720 29920 18748
rect 29914 18708 29920 18720
rect 29972 18708 29978 18760
rect 30098 18748 30104 18760
rect 30059 18720 30104 18748
rect 30098 18708 30104 18720
rect 30156 18708 30162 18760
rect 30190 18708 30196 18760
rect 30248 18748 30254 18760
rect 31021 18751 31079 18757
rect 31021 18748 31033 18751
rect 30248 18720 31033 18748
rect 30248 18708 30254 18720
rect 31021 18717 31033 18720
rect 31067 18717 31079 18751
rect 31021 18711 31079 18717
rect 31205 18751 31263 18757
rect 31205 18717 31217 18751
rect 31251 18748 31263 18751
rect 31251 18720 31754 18748
rect 31251 18717 31263 18720
rect 31205 18711 31263 18717
rect 26697 18683 26755 18689
rect 26697 18649 26709 18683
rect 26743 18680 26755 18683
rect 27522 18680 27528 18692
rect 26743 18652 27528 18680
rect 26743 18649 26755 18652
rect 26697 18643 26755 18649
rect 27522 18640 27528 18652
rect 27580 18640 27586 18692
rect 27614 18640 27620 18692
rect 27672 18680 27678 18692
rect 28261 18683 28319 18689
rect 28261 18680 28273 18683
rect 27672 18652 28273 18680
rect 27672 18640 27678 18652
rect 28261 18649 28273 18652
rect 28307 18649 28319 18683
rect 29638 18680 29644 18692
rect 28261 18643 28319 18649
rect 29288 18652 29644 18680
rect 29288 18612 29316 18652
rect 29638 18640 29644 18652
rect 29696 18640 29702 18692
rect 25056 18584 29316 18612
rect 29362 18572 29368 18624
rect 29420 18612 29426 18624
rect 29549 18615 29607 18621
rect 29549 18612 29561 18615
rect 29420 18584 29561 18612
rect 29420 18572 29426 18584
rect 29549 18581 29561 18584
rect 29595 18581 29607 18615
rect 29748 18612 29776 18708
rect 29825 18683 29883 18689
rect 29825 18649 29837 18683
rect 29871 18680 29883 18683
rect 31386 18680 31392 18692
rect 29871 18652 31392 18680
rect 29871 18649 29883 18652
rect 29825 18643 29883 18649
rect 31386 18640 31392 18652
rect 31444 18640 31450 18692
rect 31726 18624 31754 18720
rect 31846 18708 31852 18760
rect 31904 18748 31910 18760
rect 33594 18748 33600 18760
rect 31904 18720 31949 18748
rect 33555 18720 33600 18748
rect 31904 18708 31910 18720
rect 33594 18708 33600 18720
rect 33652 18708 33658 18760
rect 33689 18751 33747 18757
rect 33689 18717 33701 18751
rect 33735 18717 33747 18751
rect 33689 18711 33747 18717
rect 33873 18751 33931 18757
rect 33873 18717 33885 18751
rect 33919 18717 33931 18751
rect 33873 18711 33931 18717
rect 32306 18640 32312 18692
rect 32364 18680 32370 18692
rect 32677 18683 32735 18689
rect 32677 18680 32689 18683
rect 32364 18652 32689 18680
rect 32364 18640 32370 18652
rect 32677 18649 32689 18652
rect 32723 18649 32735 18683
rect 33704 18680 33732 18711
rect 32677 18643 32735 18649
rect 33060 18652 33732 18680
rect 33888 18680 33916 18711
rect 33962 18708 33968 18760
rect 34020 18748 34026 18760
rect 35710 18748 35716 18760
rect 34020 18720 34065 18748
rect 34256 18720 35716 18748
rect 34020 18708 34026 18720
rect 34256 18680 34284 18720
rect 35710 18708 35716 18720
rect 35768 18708 35774 18760
rect 35989 18751 36047 18757
rect 35989 18717 36001 18751
rect 36035 18748 36047 18751
rect 36354 18748 36360 18760
rect 36035 18720 36360 18748
rect 36035 18717 36047 18720
rect 35989 18711 36047 18717
rect 36354 18708 36360 18720
rect 36412 18708 36418 18760
rect 38488 18748 38516 18788
rect 40310 18776 40316 18788
rect 40368 18776 40374 18828
rect 40773 18819 40831 18825
rect 40773 18785 40785 18819
rect 40819 18816 40831 18819
rect 40819 18788 41920 18816
rect 40819 18785 40831 18788
rect 40773 18779 40831 18785
rect 40405 18751 40463 18757
rect 40405 18748 40417 18751
rect 38488 18720 40417 18748
rect 40405 18717 40417 18720
rect 40451 18748 40463 18751
rect 40678 18748 40684 18760
rect 40451 18720 40684 18748
rect 40451 18717 40463 18720
rect 40405 18711 40463 18717
rect 40678 18708 40684 18720
rect 40736 18708 40742 18760
rect 41690 18748 41696 18760
rect 41651 18720 41696 18748
rect 41690 18708 41696 18720
rect 41748 18708 41754 18760
rect 41892 18757 41920 18788
rect 49602 18776 49608 18828
rect 49660 18816 49666 18828
rect 49660 18788 50476 18816
rect 49660 18776 49666 18788
rect 41877 18751 41935 18757
rect 41877 18717 41889 18751
rect 41923 18748 41935 18751
rect 42521 18751 42579 18757
rect 42521 18748 42533 18751
rect 41923 18720 42533 18748
rect 41923 18717 41935 18720
rect 41877 18711 41935 18717
rect 42521 18717 42533 18720
rect 42567 18717 42579 18751
rect 42521 18711 42579 18717
rect 45094 18708 45100 18760
rect 45152 18748 45158 18760
rect 45833 18751 45891 18757
rect 45833 18748 45845 18751
rect 45152 18720 45845 18748
rect 45152 18708 45158 18720
rect 45833 18717 45845 18720
rect 45879 18717 45891 18751
rect 46014 18748 46020 18760
rect 45975 18720 46020 18748
rect 45833 18711 45891 18717
rect 46014 18708 46020 18720
rect 46072 18708 46078 18760
rect 50154 18748 50160 18760
rect 50115 18720 50160 18748
rect 50154 18708 50160 18720
rect 50212 18708 50218 18760
rect 50448 18757 50476 18788
rect 50540 18757 50568 18856
rect 52546 18844 52552 18896
rect 52604 18884 52610 18896
rect 52604 18856 53512 18884
rect 52604 18844 52610 18856
rect 50801 18819 50859 18825
rect 50801 18785 50813 18819
rect 50847 18785 50859 18819
rect 50801 18779 50859 18785
rect 52288 18788 53328 18816
rect 50341 18751 50399 18757
rect 50341 18717 50353 18751
rect 50387 18717 50399 18751
rect 50341 18711 50399 18717
rect 50433 18751 50491 18757
rect 50433 18717 50445 18751
rect 50479 18717 50491 18751
rect 50433 18711 50491 18717
rect 50525 18751 50583 18757
rect 50525 18717 50537 18751
rect 50571 18717 50583 18751
rect 50816 18748 50844 18779
rect 52288 18757 52316 18788
rect 52273 18751 52331 18757
rect 52273 18748 52285 18751
rect 50816 18720 52285 18748
rect 50525 18711 50583 18717
rect 52273 18717 52285 18720
rect 52319 18717 52331 18751
rect 52546 18748 52552 18760
rect 52507 18720 52552 18748
rect 52273 18711 52331 18717
rect 33888 18652 34284 18680
rect 31294 18612 31300 18624
rect 29748 18584 31300 18612
rect 29549 18575 29607 18581
rect 31294 18572 31300 18584
rect 31352 18572 31358 18624
rect 31726 18584 31760 18624
rect 31754 18572 31760 18584
rect 31812 18612 31818 18624
rect 31812 18584 31857 18612
rect 31812 18572 31818 18584
rect 32398 18572 32404 18624
rect 32456 18612 32462 18624
rect 33060 18621 33088 18652
rect 32877 18615 32935 18621
rect 32877 18612 32889 18615
rect 32456 18584 32889 18612
rect 32456 18572 32462 18584
rect 32877 18581 32889 18584
rect 32923 18581 32935 18615
rect 32877 18575 32935 18581
rect 33045 18615 33103 18621
rect 33045 18581 33057 18615
rect 33091 18581 33103 18615
rect 33045 18575 33103 18581
rect 33134 18572 33140 18624
rect 33192 18612 33198 18624
rect 33888 18612 33916 18652
rect 34330 18640 34336 18692
rect 34388 18680 34394 18692
rect 36262 18680 36268 18692
rect 34388 18652 36268 18680
rect 34388 18640 34394 18652
rect 36262 18640 36268 18652
rect 36320 18640 36326 18692
rect 41708 18680 41736 18708
rect 42337 18683 42395 18689
rect 42337 18680 42349 18683
rect 41708 18652 42349 18680
rect 42337 18649 42349 18652
rect 42383 18649 42395 18683
rect 42337 18643 42395 18649
rect 49694 18640 49700 18692
rect 49752 18680 49758 18692
rect 50356 18680 50384 18711
rect 52546 18708 52552 18720
rect 52604 18708 52610 18760
rect 52641 18751 52699 18757
rect 52641 18717 52653 18751
rect 52687 18717 52699 18751
rect 53190 18748 53196 18760
rect 53151 18720 53196 18748
rect 52641 18711 52699 18717
rect 50614 18680 50620 18692
rect 49752 18652 50620 18680
rect 49752 18640 49758 18652
rect 50614 18640 50620 18652
rect 50672 18640 50678 18692
rect 52656 18680 52684 18711
rect 53190 18708 53196 18720
rect 53248 18708 53254 18760
rect 53300 18757 53328 18788
rect 53484 18760 53512 18856
rect 56778 18816 56784 18828
rect 56739 18788 56784 18816
rect 56778 18776 56784 18788
rect 56836 18776 56842 18828
rect 57330 18816 57336 18828
rect 57291 18788 57336 18816
rect 57330 18776 57336 18788
rect 57388 18776 57394 18828
rect 53285 18751 53343 18757
rect 53285 18717 53297 18751
rect 53331 18717 53343 18751
rect 53466 18748 53472 18760
rect 53427 18720 53472 18748
rect 53285 18711 53343 18717
rect 53466 18708 53472 18720
rect 53524 18708 53530 18760
rect 53561 18751 53619 18757
rect 53561 18717 53573 18751
rect 53607 18717 53619 18751
rect 56594 18748 56600 18760
rect 56555 18720 56600 18748
rect 53561 18711 53619 18717
rect 53374 18680 53380 18692
rect 52656 18652 53380 18680
rect 53374 18640 53380 18652
rect 53432 18680 53438 18692
rect 53576 18680 53604 18711
rect 56594 18708 56600 18720
rect 56652 18708 56658 18760
rect 57882 18748 57888 18760
rect 57843 18720 57888 18748
rect 57882 18708 57888 18720
rect 57940 18708 57946 18760
rect 58069 18751 58127 18757
rect 58069 18717 58081 18751
rect 58115 18717 58127 18751
rect 58069 18711 58127 18717
rect 53432 18652 53604 18680
rect 53432 18640 53438 18652
rect 56686 18640 56692 18692
rect 56744 18680 56750 18692
rect 58084 18680 58112 18711
rect 56744 18652 58112 18680
rect 56744 18640 56750 18652
rect 33192 18584 33916 18612
rect 33192 18572 33198 18584
rect 34514 18572 34520 18624
rect 34572 18612 34578 18624
rect 35894 18612 35900 18624
rect 34572 18584 35900 18612
rect 34572 18572 34578 18584
rect 35894 18572 35900 18584
rect 35952 18612 35958 18624
rect 36081 18615 36139 18621
rect 36081 18612 36093 18615
rect 35952 18584 36093 18612
rect 35952 18572 35958 18584
rect 36081 18581 36093 18584
rect 36127 18581 36139 18615
rect 52730 18612 52736 18624
rect 52691 18584 52736 18612
rect 36081 18575 36139 18581
rect 52730 18572 52736 18584
rect 52788 18572 52794 18624
rect 57790 18572 57796 18624
rect 57848 18612 57854 18624
rect 57977 18615 58035 18621
rect 57977 18612 57989 18615
rect 57848 18584 57989 18612
rect 57848 18572 57854 18584
rect 57977 18581 57989 18584
rect 58023 18581 58035 18615
rect 57977 18575 58035 18581
rect 1104 18522 58880 18544
rect 1104 18470 19574 18522
rect 19626 18470 19638 18522
rect 19690 18470 19702 18522
rect 19754 18470 19766 18522
rect 19818 18470 19830 18522
rect 19882 18470 50294 18522
rect 50346 18470 50358 18522
rect 50410 18470 50422 18522
rect 50474 18470 50486 18522
rect 50538 18470 50550 18522
rect 50602 18470 58880 18522
rect 1104 18448 58880 18470
rect 2406 18368 2412 18420
rect 2464 18408 2470 18420
rect 2777 18411 2835 18417
rect 2777 18408 2789 18411
rect 2464 18380 2789 18408
rect 2464 18368 2470 18380
rect 2777 18377 2789 18380
rect 2823 18377 2835 18411
rect 2777 18371 2835 18377
rect 6917 18411 6975 18417
rect 6917 18377 6929 18411
rect 6963 18408 6975 18411
rect 7558 18408 7564 18420
rect 6963 18380 7564 18408
rect 6963 18377 6975 18380
rect 6917 18371 6975 18377
rect 7558 18368 7564 18380
rect 7616 18368 7622 18420
rect 15194 18408 15200 18420
rect 14476 18380 15200 18408
rect 1578 18300 1584 18352
rect 1636 18340 1642 18352
rect 1857 18343 1915 18349
rect 1857 18340 1869 18343
rect 1636 18312 1869 18340
rect 1636 18300 1642 18312
rect 1857 18309 1869 18312
rect 1903 18309 1915 18343
rect 1857 18303 1915 18309
rect 2038 18272 2044 18284
rect 1999 18244 2044 18272
rect 2038 18232 2044 18244
rect 2096 18232 2102 18284
rect 2774 18232 2780 18284
rect 2832 18272 2838 18284
rect 3050 18272 3056 18284
rect 2832 18244 2877 18272
rect 3011 18244 3056 18272
rect 2832 18232 2838 18244
rect 3050 18232 3056 18244
rect 3108 18232 3114 18284
rect 7009 18275 7067 18281
rect 7009 18241 7021 18275
rect 7055 18272 7067 18275
rect 7190 18272 7196 18284
rect 7055 18244 7196 18272
rect 7055 18241 7067 18244
rect 7009 18235 7067 18241
rect 7190 18232 7196 18244
rect 7248 18232 7254 18284
rect 7650 18272 7656 18284
rect 7611 18244 7656 18272
rect 7650 18232 7656 18244
rect 7708 18232 7714 18284
rect 7834 18272 7840 18284
rect 7795 18244 7840 18272
rect 7834 18232 7840 18244
rect 7892 18232 7898 18284
rect 8018 18232 8024 18284
rect 8076 18272 8082 18284
rect 8297 18275 8355 18281
rect 8297 18272 8309 18275
rect 8076 18244 8309 18272
rect 8076 18232 8082 18244
rect 8297 18241 8309 18244
rect 8343 18241 8355 18275
rect 8297 18235 8355 18241
rect 10686 18232 10692 18284
rect 10744 18272 10750 18284
rect 10965 18275 11023 18281
rect 10965 18272 10977 18275
rect 10744 18244 10977 18272
rect 10744 18232 10750 18244
rect 10965 18241 10977 18244
rect 11011 18272 11023 18275
rect 11609 18275 11667 18281
rect 11609 18272 11621 18275
rect 11011 18244 11621 18272
rect 11011 18241 11023 18244
rect 10965 18235 11023 18241
rect 11609 18241 11621 18244
rect 11655 18241 11667 18275
rect 12802 18272 12808 18284
rect 12282 18244 12808 18272
rect 11609 18235 11667 18241
rect 12802 18232 12808 18244
rect 12860 18232 12866 18284
rect 14476 18281 14504 18380
rect 15194 18368 15200 18380
rect 15252 18368 15258 18420
rect 15286 18368 15292 18420
rect 15344 18408 15350 18420
rect 15657 18411 15715 18417
rect 15657 18408 15669 18411
rect 15344 18380 15669 18408
rect 15344 18368 15350 18380
rect 15657 18377 15669 18380
rect 15703 18408 15715 18411
rect 15930 18408 15936 18420
rect 15703 18380 15936 18408
rect 15703 18377 15715 18380
rect 15657 18371 15715 18377
rect 15930 18368 15936 18380
rect 15988 18368 15994 18420
rect 16114 18368 16120 18420
rect 16172 18408 16178 18420
rect 18230 18408 18236 18420
rect 16172 18380 18236 18408
rect 16172 18368 16178 18380
rect 18230 18368 18236 18380
rect 18288 18368 18294 18420
rect 18414 18368 18420 18420
rect 18472 18408 18478 18420
rect 22002 18408 22008 18420
rect 18472 18380 22008 18408
rect 18472 18368 18478 18380
rect 22002 18368 22008 18380
rect 22060 18368 22066 18420
rect 22094 18368 22100 18420
rect 22152 18408 22158 18420
rect 23106 18408 23112 18420
rect 22152 18380 23112 18408
rect 22152 18368 22158 18380
rect 23106 18368 23112 18380
rect 23164 18408 23170 18420
rect 23164 18380 24256 18408
rect 23164 18368 23170 18380
rect 14642 18340 14648 18352
rect 14603 18312 14648 18340
rect 14642 18300 14648 18312
rect 14700 18340 14706 18352
rect 15102 18340 15108 18352
rect 14700 18312 15108 18340
rect 14700 18300 14706 18312
rect 15102 18300 15108 18312
rect 15160 18300 15166 18352
rect 18046 18300 18052 18352
rect 18104 18340 18110 18352
rect 18104 18312 19288 18340
rect 18104 18300 18110 18312
rect 14461 18275 14519 18281
rect 14461 18241 14473 18275
rect 14507 18241 14519 18275
rect 14734 18272 14740 18284
rect 14695 18244 14740 18272
rect 14461 18235 14519 18241
rect 14734 18232 14740 18244
rect 14792 18232 14798 18284
rect 14826 18232 14832 18284
rect 14884 18272 14890 18284
rect 15473 18275 15531 18281
rect 15473 18272 15485 18275
rect 14884 18244 15485 18272
rect 14884 18232 14890 18244
rect 15473 18241 15485 18244
rect 15519 18241 15531 18275
rect 15473 18235 15531 18241
rect 17773 18275 17831 18281
rect 17773 18241 17785 18275
rect 17819 18272 17831 18275
rect 17954 18272 17960 18284
rect 17819 18244 17960 18272
rect 17819 18241 17831 18244
rect 17773 18235 17831 18241
rect 17954 18232 17960 18244
rect 18012 18272 18018 18284
rect 18322 18272 18328 18284
rect 18012 18244 18328 18272
rect 18012 18232 18018 18244
rect 18322 18232 18328 18244
rect 18380 18232 18386 18284
rect 19260 18281 19288 18312
rect 20162 18300 20168 18352
rect 20220 18340 20226 18352
rect 22925 18343 22983 18349
rect 22925 18340 22937 18343
rect 20220 18312 22937 18340
rect 20220 18300 20226 18312
rect 22925 18309 22937 18312
rect 22971 18340 22983 18343
rect 24118 18340 24124 18352
rect 22971 18312 24124 18340
rect 22971 18309 22983 18312
rect 22925 18303 22983 18309
rect 24118 18300 24124 18312
rect 24176 18300 24182 18352
rect 24228 18340 24256 18380
rect 26234 18368 26240 18420
rect 26292 18408 26298 18420
rect 26329 18411 26387 18417
rect 26329 18408 26341 18411
rect 26292 18380 26341 18408
rect 26292 18368 26298 18380
rect 26329 18377 26341 18380
rect 26375 18377 26387 18411
rect 29178 18408 29184 18420
rect 29139 18380 29184 18408
rect 26329 18371 26387 18377
rect 29178 18368 29184 18380
rect 29236 18368 29242 18420
rect 30650 18368 30656 18420
rect 30708 18408 30714 18420
rect 32125 18411 32183 18417
rect 32125 18408 32137 18411
rect 30708 18380 32137 18408
rect 30708 18368 30714 18380
rect 32125 18377 32137 18380
rect 32171 18377 32183 18411
rect 32125 18371 32183 18377
rect 32858 18368 32864 18420
rect 32916 18408 32922 18420
rect 34330 18408 34336 18420
rect 32916 18380 34336 18408
rect 32916 18368 32922 18380
rect 34330 18368 34336 18380
rect 34388 18368 34394 18420
rect 34514 18408 34520 18420
rect 34475 18380 34520 18408
rect 34514 18368 34520 18380
rect 34572 18368 34578 18420
rect 35710 18368 35716 18420
rect 35768 18408 35774 18420
rect 37366 18408 37372 18420
rect 35768 18380 37372 18408
rect 35768 18368 35774 18380
rect 37366 18368 37372 18380
rect 37424 18368 37430 18420
rect 40681 18411 40739 18417
rect 40681 18377 40693 18411
rect 40727 18408 40739 18411
rect 42702 18408 42708 18420
rect 40727 18380 42708 18408
rect 40727 18377 40739 18380
rect 40681 18371 40739 18377
rect 42702 18368 42708 18380
rect 42760 18368 42766 18420
rect 49329 18411 49387 18417
rect 49329 18377 49341 18411
rect 49375 18408 49387 18411
rect 50154 18408 50160 18420
rect 49375 18380 50160 18408
rect 49375 18377 49387 18380
rect 49329 18371 49387 18377
rect 50154 18368 50160 18380
rect 50212 18368 50218 18420
rect 53374 18408 53380 18420
rect 53335 18380 53380 18408
rect 53374 18368 53380 18380
rect 53432 18368 53438 18420
rect 56686 18408 56692 18420
rect 56647 18380 56692 18408
rect 56686 18368 56692 18380
rect 56744 18368 56750 18420
rect 57974 18408 57980 18420
rect 57935 18380 57980 18408
rect 57974 18368 57980 18380
rect 58032 18368 58038 18420
rect 24581 18343 24639 18349
rect 24581 18340 24593 18343
rect 24228 18312 24593 18340
rect 24581 18309 24593 18312
rect 24627 18309 24639 18343
rect 25038 18340 25044 18352
rect 24581 18303 24639 18309
rect 24871 18312 25044 18340
rect 19245 18275 19303 18281
rect 19245 18241 19257 18275
rect 19291 18241 19303 18275
rect 19886 18272 19892 18284
rect 19245 18235 19303 18241
rect 19628 18244 19892 18272
rect 8573 18207 8631 18213
rect 8573 18173 8585 18207
rect 8619 18204 8631 18207
rect 9950 18204 9956 18216
rect 8619 18176 9956 18204
rect 8619 18173 8631 18176
rect 8573 18167 8631 18173
rect 9950 18164 9956 18176
rect 10008 18164 10014 18216
rect 12621 18207 12679 18213
rect 12621 18173 12633 18207
rect 12667 18204 12679 18207
rect 16022 18204 16028 18216
rect 12667 18176 16028 18204
rect 12667 18173 12679 18176
rect 12621 18167 12679 18173
rect 16022 18164 16028 18176
rect 16080 18204 16086 18216
rect 17589 18207 17647 18213
rect 17589 18204 17601 18207
rect 16080 18176 17601 18204
rect 16080 18164 16086 18176
rect 17589 18173 17601 18176
rect 17635 18204 17647 18207
rect 18874 18204 18880 18216
rect 17635 18176 18880 18204
rect 17635 18173 17647 18176
rect 17589 18167 17647 18173
rect 18874 18164 18880 18176
rect 18932 18164 18938 18216
rect 18969 18207 19027 18213
rect 18969 18173 18981 18207
rect 19015 18204 19027 18207
rect 19628 18204 19656 18244
rect 19886 18232 19892 18244
rect 19944 18232 19950 18284
rect 21818 18232 21824 18284
rect 21876 18272 21882 18284
rect 23661 18275 23719 18281
rect 23661 18272 23673 18275
rect 21876 18244 23673 18272
rect 21876 18232 21882 18244
rect 23661 18241 23673 18244
rect 23707 18241 23719 18275
rect 23661 18235 23719 18241
rect 24302 18232 24308 18284
rect 24360 18272 24366 18284
rect 24871 18281 24899 18312
rect 25038 18300 25044 18312
rect 25096 18300 25102 18352
rect 29362 18340 29368 18352
rect 29323 18312 29368 18340
rect 29362 18300 29368 18312
rect 29420 18300 29426 18352
rect 30944 18312 31524 18340
rect 24443 18275 24501 18281
rect 24443 18272 24455 18275
rect 24360 18244 24455 18272
rect 24360 18232 24366 18244
rect 24443 18241 24455 18244
rect 24489 18241 24501 18275
rect 24673 18275 24731 18281
rect 24673 18272 24685 18275
rect 24443 18235 24501 18241
rect 24596 18244 24685 18272
rect 19015 18176 19656 18204
rect 19705 18207 19763 18213
rect 19015 18173 19027 18176
rect 18969 18167 19027 18173
rect 19705 18173 19717 18207
rect 19751 18173 19763 18207
rect 19705 18167 19763 18173
rect 19981 18207 20039 18213
rect 19981 18173 19993 18207
rect 20027 18204 20039 18207
rect 20438 18204 20444 18216
rect 20027 18176 20444 18204
rect 20027 18173 20039 18176
rect 19981 18167 20039 18173
rect 12986 18096 12992 18148
rect 13044 18136 13050 18148
rect 13446 18136 13452 18148
rect 13044 18108 13452 18136
rect 13044 18096 13050 18108
rect 13446 18096 13452 18108
rect 13504 18136 13510 18148
rect 17957 18139 18015 18145
rect 13504 18108 15332 18136
rect 13504 18096 13510 18108
rect 2225 18071 2283 18077
rect 2225 18037 2237 18071
rect 2271 18068 2283 18071
rect 5994 18068 6000 18080
rect 2271 18040 6000 18068
rect 2271 18037 2283 18040
rect 2225 18031 2283 18037
rect 5994 18028 6000 18040
rect 6052 18028 6058 18080
rect 7466 18028 7472 18080
rect 7524 18068 7530 18080
rect 8294 18068 8300 18080
rect 7524 18040 8300 18068
rect 7524 18028 7530 18040
rect 8294 18028 8300 18040
rect 8352 18028 8358 18080
rect 12802 18028 12808 18080
rect 12860 18068 12866 18080
rect 13081 18071 13139 18077
rect 13081 18068 13093 18071
rect 12860 18040 13093 18068
rect 12860 18028 12866 18040
rect 13081 18037 13093 18040
rect 13127 18037 13139 18071
rect 13081 18031 13139 18037
rect 15013 18071 15071 18077
rect 15013 18037 15025 18071
rect 15059 18068 15071 18071
rect 15194 18068 15200 18080
rect 15059 18040 15200 18068
rect 15059 18037 15071 18040
rect 15013 18031 15071 18037
rect 15194 18028 15200 18040
rect 15252 18028 15258 18080
rect 15304 18068 15332 18108
rect 17957 18105 17969 18139
rect 18003 18136 18015 18139
rect 19426 18136 19432 18148
rect 18003 18108 19432 18136
rect 18003 18105 18015 18108
rect 17957 18099 18015 18105
rect 19426 18096 19432 18108
rect 19484 18136 19490 18148
rect 19720 18136 19748 18167
rect 20438 18164 20444 18176
rect 20496 18164 20502 18216
rect 24210 18164 24216 18216
rect 24268 18204 24274 18216
rect 24596 18204 24624 18244
rect 24673 18241 24685 18244
rect 24719 18241 24731 18275
rect 24673 18235 24731 18241
rect 24856 18275 24914 18281
rect 24856 18241 24868 18275
rect 24902 18241 24914 18275
rect 24856 18235 24914 18241
rect 24946 18232 24952 18284
rect 25004 18272 25010 18284
rect 27801 18275 27859 18281
rect 25004 18244 25049 18272
rect 25004 18232 25010 18244
rect 27801 18241 27813 18275
rect 27847 18272 27859 18275
rect 28166 18272 28172 18284
rect 27847 18244 28172 18272
rect 27847 18241 27859 18244
rect 27801 18235 27859 18241
rect 28166 18232 28172 18244
rect 28224 18232 28230 18284
rect 28994 18232 29000 18284
rect 29052 18272 29058 18284
rect 29089 18275 29147 18281
rect 29089 18272 29101 18275
rect 29052 18244 29101 18272
rect 29052 18232 29058 18244
rect 29089 18241 29101 18244
rect 29135 18241 29147 18275
rect 30653 18275 30711 18281
rect 30653 18272 30665 18275
rect 29089 18235 29147 18241
rect 29380 18244 30665 18272
rect 25409 18207 25467 18213
rect 25409 18204 25421 18207
rect 24268 18176 25421 18204
rect 24268 18164 24274 18176
rect 25409 18173 25421 18176
rect 25455 18173 25467 18207
rect 25409 18167 25467 18173
rect 26970 18164 26976 18216
rect 27028 18204 27034 18216
rect 27525 18207 27583 18213
rect 27525 18204 27537 18207
rect 27028 18176 27537 18204
rect 27028 18164 27034 18176
rect 27525 18173 27537 18176
rect 27571 18173 27583 18207
rect 27525 18167 27583 18173
rect 29380 18145 29408 18244
rect 30653 18241 30665 18244
rect 30699 18241 30711 18275
rect 30944 18272 30972 18312
rect 30653 18235 30711 18241
rect 30760 18244 30972 18272
rect 29917 18207 29975 18213
rect 29917 18173 29929 18207
rect 29963 18204 29975 18207
rect 30377 18207 30435 18213
rect 30377 18204 30389 18207
rect 29963 18176 30389 18204
rect 29963 18173 29975 18176
rect 29917 18167 29975 18173
rect 30377 18173 30389 18176
rect 30423 18204 30435 18207
rect 30760 18204 30788 18244
rect 31018 18232 31024 18284
rect 31076 18272 31082 18284
rect 31386 18272 31392 18284
rect 31076 18244 31392 18272
rect 31076 18232 31082 18244
rect 31386 18232 31392 18244
rect 31444 18232 31450 18284
rect 31496 18272 31524 18312
rect 31754 18300 31760 18352
rect 31812 18340 31818 18352
rect 39393 18343 39451 18349
rect 31812 18312 37320 18340
rect 31812 18300 31818 18312
rect 32953 18275 33011 18281
rect 32953 18272 32965 18275
rect 31496 18244 32965 18272
rect 32953 18241 32965 18244
rect 32999 18272 33011 18275
rect 33318 18272 33324 18284
rect 32999 18244 33324 18272
rect 32999 18241 33011 18244
rect 32953 18235 33011 18241
rect 33318 18232 33324 18244
rect 33376 18232 33382 18284
rect 34330 18272 34336 18284
rect 34291 18244 34336 18272
rect 34330 18232 34336 18244
rect 34388 18232 34394 18284
rect 34422 18232 34428 18284
rect 34480 18272 34486 18284
rect 34609 18275 34667 18281
rect 34609 18272 34621 18275
rect 34480 18244 34621 18272
rect 34480 18232 34486 18244
rect 34609 18241 34621 18244
rect 34655 18241 34667 18275
rect 35986 18272 35992 18284
rect 35947 18244 35992 18272
rect 34609 18235 34667 18241
rect 35986 18232 35992 18244
rect 36044 18232 36050 18284
rect 36078 18232 36084 18284
rect 36136 18272 36142 18284
rect 37292 18281 37320 18312
rect 39393 18309 39405 18343
rect 39439 18340 39451 18343
rect 45741 18343 45799 18349
rect 39439 18312 43116 18340
rect 39439 18309 39451 18312
rect 39393 18303 39451 18309
rect 36265 18275 36323 18281
rect 36136 18244 36181 18272
rect 36136 18232 36142 18244
rect 36265 18241 36277 18275
rect 36311 18241 36323 18275
rect 36265 18235 36323 18241
rect 36357 18275 36415 18281
rect 36357 18241 36369 18275
rect 36403 18241 36415 18275
rect 36357 18235 36415 18241
rect 37277 18275 37335 18281
rect 37277 18241 37289 18275
rect 37323 18241 37335 18275
rect 37277 18235 37335 18241
rect 38749 18275 38807 18281
rect 38749 18241 38761 18275
rect 38795 18272 38807 18275
rect 38838 18272 38844 18284
rect 38795 18244 38844 18272
rect 38795 18241 38807 18244
rect 38749 18235 38807 18241
rect 30423 18176 30788 18204
rect 30837 18207 30895 18213
rect 30423 18173 30435 18176
rect 30377 18167 30435 18173
rect 30837 18173 30849 18207
rect 30883 18204 30895 18207
rect 30883 18176 35296 18204
rect 30883 18173 30895 18176
rect 30837 18167 30895 18173
rect 29365 18139 29423 18145
rect 19484 18108 19748 18136
rect 23400 18108 28994 18136
rect 19484 18096 19490 18108
rect 23400 18068 23428 18108
rect 15304 18040 23428 18068
rect 23474 18028 23480 18080
rect 23532 18068 23538 18080
rect 23569 18071 23627 18077
rect 23569 18068 23581 18071
rect 23532 18040 23581 18068
rect 23532 18028 23538 18040
rect 23569 18037 23581 18040
rect 23615 18037 23627 18071
rect 23569 18031 23627 18037
rect 24305 18071 24363 18077
rect 24305 18037 24317 18071
rect 24351 18068 24363 18071
rect 25682 18068 25688 18080
rect 24351 18040 25688 18068
rect 24351 18037 24363 18040
rect 24305 18031 24363 18037
rect 25682 18028 25688 18040
rect 25740 18028 25746 18080
rect 26970 18068 26976 18080
rect 26931 18040 26976 18068
rect 26970 18028 26976 18040
rect 27028 18028 27034 18080
rect 28966 18068 28994 18108
rect 29365 18105 29377 18139
rect 29411 18105 29423 18139
rect 29365 18099 29423 18105
rect 29932 18068 29960 18167
rect 32784 18108 32996 18136
rect 28966 18040 29960 18068
rect 30006 18028 30012 18080
rect 30064 18068 30070 18080
rect 30469 18071 30527 18077
rect 30469 18068 30481 18071
rect 30064 18040 30481 18068
rect 30064 18028 30070 18040
rect 30469 18037 30481 18040
rect 30515 18037 30527 18071
rect 31478 18068 31484 18080
rect 31391 18040 31484 18068
rect 30469 18031 30527 18037
rect 31478 18028 31484 18040
rect 31536 18068 31542 18080
rect 32784 18068 32812 18108
rect 31536 18040 32812 18068
rect 32968 18068 32996 18108
rect 33594 18096 33600 18148
rect 33652 18136 33658 18148
rect 34333 18139 34391 18145
rect 34333 18136 34345 18139
rect 33652 18108 34345 18136
rect 33652 18096 33658 18108
rect 34333 18105 34345 18108
rect 34379 18105 34391 18139
rect 34333 18099 34391 18105
rect 33962 18068 33968 18080
rect 32968 18040 33968 18068
rect 31536 18028 31542 18040
rect 33962 18028 33968 18040
rect 34020 18028 34026 18080
rect 35268 18068 35296 18176
rect 35710 18164 35716 18216
rect 35768 18204 35774 18216
rect 36280 18204 36308 18235
rect 35768 18176 36308 18204
rect 35768 18164 35774 18176
rect 35802 18096 35808 18148
rect 35860 18136 35866 18148
rect 36372 18136 36400 18235
rect 38838 18232 38844 18244
rect 38896 18232 38902 18284
rect 40310 18232 40316 18284
rect 40368 18272 40374 18284
rect 40497 18275 40555 18281
rect 40497 18272 40509 18275
rect 40368 18244 40509 18272
rect 40368 18232 40374 18244
rect 40497 18241 40509 18244
rect 40543 18241 40555 18275
rect 40678 18272 40684 18284
rect 40639 18244 40684 18272
rect 40497 18235 40555 18241
rect 40678 18232 40684 18244
rect 40736 18232 40742 18284
rect 43088 18272 43116 18312
rect 45741 18309 45753 18343
rect 45787 18340 45799 18343
rect 46014 18340 46020 18352
rect 45787 18312 46020 18340
rect 45787 18309 45799 18312
rect 45741 18303 45799 18309
rect 46014 18300 46020 18312
rect 46072 18300 46078 18352
rect 44726 18272 44732 18284
rect 43088 18244 44732 18272
rect 44726 18232 44732 18244
rect 44784 18272 44790 18284
rect 44784 18244 44850 18272
rect 44784 18232 44790 18244
rect 48774 18232 48780 18284
rect 48832 18272 48838 18284
rect 48869 18275 48927 18281
rect 48869 18272 48881 18275
rect 48832 18244 48881 18272
rect 48832 18232 48838 18244
rect 48869 18241 48881 18244
rect 48915 18241 48927 18275
rect 48869 18235 48927 18241
rect 48958 18232 48964 18284
rect 49016 18272 49022 18284
rect 49016 18244 49061 18272
rect 49016 18232 49022 18244
rect 49142 18232 49148 18284
rect 49200 18272 49206 18284
rect 53466 18272 53472 18284
rect 49200 18244 49245 18272
rect 53427 18244 53472 18272
rect 49200 18232 49206 18244
rect 53466 18232 53472 18244
rect 53524 18232 53530 18284
rect 53650 18272 53656 18284
rect 53611 18244 53656 18272
rect 53650 18232 53656 18244
rect 53708 18232 53714 18284
rect 56594 18272 56600 18284
rect 56555 18244 56600 18272
rect 56594 18232 56600 18244
rect 56652 18232 56658 18284
rect 56778 18272 56784 18284
rect 56739 18244 56784 18272
rect 56778 18232 56784 18244
rect 56836 18232 56842 18284
rect 57698 18232 57704 18284
rect 57756 18272 57762 18284
rect 57885 18275 57943 18281
rect 57885 18272 57897 18275
rect 57756 18244 57897 18272
rect 57756 18232 57762 18244
rect 57885 18241 57897 18244
rect 57931 18241 57943 18275
rect 57885 18235 57943 18241
rect 58069 18275 58127 18281
rect 58069 18241 58081 18275
rect 58115 18241 58127 18275
rect 58069 18235 58127 18241
rect 38473 18207 38531 18213
rect 38473 18204 38485 18207
rect 35860 18108 36400 18136
rect 36464 18176 38485 18204
rect 35860 18096 35866 18108
rect 36464 18068 36492 18176
rect 38473 18173 38485 18176
rect 38519 18173 38531 18207
rect 38473 18167 38531 18173
rect 44913 18207 44971 18213
rect 44913 18173 44925 18207
rect 44959 18173 44971 18207
rect 44913 18167 44971 18173
rect 36541 18139 36599 18145
rect 36541 18105 36553 18139
rect 36587 18136 36599 18139
rect 44928 18136 44956 18167
rect 57054 18164 57060 18216
rect 57112 18204 57118 18216
rect 57790 18204 57796 18216
rect 57112 18176 57796 18204
rect 57112 18164 57118 18176
rect 57790 18164 57796 18176
rect 57848 18204 57854 18216
rect 58084 18204 58112 18235
rect 57848 18176 58112 18204
rect 57848 18164 57854 18176
rect 45094 18136 45100 18148
rect 36587 18108 45100 18136
rect 36587 18105 36599 18108
rect 36541 18099 36599 18105
rect 45094 18096 45100 18108
rect 45152 18096 45158 18148
rect 37458 18068 37464 18080
rect 35268 18040 36492 18068
rect 37419 18040 37464 18068
rect 37458 18028 37464 18040
rect 37516 18028 37522 18080
rect 53193 18071 53251 18077
rect 53193 18037 53205 18071
rect 53239 18068 53251 18071
rect 53374 18068 53380 18080
rect 53239 18040 53380 18068
rect 53239 18037 53251 18040
rect 53193 18031 53251 18037
rect 53374 18028 53380 18040
rect 53432 18028 53438 18080
rect 1104 17978 58880 18000
rect 1104 17926 4214 17978
rect 4266 17926 4278 17978
rect 4330 17926 4342 17978
rect 4394 17926 4406 17978
rect 4458 17926 4470 17978
rect 4522 17926 34934 17978
rect 34986 17926 34998 17978
rect 35050 17926 35062 17978
rect 35114 17926 35126 17978
rect 35178 17926 35190 17978
rect 35242 17926 58880 17978
rect 1104 17904 58880 17926
rect 2685 17867 2743 17873
rect 2685 17833 2697 17867
rect 2731 17864 2743 17867
rect 3970 17864 3976 17876
rect 2731 17836 3976 17864
rect 2731 17833 2743 17836
rect 2685 17827 2743 17833
rect 3970 17824 3976 17836
rect 4028 17824 4034 17876
rect 7006 17864 7012 17876
rect 6967 17836 7012 17864
rect 7006 17824 7012 17836
rect 7064 17824 7070 17876
rect 7650 17864 7656 17876
rect 7611 17836 7656 17864
rect 7650 17824 7656 17836
rect 7708 17824 7714 17876
rect 8021 17867 8079 17873
rect 8021 17833 8033 17867
rect 8067 17864 8079 17867
rect 12618 17864 12624 17876
rect 8067 17836 12624 17864
rect 8067 17833 8079 17836
rect 8021 17827 8079 17833
rect 12618 17824 12624 17836
rect 12676 17824 12682 17876
rect 14458 17824 14464 17876
rect 14516 17864 14522 17876
rect 20714 17864 20720 17876
rect 14516 17836 20720 17864
rect 14516 17824 14522 17836
rect 20714 17824 20720 17836
rect 20772 17824 20778 17876
rect 21913 17867 21971 17873
rect 21913 17833 21925 17867
rect 21959 17864 21971 17867
rect 22094 17864 22100 17876
rect 21959 17836 22100 17864
rect 21959 17833 21971 17836
rect 21913 17827 21971 17833
rect 22094 17824 22100 17836
rect 22152 17824 22158 17876
rect 23198 17824 23204 17876
rect 23256 17864 23262 17876
rect 23750 17864 23756 17876
rect 23256 17836 23756 17864
rect 23256 17824 23262 17836
rect 23750 17824 23756 17836
rect 23808 17824 23814 17876
rect 24946 17864 24952 17876
rect 24907 17836 24952 17864
rect 24946 17824 24952 17836
rect 25004 17824 25010 17876
rect 27617 17867 27675 17873
rect 27617 17833 27629 17867
rect 27663 17864 27675 17867
rect 30190 17864 30196 17876
rect 27663 17836 30196 17864
rect 27663 17833 27675 17836
rect 27617 17827 27675 17833
rect 30190 17824 30196 17836
rect 30248 17824 30254 17876
rect 31849 17867 31907 17873
rect 31849 17833 31861 17867
rect 31895 17864 31907 17867
rect 33045 17867 33103 17873
rect 33045 17864 33057 17867
rect 31895 17836 33057 17864
rect 31895 17833 31907 17836
rect 31849 17827 31907 17833
rect 33045 17833 33057 17836
rect 33091 17864 33103 17867
rect 33226 17864 33232 17876
rect 33091 17836 33232 17864
rect 33091 17833 33103 17836
rect 33045 17827 33103 17833
rect 33226 17824 33232 17836
rect 33284 17824 33290 17876
rect 33410 17864 33416 17876
rect 33371 17836 33416 17864
rect 33410 17824 33416 17836
rect 33468 17824 33474 17876
rect 36173 17867 36231 17873
rect 36173 17833 36185 17867
rect 36219 17864 36231 17867
rect 36262 17864 36268 17876
rect 36219 17836 36268 17864
rect 36219 17833 36231 17836
rect 36173 17827 36231 17833
rect 36262 17824 36268 17836
rect 36320 17824 36326 17876
rect 45094 17864 45100 17876
rect 45055 17836 45100 17864
rect 45094 17824 45100 17836
rect 45152 17824 45158 17876
rect 48409 17867 48467 17873
rect 48409 17833 48421 17867
rect 48455 17864 48467 17867
rect 49694 17864 49700 17876
rect 48455 17836 49700 17864
rect 48455 17833 48467 17836
rect 48409 17827 48467 17833
rect 49694 17824 49700 17836
rect 49752 17824 49758 17876
rect 52730 17824 52736 17876
rect 52788 17864 52794 17876
rect 53466 17864 53472 17876
rect 52788 17836 53472 17864
rect 52788 17824 52794 17836
rect 53466 17824 53472 17836
rect 53524 17864 53530 17876
rect 53561 17867 53619 17873
rect 53561 17864 53573 17867
rect 53524 17836 53573 17864
rect 53524 17824 53530 17836
rect 53561 17833 53573 17836
rect 53607 17833 53619 17867
rect 56962 17864 56968 17876
rect 56923 17836 56968 17864
rect 53561 17827 53619 17833
rect 56962 17824 56968 17836
rect 57020 17824 57026 17876
rect 7190 17796 7196 17808
rect 7103 17768 7196 17796
rect 7190 17756 7196 17768
rect 7248 17796 7254 17808
rect 7248 17768 9168 17796
rect 7248 17756 7254 17768
rect 3970 17688 3976 17740
rect 4028 17728 4034 17740
rect 6181 17731 6239 17737
rect 4028 17700 5212 17728
rect 4028 17688 4034 17700
rect 4982 17660 4988 17672
rect 4943 17632 4988 17660
rect 4982 17620 4988 17632
rect 5040 17620 5046 17672
rect 5184 17669 5212 17700
rect 6181 17697 6193 17731
rect 6227 17728 6239 17731
rect 6227 17700 7880 17728
rect 6227 17697 6239 17700
rect 6181 17691 6239 17697
rect 5169 17663 5227 17669
rect 5169 17629 5181 17663
rect 5215 17629 5227 17663
rect 5169 17623 5227 17629
rect 5813 17663 5871 17669
rect 5813 17629 5825 17663
rect 5859 17629 5871 17663
rect 5994 17660 6000 17672
rect 5955 17632 6000 17660
rect 5813 17623 5871 17629
rect 1578 17552 1584 17604
rect 1636 17592 1642 17604
rect 2038 17592 2044 17604
rect 1636 17564 2044 17592
rect 1636 17552 1642 17564
rect 2038 17552 2044 17564
rect 2096 17592 2102 17604
rect 2409 17595 2467 17601
rect 2409 17592 2421 17595
rect 2096 17564 2421 17592
rect 2096 17552 2102 17564
rect 2409 17561 2421 17564
rect 2455 17561 2467 17595
rect 2409 17555 2467 17561
rect 5353 17595 5411 17601
rect 5353 17561 5365 17595
rect 5399 17592 5411 17595
rect 5828 17592 5856 17623
rect 5994 17620 6000 17632
rect 6052 17620 6058 17672
rect 6840 17601 6868 17700
rect 7653 17663 7711 17669
rect 7653 17629 7665 17663
rect 7699 17660 7711 17663
rect 7742 17660 7748 17672
rect 7699 17632 7748 17660
rect 7699 17629 7711 17632
rect 7653 17623 7711 17629
rect 7742 17620 7748 17632
rect 7800 17620 7806 17672
rect 7852 17669 7880 17700
rect 7837 17663 7895 17669
rect 7837 17629 7849 17663
rect 7883 17660 7895 17663
rect 8018 17660 8024 17672
rect 7883 17632 8024 17660
rect 7883 17629 7895 17632
rect 7837 17623 7895 17629
rect 8018 17620 8024 17632
rect 8076 17620 8082 17672
rect 9140 17669 9168 17768
rect 14366 17756 14372 17808
rect 14424 17796 14430 17808
rect 19978 17796 19984 17808
rect 14424 17768 19984 17796
rect 14424 17756 14430 17768
rect 19978 17756 19984 17768
rect 20036 17756 20042 17808
rect 24762 17796 24768 17808
rect 23308 17768 24768 17796
rect 12434 17688 12440 17740
rect 12492 17728 12498 17740
rect 13354 17728 13360 17740
rect 12492 17700 13360 17728
rect 12492 17688 12498 17700
rect 13354 17688 13360 17700
rect 13412 17688 13418 17740
rect 16666 17688 16672 17740
rect 16724 17728 16730 17740
rect 17589 17731 17647 17737
rect 17589 17728 17601 17731
rect 16724 17700 17601 17728
rect 16724 17688 16730 17700
rect 17589 17697 17601 17700
rect 17635 17728 17647 17731
rect 19426 17728 19432 17740
rect 17635 17700 19432 17728
rect 17635 17697 17647 17700
rect 17589 17691 17647 17697
rect 19426 17688 19432 17700
rect 19484 17688 19490 17740
rect 19705 17731 19763 17737
rect 19705 17697 19717 17731
rect 19751 17728 19763 17731
rect 20530 17728 20536 17740
rect 19751 17700 20536 17728
rect 19751 17697 19763 17700
rect 19705 17691 19763 17697
rect 20530 17688 20536 17700
rect 20588 17688 20594 17740
rect 8941 17663 8999 17669
rect 8941 17629 8953 17663
rect 8987 17629 8999 17663
rect 8941 17623 8999 17629
rect 9125 17663 9183 17669
rect 9125 17629 9137 17663
rect 9171 17629 9183 17663
rect 12618 17660 12624 17672
rect 12579 17632 12624 17660
rect 9125 17623 9183 17629
rect 6825 17595 6883 17601
rect 5399 17564 6040 17592
rect 5399 17561 5411 17564
rect 5353 17555 5411 17561
rect 6012 17524 6040 17564
rect 6825 17561 6837 17595
rect 6871 17561 6883 17595
rect 6825 17555 6883 17561
rect 7041 17595 7099 17601
rect 7041 17561 7053 17595
rect 7087 17592 7099 17595
rect 7282 17592 7288 17604
rect 7087 17564 7288 17592
rect 7087 17561 7099 17564
rect 7041 17555 7099 17561
rect 7282 17552 7288 17564
rect 7340 17552 7346 17604
rect 7760 17592 7788 17620
rect 8956 17592 8984 17623
rect 12618 17620 12624 17632
rect 12676 17620 12682 17672
rect 13722 17620 13728 17672
rect 13780 17660 13786 17672
rect 14277 17663 14335 17669
rect 14277 17660 14289 17663
rect 13780 17632 14289 17660
rect 13780 17620 13786 17632
rect 14277 17629 14289 17632
rect 14323 17629 14335 17663
rect 15194 17660 15200 17672
rect 15155 17632 15200 17660
rect 14277 17623 14335 17629
rect 15194 17620 15200 17632
rect 15252 17620 15258 17672
rect 17773 17663 17831 17669
rect 17773 17629 17785 17663
rect 17819 17660 17831 17663
rect 18506 17660 18512 17672
rect 17819 17632 18512 17660
rect 17819 17629 17831 17632
rect 17773 17623 17831 17629
rect 18506 17620 18512 17632
rect 18564 17620 18570 17672
rect 18598 17620 18604 17672
rect 18656 17660 18662 17672
rect 19521 17663 19579 17669
rect 19521 17660 19533 17663
rect 18656 17632 19533 17660
rect 18656 17620 18662 17632
rect 19521 17629 19533 17632
rect 19567 17629 19579 17663
rect 19521 17623 19579 17629
rect 20070 17620 20076 17672
rect 20128 17660 20134 17672
rect 20165 17663 20223 17669
rect 20165 17660 20177 17663
rect 20128 17632 20177 17660
rect 20128 17620 20134 17632
rect 20165 17629 20177 17632
rect 20211 17629 20223 17663
rect 20165 17623 20223 17629
rect 20258 17663 20316 17669
rect 20258 17629 20270 17663
rect 20304 17629 20316 17663
rect 20258 17623 20316 17629
rect 15010 17592 15016 17604
rect 7760 17564 8984 17592
rect 14971 17564 15016 17592
rect 15010 17552 15016 17564
rect 15068 17552 15074 17604
rect 15562 17592 15568 17604
rect 15523 17564 15568 17592
rect 15562 17552 15568 17564
rect 15620 17552 15626 17604
rect 18230 17552 18236 17604
rect 18288 17592 18294 17604
rect 20272 17592 20300 17623
rect 20622 17620 20628 17672
rect 20680 17669 20686 17672
rect 20680 17660 20688 17669
rect 20680 17632 20725 17660
rect 20680 17623 20688 17632
rect 20680 17620 20686 17623
rect 21910 17620 21916 17672
rect 21968 17660 21974 17672
rect 23308 17669 23336 17768
rect 24762 17756 24768 17768
rect 24820 17756 24826 17808
rect 36078 17756 36084 17808
rect 36136 17796 36142 17808
rect 36357 17799 36415 17805
rect 36357 17796 36369 17799
rect 36136 17768 36369 17796
rect 36136 17756 36142 17768
rect 36357 17765 36369 17768
rect 36403 17765 36415 17799
rect 36357 17759 36415 17765
rect 41325 17799 41383 17805
rect 41325 17765 41337 17799
rect 41371 17796 41383 17799
rect 41690 17796 41696 17808
rect 41371 17768 41696 17796
rect 41371 17765 41383 17768
rect 41325 17759 41383 17765
rect 41690 17756 41696 17768
rect 41748 17756 41754 17808
rect 24670 17688 24676 17740
rect 24728 17688 24734 17740
rect 26234 17688 26240 17740
rect 26292 17728 26298 17740
rect 26973 17731 27031 17737
rect 26973 17728 26985 17731
rect 26292 17700 26985 17728
rect 26292 17688 26298 17700
rect 26973 17697 26985 17700
rect 27019 17697 27031 17731
rect 26973 17691 27031 17697
rect 40218 17688 40224 17740
rect 40276 17728 40282 17740
rect 40865 17731 40923 17737
rect 40865 17728 40877 17731
rect 40276 17700 40877 17728
rect 40276 17688 40282 17700
rect 40865 17697 40877 17700
rect 40911 17697 40923 17731
rect 40865 17691 40923 17697
rect 43990 17688 43996 17740
rect 44048 17728 44054 17740
rect 44269 17731 44327 17737
rect 44269 17728 44281 17731
rect 44048 17700 44281 17728
rect 44048 17688 44054 17700
rect 44269 17697 44281 17700
rect 44315 17697 44327 17731
rect 44269 17691 44327 17697
rect 44453 17731 44511 17737
rect 44453 17697 44465 17731
rect 44499 17728 44511 17731
rect 45370 17728 45376 17740
rect 44499 17700 45376 17728
rect 44499 17697 44511 17700
rect 44453 17691 44511 17697
rect 45370 17688 45376 17700
rect 45428 17728 45434 17740
rect 45465 17731 45523 17737
rect 45465 17728 45477 17731
rect 45428 17700 45477 17728
rect 45428 17688 45434 17700
rect 45465 17697 45477 17700
rect 45511 17697 45523 17731
rect 53650 17728 53656 17740
rect 53611 17700 53656 17728
rect 45465 17691 45523 17697
rect 53650 17688 53656 17700
rect 53708 17688 53714 17740
rect 57054 17728 57060 17740
rect 57015 17700 57060 17728
rect 57054 17688 57060 17700
rect 57112 17688 57118 17740
rect 22649 17663 22707 17669
rect 22649 17660 22661 17663
rect 21968 17632 22661 17660
rect 21968 17620 21974 17632
rect 22649 17629 22661 17632
rect 22695 17629 22707 17663
rect 22649 17623 22707 17629
rect 23293 17663 23351 17669
rect 23293 17629 23305 17663
rect 23339 17629 23351 17663
rect 23293 17623 23351 17629
rect 23661 17663 23719 17669
rect 23661 17629 23673 17663
rect 23707 17660 23719 17663
rect 23750 17660 23756 17672
rect 23707 17632 23756 17660
rect 23707 17629 23719 17632
rect 23661 17623 23719 17629
rect 20438 17592 20444 17604
rect 18288 17564 20300 17592
rect 20399 17564 20444 17592
rect 18288 17552 18294 17564
rect 20438 17552 20444 17564
rect 20496 17552 20502 17604
rect 20533 17595 20591 17601
rect 20533 17561 20545 17595
rect 20579 17592 20591 17595
rect 20714 17592 20720 17604
rect 20579 17564 20720 17592
rect 20579 17561 20591 17564
rect 20533 17555 20591 17561
rect 20714 17552 20720 17564
rect 20772 17552 20778 17604
rect 22005 17595 22063 17601
rect 22005 17561 22017 17595
rect 22051 17592 22063 17595
rect 23308 17592 23336 17623
rect 23750 17620 23756 17632
rect 23808 17620 23814 17672
rect 24397 17663 24455 17669
rect 24397 17629 24409 17663
rect 24443 17660 24455 17663
rect 24688 17660 24716 17688
rect 24443 17632 24716 17660
rect 24765 17663 24823 17669
rect 24443 17629 24455 17632
rect 24397 17623 24455 17629
rect 24765 17629 24777 17663
rect 24811 17660 24823 17663
rect 24854 17660 24860 17672
rect 24811 17632 24860 17660
rect 24811 17629 24823 17632
rect 24765 17623 24823 17629
rect 23474 17592 23480 17604
rect 22051 17564 23336 17592
rect 23435 17564 23480 17592
rect 22051 17561 22063 17564
rect 22005 17555 22063 17561
rect 23474 17552 23480 17564
rect 23532 17552 23538 17604
rect 23569 17595 23627 17601
rect 23569 17561 23581 17595
rect 23615 17592 23627 17595
rect 24412 17592 24440 17623
rect 24854 17620 24860 17632
rect 24912 17620 24918 17672
rect 25869 17663 25927 17669
rect 25869 17629 25881 17663
rect 25915 17660 25927 17663
rect 26418 17660 26424 17672
rect 25915 17632 26424 17660
rect 25915 17629 25927 17632
rect 25869 17623 25927 17629
rect 26418 17620 26424 17632
rect 26476 17660 26482 17672
rect 27157 17663 27215 17669
rect 27157 17660 27169 17663
rect 26476 17632 27169 17660
rect 26476 17620 26482 17632
rect 27157 17629 27169 17632
rect 27203 17660 27215 17663
rect 28169 17663 28227 17669
rect 28169 17660 28181 17663
rect 27203 17632 28181 17660
rect 27203 17629 27215 17632
rect 27157 17623 27215 17629
rect 28169 17629 28181 17632
rect 28215 17660 28227 17663
rect 28813 17663 28871 17669
rect 28813 17660 28825 17663
rect 28215 17632 28825 17660
rect 28215 17629 28227 17632
rect 28169 17623 28227 17629
rect 28813 17629 28825 17632
rect 28859 17629 28871 17663
rect 28813 17623 28871 17629
rect 30009 17663 30067 17669
rect 30009 17629 30021 17663
rect 30055 17660 30067 17663
rect 30098 17660 30104 17672
rect 30055 17632 30104 17660
rect 30055 17629 30067 17632
rect 30009 17623 30067 17629
rect 30098 17620 30104 17632
rect 30156 17620 30162 17672
rect 30650 17660 30656 17672
rect 30611 17632 30656 17660
rect 30650 17620 30656 17632
rect 30708 17620 30714 17672
rect 32309 17663 32367 17669
rect 32309 17629 32321 17663
rect 32355 17660 32367 17663
rect 32398 17660 32404 17672
rect 32355 17632 32404 17660
rect 32355 17629 32367 17632
rect 32309 17623 32367 17629
rect 32398 17620 32404 17632
rect 32456 17620 32462 17672
rect 33045 17663 33103 17669
rect 33045 17629 33057 17663
rect 33091 17629 33103 17663
rect 33045 17623 33103 17629
rect 33229 17663 33287 17669
rect 33229 17629 33241 17663
rect 33275 17660 33287 17663
rect 33410 17660 33416 17672
rect 33275 17632 33416 17660
rect 33275 17629 33287 17632
rect 33229 17623 33287 17629
rect 24578 17592 24584 17604
rect 23615 17564 24440 17592
rect 24539 17564 24584 17592
rect 23615 17561 23627 17564
rect 23569 17555 23627 17561
rect 24578 17552 24584 17564
rect 24636 17552 24642 17604
rect 24673 17595 24731 17601
rect 24673 17561 24685 17595
rect 24719 17592 24731 17595
rect 24946 17592 24952 17604
rect 24719 17564 24952 17592
rect 24719 17561 24731 17564
rect 24673 17555 24731 17561
rect 24946 17552 24952 17564
rect 25004 17592 25010 17604
rect 25958 17592 25964 17604
rect 25004 17564 25964 17592
rect 25004 17552 25010 17564
rect 25958 17552 25964 17564
rect 26016 17552 26022 17604
rect 26970 17592 26976 17604
rect 26344 17564 26976 17592
rect 26344 17536 26372 17564
rect 26970 17552 26976 17564
rect 27028 17592 27034 17604
rect 27249 17595 27307 17601
rect 27249 17592 27261 17595
rect 27028 17564 27261 17592
rect 27028 17552 27034 17564
rect 27249 17561 27261 17564
rect 27295 17561 27307 17595
rect 27249 17555 27307 17561
rect 28626 17552 28632 17604
rect 28684 17592 28690 17604
rect 30193 17595 30251 17601
rect 30193 17592 30205 17595
rect 28684 17564 30205 17592
rect 28684 17552 28690 17564
rect 30193 17561 30205 17564
rect 30239 17561 30251 17595
rect 30193 17555 30251 17561
rect 32582 17552 32588 17604
rect 32640 17592 32646 17604
rect 33060 17592 33088 17623
rect 33410 17620 33416 17632
rect 33468 17620 33474 17672
rect 40494 17620 40500 17672
rect 40552 17660 40558 17672
rect 40957 17663 41015 17669
rect 40957 17660 40969 17663
rect 40552 17632 40969 17660
rect 40552 17620 40558 17632
rect 40957 17629 40969 17632
rect 41003 17629 41015 17663
rect 44174 17660 44180 17672
rect 44135 17632 44180 17660
rect 40957 17623 41015 17629
rect 44174 17620 44180 17632
rect 44232 17620 44238 17672
rect 44726 17620 44732 17672
rect 44784 17660 44790 17672
rect 45005 17663 45063 17669
rect 45005 17660 45017 17663
rect 44784 17632 45017 17660
rect 44784 17620 44790 17632
rect 45005 17629 45017 17632
rect 45051 17629 45063 17663
rect 48225 17663 48283 17669
rect 48225 17660 48237 17663
rect 45005 17623 45063 17629
rect 45526 17632 48237 17660
rect 33873 17595 33931 17601
rect 33873 17592 33885 17595
rect 32640 17564 33885 17592
rect 32640 17552 32646 17564
rect 33873 17561 33885 17564
rect 33919 17561 33931 17595
rect 33873 17555 33931 17561
rect 35894 17552 35900 17604
rect 35952 17592 35958 17604
rect 35989 17595 36047 17601
rect 35989 17592 36001 17595
rect 35952 17564 36001 17592
rect 35952 17552 35958 17564
rect 35989 17561 36001 17564
rect 36035 17561 36047 17595
rect 35989 17555 36047 17561
rect 36205 17595 36263 17601
rect 36205 17561 36217 17595
rect 36251 17592 36263 17595
rect 36538 17592 36544 17604
rect 36251 17564 36544 17592
rect 36251 17561 36263 17564
rect 36205 17555 36263 17561
rect 36538 17552 36544 17564
rect 36596 17592 36602 17604
rect 36909 17595 36967 17601
rect 36909 17592 36921 17595
rect 36596 17564 36921 17592
rect 36596 17552 36602 17564
rect 36909 17561 36921 17564
rect 36955 17592 36967 17595
rect 44082 17592 44088 17604
rect 36955 17564 44088 17592
rect 36955 17561 36967 17564
rect 36909 17555 36967 17561
rect 44082 17552 44088 17564
rect 44140 17552 44146 17604
rect 44453 17595 44511 17601
rect 44453 17561 44465 17595
rect 44499 17592 44511 17595
rect 45526 17592 45554 17632
rect 48225 17629 48237 17632
rect 48271 17660 48283 17663
rect 48958 17660 48964 17672
rect 48271 17632 48964 17660
rect 48271 17629 48283 17632
rect 48225 17623 48283 17629
rect 48958 17620 48964 17632
rect 49016 17660 49022 17672
rect 49329 17663 49387 17669
rect 49329 17660 49341 17663
rect 49016 17632 49341 17660
rect 49016 17620 49022 17632
rect 49329 17629 49341 17632
rect 49375 17629 49387 17663
rect 49329 17623 49387 17629
rect 49421 17663 49479 17669
rect 49421 17629 49433 17663
rect 49467 17629 49479 17663
rect 49421 17623 49479 17629
rect 48314 17592 48320 17604
rect 44499 17564 45554 17592
rect 48275 17564 48320 17592
rect 44499 17561 44511 17564
rect 44453 17555 44511 17561
rect 48314 17552 48320 17564
rect 48372 17552 48378 17604
rect 48498 17592 48504 17604
rect 48459 17564 48504 17592
rect 48498 17552 48504 17564
rect 48556 17592 48562 17604
rect 49142 17592 49148 17604
rect 48556 17564 49148 17592
rect 48556 17552 48562 17564
rect 49142 17552 49148 17564
rect 49200 17592 49206 17604
rect 49436 17592 49464 17623
rect 53374 17620 53380 17672
rect 53432 17660 53438 17672
rect 53929 17663 53987 17669
rect 53929 17660 53941 17663
rect 53432 17632 53941 17660
rect 53432 17620 53438 17632
rect 53929 17629 53941 17632
rect 53975 17629 53987 17663
rect 53929 17623 53987 17629
rect 56686 17620 56692 17672
rect 56744 17660 56750 17672
rect 56781 17663 56839 17669
rect 56781 17660 56793 17663
rect 56744 17632 56793 17660
rect 56744 17620 56750 17632
rect 56781 17629 56793 17632
rect 56827 17629 56839 17663
rect 56781 17623 56839 17629
rect 56873 17663 56931 17669
rect 56873 17629 56885 17663
rect 56919 17660 56931 17663
rect 56962 17660 56968 17672
rect 56919 17632 56968 17660
rect 56919 17629 56931 17632
rect 56873 17623 56931 17629
rect 56962 17620 56968 17632
rect 57020 17620 57026 17672
rect 58066 17660 58072 17672
rect 58027 17632 58072 17660
rect 58066 17620 58072 17632
rect 58124 17620 58130 17672
rect 49200 17564 49464 17592
rect 49200 17552 49206 17564
rect 56318 17552 56324 17604
rect 56376 17592 56382 17604
rect 57701 17595 57759 17601
rect 57701 17592 57713 17595
rect 56376 17564 57713 17592
rect 56376 17552 56382 17564
rect 57701 17561 57713 17564
rect 57747 17561 57759 17595
rect 57701 17555 57759 17561
rect 8202 17524 8208 17536
rect 6012 17496 8208 17524
rect 8202 17484 8208 17496
rect 8260 17484 8266 17536
rect 8938 17524 8944 17536
rect 8899 17496 8944 17524
rect 8938 17484 8944 17496
rect 8996 17484 9002 17536
rect 12805 17527 12863 17533
rect 12805 17493 12817 17527
rect 12851 17524 12863 17527
rect 13998 17524 14004 17536
rect 12851 17496 14004 17524
rect 12851 17493 12863 17496
rect 12805 17487 12863 17493
rect 13998 17484 14004 17496
rect 14056 17484 14062 17536
rect 14461 17527 14519 17533
rect 14461 17493 14473 17527
rect 14507 17524 14519 17527
rect 16942 17524 16948 17536
rect 14507 17496 16948 17524
rect 14507 17493 14519 17496
rect 14461 17487 14519 17493
rect 16942 17484 16948 17496
rect 17000 17484 17006 17536
rect 18322 17524 18328 17536
rect 18283 17496 18328 17524
rect 18322 17484 18328 17496
rect 18380 17484 18386 17536
rect 20806 17524 20812 17536
rect 20767 17496 20812 17524
rect 20806 17484 20812 17496
rect 20864 17484 20870 17536
rect 22741 17527 22799 17533
rect 22741 17493 22753 17527
rect 22787 17524 22799 17527
rect 23198 17524 23204 17536
rect 22787 17496 23204 17524
rect 22787 17493 22799 17496
rect 22741 17487 22799 17493
rect 23198 17484 23204 17496
rect 23256 17484 23262 17536
rect 23842 17524 23848 17536
rect 23803 17496 23848 17524
rect 23842 17484 23848 17496
rect 23900 17484 23906 17536
rect 26326 17524 26332 17536
rect 26287 17496 26332 17524
rect 26326 17484 26332 17496
rect 26384 17484 26390 17536
rect 28261 17527 28319 17533
rect 28261 17493 28273 17527
rect 28307 17524 28319 17527
rect 28718 17524 28724 17536
rect 28307 17496 28724 17524
rect 28307 17493 28319 17496
rect 28261 17487 28319 17493
rect 28718 17484 28724 17496
rect 28776 17484 28782 17536
rect 30834 17524 30840 17536
rect 30795 17496 30840 17524
rect 30834 17484 30840 17496
rect 30892 17484 30898 17536
rect 32493 17527 32551 17533
rect 32493 17493 32505 17527
rect 32539 17524 32551 17527
rect 33778 17524 33784 17536
rect 32539 17496 33784 17524
rect 32539 17493 32551 17496
rect 32493 17487 32551 17493
rect 33778 17484 33784 17496
rect 33836 17524 33842 17536
rect 34422 17524 34428 17536
rect 33836 17496 34428 17524
rect 33836 17484 33842 17496
rect 34422 17484 34428 17496
rect 34480 17484 34486 17536
rect 40218 17524 40224 17536
rect 40179 17496 40224 17524
rect 40218 17484 40224 17496
rect 40276 17484 40282 17536
rect 48332 17524 48360 17552
rect 48774 17524 48780 17536
rect 48332 17496 48780 17524
rect 48774 17484 48780 17496
rect 48832 17524 48838 17536
rect 48961 17527 49019 17533
rect 48961 17524 48973 17527
rect 48832 17496 48973 17524
rect 48832 17484 48838 17496
rect 48961 17493 48973 17496
rect 49007 17493 49019 17527
rect 48961 17487 49019 17493
rect 49605 17527 49663 17533
rect 49605 17493 49617 17527
rect 49651 17524 49663 17527
rect 52546 17524 52552 17536
rect 49651 17496 52552 17524
rect 49651 17493 49663 17496
rect 49605 17487 49663 17493
rect 52546 17484 52552 17496
rect 52604 17484 52610 17536
rect 53377 17527 53435 17533
rect 53377 17493 53389 17527
rect 53423 17524 53435 17527
rect 53558 17524 53564 17536
rect 53423 17496 53564 17524
rect 53423 17493 53435 17496
rect 53377 17487 53435 17493
rect 53558 17484 53564 17496
rect 53616 17484 53622 17536
rect 1104 17434 58880 17456
rect 1104 17382 19574 17434
rect 19626 17382 19638 17434
rect 19690 17382 19702 17434
rect 19754 17382 19766 17434
rect 19818 17382 19830 17434
rect 19882 17382 50294 17434
rect 50346 17382 50358 17434
rect 50410 17382 50422 17434
rect 50474 17382 50486 17434
rect 50538 17382 50550 17434
rect 50602 17382 58880 17434
rect 1104 17360 58880 17382
rect 3050 17280 3056 17332
rect 3108 17320 3114 17332
rect 3329 17323 3387 17329
rect 3329 17320 3341 17323
rect 3108 17292 3341 17320
rect 3108 17280 3114 17292
rect 3329 17289 3341 17292
rect 3375 17320 3387 17323
rect 3510 17320 3516 17332
rect 3375 17292 3516 17320
rect 3375 17289 3387 17292
rect 3329 17283 3387 17289
rect 3510 17280 3516 17292
rect 3568 17280 3574 17332
rect 8323 17323 8381 17329
rect 8323 17289 8335 17323
rect 8369 17320 8381 17323
rect 8938 17320 8944 17332
rect 8369 17292 8944 17320
rect 8369 17289 8381 17292
rect 8323 17283 8381 17289
rect 8938 17280 8944 17292
rect 8996 17280 9002 17332
rect 9122 17280 9128 17332
rect 9180 17320 9186 17332
rect 16574 17320 16580 17332
rect 9180 17292 16580 17320
rect 9180 17280 9186 17292
rect 16574 17280 16580 17292
rect 16632 17280 16638 17332
rect 20070 17320 20076 17332
rect 20031 17292 20076 17320
rect 20070 17280 20076 17292
rect 20128 17280 20134 17332
rect 20346 17280 20352 17332
rect 20404 17280 20410 17332
rect 24578 17280 24584 17332
rect 24636 17320 24642 17332
rect 28350 17320 28356 17332
rect 24636 17292 28356 17320
rect 24636 17280 24642 17292
rect 28350 17280 28356 17292
rect 28408 17320 28414 17332
rect 28408 17292 28580 17320
rect 28408 17280 28414 17292
rect 4982 17212 4988 17264
rect 5040 17252 5046 17264
rect 7466 17252 7472 17264
rect 5040 17224 7472 17252
rect 5040 17212 5046 17224
rect 7466 17212 7472 17224
rect 7524 17212 7530 17264
rect 7653 17255 7711 17261
rect 7653 17221 7665 17255
rect 7699 17252 7711 17255
rect 8018 17252 8024 17264
rect 7699 17224 8024 17252
rect 7699 17221 7711 17224
rect 7653 17215 7711 17221
rect 8018 17212 8024 17224
rect 8076 17212 8082 17264
rect 8113 17255 8171 17261
rect 8113 17221 8125 17255
rect 8159 17252 8171 17255
rect 8202 17252 8208 17264
rect 8159 17224 8208 17252
rect 8159 17221 8171 17224
rect 8113 17215 8171 17221
rect 8202 17212 8208 17224
rect 8260 17212 8266 17264
rect 9033 17255 9091 17261
rect 9033 17221 9045 17255
rect 9079 17252 9091 17255
rect 10410 17252 10416 17264
rect 9079 17224 10416 17252
rect 9079 17221 9091 17224
rect 9033 17215 9091 17221
rect 10410 17212 10416 17224
rect 10468 17252 10474 17264
rect 10468 17224 10824 17252
rect 10468 17212 10474 17224
rect 8941 17187 8999 17193
rect 8941 17184 8953 17187
rect 8312 17156 8953 17184
rect 2866 17116 2872 17128
rect 2827 17088 2872 17116
rect 2866 17076 2872 17088
rect 2924 17076 2930 17128
rect 7282 17116 7288 17128
rect 7195 17088 7288 17116
rect 7282 17076 7288 17088
rect 7340 17116 7346 17128
rect 8312 17116 8340 17156
rect 8941 17153 8953 17156
rect 8987 17153 8999 17187
rect 9125 17187 9183 17193
rect 9125 17184 9137 17187
rect 8941 17147 8999 17153
rect 9048 17156 9137 17184
rect 9048 17128 9076 17156
rect 9125 17153 9137 17156
rect 9171 17153 9183 17187
rect 9950 17184 9956 17196
rect 9911 17156 9956 17184
rect 9125 17147 9183 17153
rect 9950 17144 9956 17156
rect 10008 17144 10014 17196
rect 10134 17144 10140 17196
rect 10192 17184 10198 17196
rect 10796 17193 10824 17224
rect 12894 17212 12900 17264
rect 12952 17252 12958 17264
rect 13722 17252 13728 17264
rect 12952 17224 13728 17252
rect 12952 17212 12958 17224
rect 13722 17212 13728 17224
rect 13780 17252 13786 17264
rect 14277 17255 14335 17261
rect 14277 17252 14289 17255
rect 13780 17224 14289 17252
rect 13780 17212 13786 17224
rect 14277 17221 14289 17224
rect 14323 17252 14335 17255
rect 20364 17252 20392 17280
rect 21177 17255 21235 17261
rect 21177 17252 21189 17255
rect 14323 17224 15516 17252
rect 14323 17221 14335 17224
rect 14277 17215 14335 17221
rect 10229 17187 10287 17193
rect 10229 17184 10241 17187
rect 10192 17156 10241 17184
rect 10192 17144 10198 17156
rect 10229 17153 10241 17156
rect 10275 17153 10287 17187
rect 10229 17147 10287 17153
rect 10781 17187 10839 17193
rect 10781 17153 10793 17187
rect 10827 17153 10839 17187
rect 14090 17184 14096 17196
rect 14051 17156 14096 17184
rect 10781 17147 10839 17153
rect 14090 17144 14096 17156
rect 14148 17144 14154 17196
rect 14366 17184 14372 17196
rect 14279 17156 14372 17184
rect 14366 17144 14372 17156
rect 14424 17144 14430 17196
rect 14461 17187 14519 17193
rect 14461 17153 14473 17187
rect 14507 17184 14519 17187
rect 14550 17184 14556 17196
rect 14507 17156 14556 17184
rect 14507 17153 14519 17156
rect 14461 17147 14519 17153
rect 14550 17144 14556 17156
rect 14608 17144 14614 17196
rect 14734 17144 14740 17196
rect 14792 17184 14798 17196
rect 15105 17187 15163 17193
rect 15105 17184 15117 17187
rect 14792 17156 15117 17184
rect 14792 17144 14798 17156
rect 15105 17153 15117 17156
rect 15151 17153 15163 17187
rect 15105 17147 15163 17153
rect 15194 17144 15200 17196
rect 15252 17184 15258 17196
rect 15488 17193 15516 17224
rect 18248 17224 19840 17252
rect 20364 17224 21189 17252
rect 18248 17193 18276 17224
rect 15289 17187 15347 17193
rect 15289 17184 15301 17187
rect 15252 17156 15301 17184
rect 15252 17144 15258 17156
rect 15289 17153 15301 17156
rect 15335 17153 15347 17187
rect 15289 17147 15347 17153
rect 15381 17187 15439 17193
rect 15381 17153 15393 17187
rect 15427 17153 15439 17187
rect 15381 17147 15439 17153
rect 15473 17187 15531 17193
rect 15473 17153 15485 17187
rect 15519 17153 15531 17187
rect 15473 17147 15531 17153
rect 18233 17187 18291 17193
rect 18233 17153 18245 17187
rect 18279 17153 18291 17187
rect 18233 17147 18291 17153
rect 7340 17088 8340 17116
rect 7340 17076 7346 17088
rect 9030 17076 9036 17128
rect 9088 17076 9094 17128
rect 9968 17116 9996 17144
rect 12434 17116 12440 17128
rect 9968 17088 12440 17116
rect 12434 17076 12440 17088
rect 12492 17076 12498 17128
rect 13633 17119 13691 17125
rect 13633 17085 13645 17119
rect 13679 17116 13691 17119
rect 14384 17116 14412 17144
rect 13679 17088 14412 17116
rect 13679 17085 13691 17088
rect 13633 17079 13691 17085
rect 3237 17051 3295 17057
rect 3237 17017 3249 17051
rect 3283 17048 3295 17051
rect 3418 17048 3424 17060
rect 3283 17020 3424 17048
rect 3283 17017 3295 17020
rect 3237 17011 3295 17017
rect 3418 17008 3424 17020
rect 3476 17008 3482 17060
rect 8202 17008 8208 17060
rect 8260 17048 8266 17060
rect 10873 17051 10931 17057
rect 8260 17020 9674 17048
rect 8260 17008 8266 17020
rect 1673 16983 1731 16989
rect 1673 16949 1685 16983
rect 1719 16980 1731 16983
rect 1854 16980 1860 16992
rect 1719 16952 1860 16980
rect 1719 16949 1731 16952
rect 1673 16943 1731 16949
rect 1854 16940 1860 16952
rect 1912 16940 1918 16992
rect 7834 16940 7840 16992
rect 7892 16980 7898 16992
rect 8297 16983 8355 16989
rect 8297 16980 8309 16983
rect 7892 16952 8309 16980
rect 7892 16940 7898 16952
rect 8297 16949 8309 16952
rect 8343 16949 8355 16983
rect 8478 16980 8484 16992
rect 8439 16952 8484 16980
rect 8297 16943 8355 16949
rect 8478 16940 8484 16952
rect 8536 16940 8542 16992
rect 9646 16980 9674 17020
rect 10873 17017 10885 17051
rect 10919 17048 10931 17051
rect 15286 17048 15292 17060
rect 10919 17020 15292 17048
rect 10919 17017 10931 17020
rect 10873 17011 10931 17017
rect 15286 17008 15292 17020
rect 15344 17008 15350 17060
rect 15396 17048 15424 17147
rect 17954 17048 17960 17060
rect 15396 17020 17960 17048
rect 17954 17008 17960 17020
rect 18012 17048 18018 17060
rect 18049 17051 18107 17057
rect 18049 17048 18061 17051
rect 18012 17020 18061 17048
rect 18012 17008 18018 17020
rect 18049 17017 18061 17020
rect 18095 17017 18107 17051
rect 19352 17048 19380 17224
rect 19518 17184 19524 17196
rect 19479 17156 19524 17184
rect 19518 17144 19524 17156
rect 19576 17144 19582 17196
rect 19702 17184 19708 17196
rect 19663 17156 19708 17184
rect 19702 17144 19708 17156
rect 19760 17144 19766 17196
rect 19812 17193 19840 17224
rect 19797 17187 19855 17193
rect 19797 17153 19809 17187
rect 19843 17153 19855 17187
rect 19797 17147 19855 17153
rect 19889 17187 19947 17193
rect 19889 17153 19901 17187
rect 19935 17184 19947 17187
rect 20162 17184 20168 17196
rect 19935 17156 20168 17184
rect 19935 17153 19947 17156
rect 19889 17147 19947 17153
rect 20162 17144 20168 17156
rect 20220 17184 20226 17196
rect 20346 17184 20352 17196
rect 20220 17156 20352 17184
rect 20220 17144 20226 17156
rect 20346 17144 20352 17156
rect 20404 17144 20410 17196
rect 20530 17184 20536 17196
rect 20491 17156 20536 17184
rect 20530 17144 20536 17156
rect 20588 17144 20594 17196
rect 20732 17193 20760 17224
rect 21177 17221 21189 17224
rect 21223 17221 21235 17255
rect 21177 17215 21235 17221
rect 22738 17212 22744 17264
rect 22796 17252 22802 17264
rect 23753 17255 23811 17261
rect 23753 17252 23765 17255
rect 22796 17224 23765 17252
rect 22796 17212 22802 17224
rect 23753 17221 23765 17224
rect 23799 17221 23811 17255
rect 24670 17252 24676 17264
rect 24631 17224 24676 17252
rect 23753 17215 23811 17221
rect 24670 17212 24676 17224
rect 24728 17212 24734 17264
rect 24854 17212 24860 17264
rect 24912 17252 24918 17264
rect 25961 17255 26019 17261
rect 25961 17252 25973 17255
rect 24912 17224 25973 17252
rect 24912 17212 24918 17224
rect 25961 17221 25973 17224
rect 26007 17221 26019 17255
rect 25961 17215 26019 17221
rect 20717 17187 20775 17193
rect 20717 17153 20729 17187
rect 20763 17153 20775 17187
rect 20717 17147 20775 17153
rect 24302 17144 24308 17196
rect 24360 17184 24366 17196
rect 28166 17184 28172 17196
rect 24360 17156 28172 17184
rect 24360 17144 24366 17156
rect 28166 17144 28172 17156
rect 28224 17144 28230 17196
rect 28353 17187 28411 17193
rect 28353 17153 28365 17187
rect 28399 17184 28411 17187
rect 28442 17184 28448 17196
rect 28399 17156 28448 17184
rect 28399 17153 28411 17156
rect 28353 17147 28411 17153
rect 28442 17144 28448 17156
rect 28500 17144 28506 17196
rect 28552 17193 28580 17292
rect 28718 17280 28724 17332
rect 28776 17280 28782 17332
rect 29914 17280 29920 17332
rect 29972 17320 29978 17332
rect 29972 17292 33456 17320
rect 29972 17280 29978 17292
rect 28629 17255 28687 17261
rect 28629 17221 28641 17255
rect 28675 17252 28687 17255
rect 28736 17252 28764 17280
rect 31220 17261 31248 17292
rect 33428 17261 33456 17292
rect 37458 17280 37464 17332
rect 37516 17320 37522 17332
rect 44266 17320 44272 17332
rect 37516 17292 44272 17320
rect 37516 17280 37522 17292
rect 31205 17255 31263 17261
rect 28675 17224 31064 17252
rect 28675 17221 28687 17224
rect 28629 17215 28687 17221
rect 31036 17196 31064 17224
rect 31205 17221 31217 17255
rect 31251 17221 31263 17255
rect 31205 17215 31263 17221
rect 31297 17255 31355 17261
rect 31297 17221 31309 17255
rect 31343 17252 31355 17255
rect 33413 17255 33471 17261
rect 31343 17224 31524 17252
rect 31343 17221 31355 17224
rect 31297 17215 31355 17221
rect 28537 17187 28595 17193
rect 28537 17153 28549 17187
rect 28583 17153 28595 17187
rect 28537 17147 28595 17153
rect 28721 17187 28779 17193
rect 28721 17153 28733 17187
rect 28767 17153 28779 17187
rect 31018 17184 31024 17196
rect 30979 17156 31024 17184
rect 28721 17147 28779 17153
rect 19426 17076 19432 17128
rect 19484 17116 19490 17128
rect 26326 17116 26332 17128
rect 19484 17088 26332 17116
rect 19484 17076 19490 17088
rect 26326 17076 26332 17088
rect 26384 17076 26390 17128
rect 28736 17116 28764 17147
rect 31018 17144 31024 17156
rect 31076 17144 31082 17196
rect 31389 17187 31447 17193
rect 31389 17153 31401 17187
rect 31435 17153 31447 17187
rect 31496 17184 31524 17224
rect 33413 17221 33425 17255
rect 33459 17252 33471 17255
rect 36446 17252 36452 17264
rect 33459 17224 36452 17252
rect 33459 17221 33471 17224
rect 33413 17215 33471 17221
rect 36446 17212 36452 17224
rect 36504 17212 36510 17264
rect 36538 17212 36544 17264
rect 36596 17252 36602 17264
rect 36596 17224 36641 17252
rect 36596 17212 36602 17224
rect 32398 17184 32404 17196
rect 31496 17156 32404 17184
rect 31389 17147 31447 17153
rect 27632 17088 28764 17116
rect 27632 17060 27660 17088
rect 31294 17076 31300 17128
rect 31352 17116 31358 17128
rect 31404 17116 31432 17147
rect 32398 17144 32404 17156
rect 32456 17184 32462 17196
rect 32493 17187 32551 17193
rect 32493 17184 32505 17187
rect 32456 17156 32505 17184
rect 32456 17144 32462 17156
rect 32493 17153 32505 17156
rect 32539 17184 32551 17187
rect 32950 17184 32956 17196
rect 32539 17156 32956 17184
rect 32539 17153 32551 17156
rect 32493 17147 32551 17153
rect 32950 17144 32956 17156
rect 33008 17184 33014 17196
rect 33229 17187 33287 17193
rect 33229 17184 33241 17187
rect 33008 17156 33241 17184
rect 33008 17144 33014 17156
rect 33229 17153 33241 17156
rect 33275 17153 33287 17187
rect 33502 17184 33508 17196
rect 33463 17156 33508 17184
rect 33229 17147 33287 17153
rect 33502 17144 33508 17156
rect 33560 17144 33566 17196
rect 33597 17187 33655 17193
rect 33597 17153 33609 17187
rect 33643 17153 33655 17187
rect 33597 17147 33655 17153
rect 33612 17116 33640 17147
rect 33686 17144 33692 17196
rect 33744 17184 33750 17196
rect 34333 17187 34391 17193
rect 34333 17184 34345 17187
rect 33744 17156 34345 17184
rect 33744 17144 33750 17156
rect 34333 17153 34345 17156
rect 34379 17184 34391 17187
rect 34422 17184 34428 17196
rect 34379 17156 34428 17184
rect 34379 17153 34391 17156
rect 34333 17147 34391 17153
rect 34422 17144 34428 17156
rect 34480 17184 34486 17196
rect 35989 17187 36047 17193
rect 35989 17184 36001 17187
rect 34480 17156 36001 17184
rect 34480 17144 34486 17156
rect 35989 17153 36001 17156
rect 36035 17184 36047 17187
rect 36556 17184 36584 17212
rect 36035 17156 36584 17184
rect 36035 17153 36047 17156
rect 35989 17147 36047 17153
rect 37366 17144 37372 17196
rect 37424 17184 37430 17196
rect 37461 17187 37519 17193
rect 37461 17184 37473 17187
rect 37424 17156 37473 17184
rect 37424 17144 37430 17156
rect 37461 17153 37473 17156
rect 37507 17153 37519 17187
rect 37660 17184 37688 17292
rect 44266 17280 44272 17292
rect 44324 17280 44330 17332
rect 45649 17323 45707 17329
rect 45649 17289 45661 17323
rect 45695 17320 45707 17323
rect 48314 17320 48320 17332
rect 45695 17292 48320 17320
rect 45695 17289 45707 17292
rect 45649 17283 45707 17289
rect 48314 17280 48320 17292
rect 48372 17280 48378 17332
rect 52917 17323 52975 17329
rect 52917 17289 52929 17323
rect 52963 17320 52975 17323
rect 53098 17320 53104 17332
rect 52963 17292 53104 17320
rect 52963 17289 52975 17292
rect 52917 17283 52975 17289
rect 53098 17280 53104 17292
rect 53156 17280 53162 17332
rect 58066 17320 58072 17332
rect 58027 17292 58072 17320
rect 58066 17280 58072 17292
rect 58124 17280 58130 17332
rect 37737 17255 37795 17261
rect 37737 17221 37749 17255
rect 37783 17252 37795 17255
rect 43898 17252 43904 17264
rect 37783 17224 43904 17252
rect 37783 17221 37795 17224
rect 37737 17215 37795 17221
rect 43898 17212 43904 17224
rect 43956 17212 43962 17264
rect 44082 17212 44088 17264
rect 44140 17252 44146 17264
rect 56318 17252 56324 17264
rect 44140 17224 56324 17252
rect 44140 17212 44146 17224
rect 56318 17212 56324 17224
rect 56376 17212 56382 17264
rect 56778 17212 56784 17264
rect 56836 17252 56842 17264
rect 57057 17255 57115 17261
rect 57057 17252 57069 17255
rect 56836 17224 57069 17252
rect 56836 17212 56842 17224
rect 57057 17221 57069 17224
rect 57103 17221 57115 17255
rect 57057 17215 57115 17221
rect 37829 17187 37887 17193
rect 37829 17184 37841 17187
rect 37660 17156 37841 17184
rect 37461 17147 37519 17153
rect 37829 17153 37841 17156
rect 37875 17153 37887 17187
rect 37829 17147 37887 17153
rect 40494 17144 40500 17196
rect 40552 17184 40558 17196
rect 40773 17187 40831 17193
rect 40773 17184 40785 17187
rect 40552 17156 40785 17184
rect 40552 17144 40558 17156
rect 40773 17153 40785 17156
rect 40819 17153 40831 17187
rect 40773 17147 40831 17153
rect 43990 17144 43996 17196
rect 44048 17184 44054 17196
rect 45281 17187 45339 17193
rect 45281 17184 45293 17187
rect 44048 17156 45293 17184
rect 44048 17144 44054 17156
rect 45281 17153 45293 17156
rect 45327 17153 45339 17187
rect 45281 17147 45339 17153
rect 45370 17144 45376 17196
rect 45428 17184 45434 17196
rect 48130 17184 48136 17196
rect 45428 17156 45473 17184
rect 48091 17156 48136 17184
rect 45428 17144 45434 17156
rect 48130 17144 48136 17156
rect 48188 17144 48194 17196
rect 49145 17187 49203 17193
rect 49145 17184 49157 17187
rect 48240 17156 49157 17184
rect 37277 17119 37335 17125
rect 37277 17116 37289 17119
rect 31352 17088 33640 17116
rect 36648 17088 37289 17116
rect 31352 17076 31358 17088
rect 21634 17048 21640 17060
rect 19352 17020 21640 17048
rect 18049 17011 18107 17017
rect 21634 17008 21640 17020
rect 21692 17008 21698 17060
rect 23290 17008 23296 17060
rect 23348 17048 23354 17060
rect 23569 17051 23627 17057
rect 23569 17048 23581 17051
rect 23348 17020 23581 17048
rect 23348 17008 23354 17020
rect 23569 17017 23581 17020
rect 23615 17017 23627 17051
rect 23569 17011 23627 17017
rect 26145 17051 26203 17057
rect 26145 17017 26157 17051
rect 26191 17048 26203 17051
rect 27614 17048 27620 17060
rect 26191 17020 27620 17048
rect 26191 17017 26203 17020
rect 26145 17011 26203 17017
rect 27614 17008 27620 17020
rect 27672 17008 27678 17060
rect 30834 17008 30840 17060
rect 30892 17048 30898 17060
rect 35342 17048 35348 17060
rect 30892 17020 35348 17048
rect 30892 17008 30898 17020
rect 35342 17008 35348 17020
rect 35400 17008 35406 17060
rect 10134 16980 10140 16992
rect 9646 16952 10140 16980
rect 10134 16940 10140 16952
rect 10192 16940 10198 16992
rect 14645 16983 14703 16989
rect 14645 16949 14657 16983
rect 14691 16980 14703 16983
rect 15010 16980 15016 16992
rect 14691 16952 15016 16980
rect 14691 16949 14703 16952
rect 14645 16943 14703 16949
rect 15010 16940 15016 16952
rect 15068 16940 15074 16992
rect 15470 16940 15476 16992
rect 15528 16980 15534 16992
rect 15657 16983 15715 16989
rect 15657 16980 15669 16983
rect 15528 16952 15669 16980
rect 15528 16940 15534 16952
rect 15657 16949 15669 16952
rect 15703 16949 15715 16983
rect 15657 16943 15715 16949
rect 16298 16940 16304 16992
rect 16356 16980 16362 16992
rect 20070 16980 20076 16992
rect 16356 16952 20076 16980
rect 16356 16940 16362 16952
rect 20070 16940 20076 16952
rect 20128 16940 20134 16992
rect 20162 16940 20168 16992
rect 20220 16980 20226 16992
rect 20533 16983 20591 16989
rect 20533 16980 20545 16983
rect 20220 16952 20545 16980
rect 20220 16940 20226 16952
rect 20533 16949 20545 16952
rect 20579 16949 20591 16983
rect 20533 16943 20591 16949
rect 24581 16983 24639 16989
rect 24581 16949 24593 16983
rect 24627 16980 24639 16983
rect 25222 16980 25228 16992
rect 24627 16952 25228 16980
rect 24627 16949 24639 16952
rect 24581 16943 24639 16949
rect 25222 16940 25228 16952
rect 25280 16980 25286 16992
rect 26786 16980 26792 16992
rect 25280 16952 26792 16980
rect 25280 16940 25286 16952
rect 26786 16940 26792 16952
rect 26844 16940 26850 16992
rect 28905 16983 28963 16989
rect 28905 16949 28917 16983
rect 28951 16980 28963 16983
rect 29178 16980 29184 16992
rect 28951 16952 29184 16980
rect 28951 16949 28963 16952
rect 28905 16943 28963 16949
rect 29178 16940 29184 16952
rect 29236 16940 29242 16992
rect 29822 16940 29828 16992
rect 29880 16980 29886 16992
rect 30006 16980 30012 16992
rect 29880 16952 30012 16980
rect 29880 16940 29886 16952
rect 30006 16940 30012 16952
rect 30064 16940 30070 16992
rect 31386 16940 31392 16992
rect 31444 16980 31450 16992
rect 31573 16983 31631 16989
rect 31573 16980 31585 16983
rect 31444 16952 31585 16980
rect 31444 16940 31450 16952
rect 31573 16949 31585 16952
rect 31619 16949 31631 16983
rect 32674 16980 32680 16992
rect 32635 16952 32680 16980
rect 31573 16943 31631 16949
rect 32674 16940 32680 16952
rect 32732 16940 32738 16992
rect 33778 16980 33784 16992
rect 33739 16952 33784 16980
rect 33778 16940 33784 16952
rect 33836 16940 33842 16992
rect 36354 16940 36360 16992
rect 36412 16980 36418 16992
rect 36648 16989 36676 17088
rect 37277 17085 37289 17088
rect 37323 17085 37335 17119
rect 40681 17119 40739 17125
rect 40681 17116 40693 17119
rect 37277 17079 37335 17085
rect 40052 17088 40693 17116
rect 40052 16992 40080 17088
rect 40681 17085 40693 17088
rect 40727 17085 40739 17119
rect 40681 17079 40739 17085
rect 48041 17119 48099 17125
rect 48041 17085 48053 17119
rect 48087 17116 48099 17119
rect 48240 17116 48268 17156
rect 49145 17153 49157 17156
rect 49191 17153 49203 17187
rect 49145 17147 49203 17153
rect 49329 17187 49387 17193
rect 49329 17153 49341 17187
rect 49375 17184 49387 17187
rect 50433 17187 50491 17193
rect 50433 17184 50445 17187
rect 49375 17156 50445 17184
rect 49375 17153 49387 17156
rect 49329 17147 49387 17153
rect 48498 17116 48504 17128
rect 48087 17088 48268 17116
rect 48459 17088 48504 17116
rect 48087 17085 48099 17088
rect 48041 17079 48099 17085
rect 41141 17051 41199 17057
rect 41141 17017 41153 17051
rect 41187 17048 41199 17051
rect 48056 17048 48084 17079
rect 48498 17076 48504 17088
rect 48556 17076 48562 17128
rect 48961 17119 49019 17125
rect 48961 17085 48973 17119
rect 49007 17085 49019 17119
rect 48961 17079 49019 17085
rect 41187 17020 48084 17048
rect 41187 17017 41199 17020
rect 41141 17011 41199 17017
rect 48130 17008 48136 17060
rect 48188 17048 48194 17060
rect 48976 17048 49004 17079
rect 48188 17020 49004 17048
rect 50080 17048 50108 17156
rect 50433 17153 50445 17156
rect 50479 17153 50491 17187
rect 50798 17184 50804 17196
rect 50759 17156 50804 17184
rect 50433 17147 50491 17153
rect 50798 17144 50804 17156
rect 50856 17184 50862 17196
rect 51261 17187 51319 17193
rect 51261 17184 51273 17187
rect 50856 17156 51273 17184
rect 50856 17144 50862 17156
rect 51261 17153 51273 17156
rect 51307 17153 51319 17187
rect 51261 17147 51319 17153
rect 52546 17144 52552 17196
rect 52604 17184 52610 17196
rect 52733 17187 52791 17193
rect 52733 17184 52745 17187
rect 52604 17156 52745 17184
rect 52604 17144 52610 17156
rect 52733 17153 52745 17156
rect 52779 17153 52791 17187
rect 52733 17147 52791 17153
rect 53009 17187 53067 17193
rect 53009 17153 53021 17187
rect 53055 17184 53067 17187
rect 53190 17184 53196 17196
rect 53055 17156 53196 17184
rect 53055 17153 53067 17156
rect 53009 17147 53067 17153
rect 53190 17144 53196 17156
rect 53248 17144 53254 17196
rect 53650 17184 53656 17196
rect 53611 17156 53656 17184
rect 53650 17144 53656 17156
rect 53708 17144 53714 17196
rect 53742 17144 53748 17196
rect 53800 17184 53806 17196
rect 54021 17187 54079 17193
rect 54021 17184 54033 17187
rect 53800 17156 54033 17184
rect 53800 17144 53806 17156
rect 54021 17153 54033 17156
rect 54067 17153 54079 17187
rect 57146 17184 57152 17196
rect 56994 17156 57152 17184
rect 54021 17147 54079 17153
rect 57146 17144 57152 17156
rect 57204 17144 57210 17196
rect 50246 17116 50252 17128
rect 50207 17088 50252 17116
rect 50246 17076 50252 17088
rect 50304 17116 50310 17128
rect 51353 17119 51411 17125
rect 51353 17116 51365 17119
rect 50304 17088 51365 17116
rect 50304 17076 50310 17088
rect 51353 17085 51365 17088
rect 51399 17085 51411 17119
rect 53466 17116 53472 17128
rect 53427 17088 53472 17116
rect 51353 17079 51411 17085
rect 53466 17076 53472 17088
rect 53524 17076 53530 17128
rect 56134 17076 56140 17128
rect 56192 17116 56198 17128
rect 56505 17119 56563 17125
rect 56505 17116 56517 17119
rect 56192 17088 56517 17116
rect 56192 17076 56198 17088
rect 56505 17085 56517 17088
rect 56551 17085 56563 17119
rect 56505 17079 56563 17085
rect 52730 17048 52736 17060
rect 50080 17020 51304 17048
rect 52691 17020 52736 17048
rect 48188 17008 48194 17020
rect 36633 16983 36691 16989
rect 36633 16980 36645 16983
rect 36412 16952 36645 16980
rect 36412 16940 36418 16952
rect 36633 16949 36645 16952
rect 36679 16949 36691 16983
rect 40034 16980 40040 16992
rect 39995 16952 40040 16980
rect 36633 16943 36691 16949
rect 40034 16940 40040 16952
rect 40092 16940 40098 16992
rect 44174 16940 44180 16992
rect 44232 16980 44238 16992
rect 45278 16980 45284 16992
rect 44232 16952 45284 16980
rect 44232 16940 44238 16952
rect 45278 16940 45284 16952
rect 45336 16940 45342 16992
rect 50709 16983 50767 16989
rect 50709 16949 50721 16983
rect 50755 16980 50767 16983
rect 51166 16980 51172 16992
rect 50755 16952 51172 16980
rect 50755 16949 50767 16952
rect 50709 16943 50767 16949
rect 51166 16940 51172 16952
rect 51224 16940 51230 16992
rect 51276 16989 51304 17020
rect 52730 17008 52736 17020
rect 52788 17008 52794 17060
rect 53929 17051 53987 17057
rect 53929 17017 53941 17051
rect 53975 17048 53987 17051
rect 56318 17048 56324 17060
rect 53975 17020 56324 17048
rect 53975 17017 53987 17020
rect 53929 17011 53987 17017
rect 56318 17008 56324 17020
rect 56376 17008 56382 17060
rect 51261 16983 51319 16989
rect 51261 16949 51273 16983
rect 51307 16949 51319 16983
rect 51626 16980 51632 16992
rect 51587 16952 51632 16980
rect 51261 16943 51319 16949
rect 51626 16940 51632 16952
rect 51684 16940 51690 16992
rect 51810 16940 51816 16992
rect 51868 16980 51874 16992
rect 56134 16980 56140 16992
rect 51868 16952 56140 16980
rect 51868 16940 51874 16952
rect 56134 16940 56140 16952
rect 56192 16940 56198 16992
rect 1104 16890 58880 16912
rect 1104 16838 4214 16890
rect 4266 16838 4278 16890
rect 4330 16838 4342 16890
rect 4394 16838 4406 16890
rect 4458 16838 4470 16890
rect 4522 16838 34934 16890
rect 34986 16838 34998 16890
rect 35050 16838 35062 16890
rect 35114 16838 35126 16890
rect 35178 16838 35190 16890
rect 35242 16838 58880 16890
rect 1104 16816 58880 16838
rect 1949 16779 2007 16785
rect 1949 16745 1961 16779
rect 1995 16776 2007 16779
rect 3326 16776 3332 16788
rect 1995 16748 3332 16776
rect 1995 16745 2007 16748
rect 1949 16739 2007 16745
rect 3326 16736 3332 16748
rect 3384 16736 3390 16788
rect 7006 16736 7012 16788
rect 7064 16776 7070 16788
rect 7834 16776 7840 16788
rect 7064 16748 7840 16776
rect 7064 16736 7070 16748
rect 7834 16736 7840 16748
rect 7892 16776 7898 16788
rect 9030 16776 9036 16788
rect 7892 16748 9036 16776
rect 7892 16736 7898 16748
rect 9030 16736 9036 16748
rect 9088 16736 9094 16788
rect 10042 16736 10048 16788
rect 10100 16776 10106 16788
rect 10413 16779 10471 16785
rect 10413 16776 10425 16779
rect 10100 16748 10425 16776
rect 10100 16736 10106 16748
rect 10413 16745 10425 16748
rect 10459 16745 10471 16779
rect 12894 16776 12900 16788
rect 12855 16748 12900 16776
rect 10413 16739 10471 16745
rect 12894 16736 12900 16748
rect 12952 16736 12958 16788
rect 13449 16779 13507 16785
rect 13449 16745 13461 16779
rect 13495 16776 13507 16779
rect 14458 16776 14464 16788
rect 13495 16748 14464 16776
rect 13495 16745 13507 16748
rect 13449 16739 13507 16745
rect 14458 16736 14464 16748
rect 14516 16736 14522 16788
rect 15565 16779 15623 16785
rect 15565 16745 15577 16779
rect 15611 16776 15623 16779
rect 33042 16776 33048 16788
rect 15611 16748 33048 16776
rect 15611 16745 15623 16748
rect 15565 16739 15623 16745
rect 33042 16736 33048 16748
rect 33100 16736 33106 16788
rect 45922 16776 45928 16788
rect 38488 16748 45928 16776
rect 2866 16708 2872 16720
rect 2827 16680 2872 16708
rect 2866 16668 2872 16680
rect 2924 16668 2930 16720
rect 5813 16711 5871 16717
rect 5813 16677 5825 16711
rect 5859 16708 5871 16711
rect 9122 16708 9128 16720
rect 5859 16680 9128 16708
rect 5859 16677 5871 16680
rect 5813 16671 5871 16677
rect 9122 16668 9128 16680
rect 9180 16668 9186 16720
rect 9493 16711 9551 16717
rect 9493 16677 9505 16711
rect 9539 16708 9551 16711
rect 9950 16708 9956 16720
rect 9539 16680 9956 16708
rect 9539 16677 9551 16680
rect 9493 16671 9551 16677
rect 9950 16668 9956 16680
rect 10008 16668 10014 16720
rect 11882 16668 11888 16720
rect 11940 16708 11946 16720
rect 11977 16711 12035 16717
rect 11977 16708 11989 16711
rect 11940 16680 11989 16708
rect 11940 16668 11946 16680
rect 11977 16677 11989 16680
rect 12023 16708 12035 16711
rect 12805 16711 12863 16717
rect 12805 16708 12817 16711
rect 12023 16680 12817 16708
rect 12023 16677 12035 16680
rect 11977 16671 12035 16677
rect 12805 16677 12817 16680
rect 12851 16708 12863 16711
rect 13538 16708 13544 16720
rect 12851 16680 13544 16708
rect 12851 16677 12863 16680
rect 12805 16671 12863 16677
rect 13538 16668 13544 16680
rect 13596 16668 13602 16720
rect 14090 16668 14096 16720
rect 14148 16708 14154 16720
rect 14148 16680 14964 16708
rect 14148 16668 14154 16680
rect 3237 16643 3295 16649
rect 3237 16609 3249 16643
rect 3283 16640 3295 16643
rect 3418 16640 3424 16652
rect 3283 16612 3424 16640
rect 3283 16609 3295 16612
rect 3237 16603 3295 16609
rect 3418 16600 3424 16612
rect 3476 16600 3482 16652
rect 4154 16572 4160 16584
rect 4115 16544 4160 16572
rect 4154 16532 4160 16544
rect 4212 16532 4218 16584
rect 4614 16572 4620 16584
rect 4575 16544 4620 16572
rect 4614 16532 4620 16544
rect 4672 16532 4678 16584
rect 7466 16532 7472 16584
rect 7524 16572 7530 16584
rect 7745 16575 7803 16581
rect 7745 16572 7757 16575
rect 7524 16544 7757 16572
rect 7524 16532 7530 16544
rect 7745 16541 7757 16544
rect 7791 16541 7803 16575
rect 7745 16535 7803 16541
rect 7929 16575 7987 16581
rect 7929 16541 7941 16575
rect 7975 16541 7987 16575
rect 7929 16535 7987 16541
rect 1854 16504 1860 16516
rect 1815 16476 1860 16504
rect 1854 16464 1860 16476
rect 1912 16464 1918 16516
rect 7285 16507 7343 16513
rect 7285 16473 7297 16507
rect 7331 16504 7343 16507
rect 7944 16504 7972 16535
rect 8478 16532 8484 16584
rect 8536 16572 8542 16584
rect 9030 16572 9036 16584
rect 8536 16544 9036 16572
rect 8536 16532 8542 16544
rect 9030 16532 9036 16544
rect 9088 16572 9094 16584
rect 9401 16575 9459 16581
rect 9401 16572 9413 16575
rect 9088 16544 9413 16572
rect 9088 16532 9094 16544
rect 9401 16541 9413 16544
rect 9447 16541 9459 16575
rect 9401 16535 9459 16541
rect 9493 16575 9551 16581
rect 9493 16541 9505 16575
rect 9539 16541 9551 16575
rect 9493 16535 9551 16541
rect 8202 16504 8208 16516
rect 7331 16476 8208 16504
rect 7331 16473 7343 16476
rect 7285 16467 7343 16473
rect 8202 16464 8208 16476
rect 8260 16464 8266 16516
rect 9214 16504 9220 16516
rect 9175 16476 9220 16504
rect 9214 16464 9220 16476
rect 9272 16464 9278 16516
rect 9306 16464 9312 16516
rect 9364 16504 9370 16516
rect 9508 16504 9536 16535
rect 9674 16532 9680 16584
rect 9732 16572 9738 16584
rect 14185 16575 14243 16581
rect 9732 16544 13860 16572
rect 9732 16532 9738 16544
rect 9364 16476 9536 16504
rect 9364 16464 9370 16476
rect 10134 16464 10140 16516
rect 10192 16504 10198 16516
rect 10229 16507 10287 16513
rect 10229 16504 10241 16507
rect 10192 16476 10241 16504
rect 10192 16464 10198 16476
rect 10229 16473 10241 16476
rect 10275 16473 10287 16507
rect 10410 16504 10416 16516
rect 10371 16476 10416 16504
rect 10229 16467 10287 16473
rect 10410 16464 10416 16476
rect 10468 16464 10474 16516
rect 12434 16464 12440 16516
rect 12492 16504 12498 16516
rect 13832 16504 13860 16544
rect 14185 16541 14197 16575
rect 14231 16572 14243 16575
rect 14292 16572 14320 16680
rect 14826 16640 14832 16652
rect 14231 16544 14320 16572
rect 14384 16612 14832 16640
rect 14231 16541 14243 16544
rect 14185 16535 14243 16541
rect 14384 16513 14412 16612
rect 14826 16600 14832 16612
rect 14884 16600 14890 16652
rect 14936 16640 14964 16680
rect 15286 16668 15292 16720
rect 15344 16708 15350 16720
rect 15344 16680 19472 16708
rect 15344 16668 15350 16680
rect 14936 16612 15608 16640
rect 14550 16572 14556 16584
rect 14511 16544 14556 16572
rect 14550 16532 14556 16544
rect 14608 16532 14614 16584
rect 15470 16572 15476 16584
rect 15431 16544 15476 16572
rect 15470 16532 15476 16544
rect 15528 16532 15534 16584
rect 15580 16572 15608 16612
rect 16114 16600 16120 16652
rect 16172 16640 16178 16652
rect 16853 16643 16911 16649
rect 16853 16640 16865 16643
rect 16172 16612 16865 16640
rect 16172 16600 16178 16612
rect 16853 16609 16865 16612
rect 16899 16609 16911 16643
rect 19444 16640 19472 16680
rect 19518 16668 19524 16720
rect 19576 16708 19582 16720
rect 20717 16711 20775 16717
rect 20717 16708 20729 16711
rect 19576 16680 20024 16708
rect 19576 16668 19582 16680
rect 19702 16640 19708 16652
rect 19444 16612 19564 16640
rect 19663 16612 19708 16640
rect 16853 16603 16911 16609
rect 16666 16572 16672 16584
rect 15580 16544 16672 16572
rect 16666 16532 16672 16544
rect 16724 16532 16730 16584
rect 19536 16572 19564 16612
rect 19702 16600 19708 16612
rect 19760 16600 19766 16652
rect 19794 16572 19800 16584
rect 19536 16544 19800 16572
rect 19794 16532 19800 16544
rect 19852 16532 19858 16584
rect 19996 16581 20024 16680
rect 20272 16680 20729 16708
rect 19889 16575 19947 16581
rect 19889 16541 19901 16575
rect 19935 16541 19947 16575
rect 19889 16535 19947 16541
rect 19981 16575 20039 16581
rect 19981 16541 19993 16575
rect 20027 16541 20039 16575
rect 20162 16572 20168 16584
rect 20123 16544 20168 16572
rect 19981 16535 20039 16541
rect 14369 16507 14427 16513
rect 14369 16504 14381 16507
rect 12492 16476 12537 16504
rect 13832 16476 14381 16504
rect 12492 16464 12498 16476
rect 14369 16473 14381 16476
rect 14415 16473 14427 16507
rect 14369 16467 14427 16473
rect 14458 16464 14464 16516
rect 14516 16504 14522 16516
rect 15289 16507 15347 16513
rect 14516 16476 14561 16504
rect 14516 16464 14522 16476
rect 15289 16473 15301 16507
rect 15335 16473 15347 16507
rect 19904 16504 19932 16535
rect 20162 16532 20168 16544
rect 20220 16532 20226 16584
rect 20272 16581 20300 16680
rect 20717 16677 20729 16680
rect 20763 16677 20775 16711
rect 20717 16671 20775 16677
rect 23845 16711 23903 16717
rect 23845 16677 23857 16711
rect 23891 16677 23903 16711
rect 23845 16671 23903 16677
rect 24857 16711 24915 16717
rect 24857 16677 24869 16711
rect 24903 16708 24915 16711
rect 27065 16711 27123 16717
rect 24903 16680 27016 16708
rect 24903 16677 24915 16680
rect 24857 16671 24915 16677
rect 23860 16640 23888 16671
rect 26988 16640 27016 16680
rect 27065 16677 27077 16711
rect 27111 16708 27123 16711
rect 27111 16680 36216 16708
rect 27111 16677 27123 16680
rect 27065 16671 27123 16677
rect 27706 16640 27712 16652
rect 23860 16612 23980 16640
rect 26988 16612 27712 16640
rect 20257 16575 20315 16581
rect 20257 16541 20269 16575
rect 20303 16541 20315 16575
rect 20257 16535 20315 16541
rect 20346 16532 20352 16584
rect 20404 16572 20410 16584
rect 20901 16575 20959 16581
rect 20901 16572 20913 16575
rect 20404 16544 20913 16572
rect 20404 16532 20410 16544
rect 20901 16541 20913 16544
rect 20947 16541 20959 16575
rect 21266 16572 21272 16584
rect 21227 16544 21272 16572
rect 20901 16535 20959 16541
rect 21266 16532 21272 16544
rect 21324 16532 21330 16584
rect 23290 16532 23296 16584
rect 23348 16572 23354 16584
rect 23569 16575 23627 16581
rect 23569 16572 23581 16575
rect 23348 16544 23581 16572
rect 23348 16532 23354 16544
rect 23569 16541 23581 16544
rect 23615 16541 23627 16575
rect 23842 16572 23848 16584
rect 23803 16544 23848 16572
rect 23569 16535 23627 16541
rect 23842 16532 23848 16544
rect 23900 16532 23906 16584
rect 20438 16504 20444 16516
rect 19904 16476 20444 16504
rect 15289 16467 15347 16473
rect 2774 16396 2780 16448
rect 2832 16436 2838 16448
rect 10594 16436 10600 16448
rect 2832 16408 2877 16436
rect 10555 16408 10600 16436
rect 2832 16396 2838 16408
rect 10594 16396 10600 16408
rect 10652 16396 10658 16448
rect 14737 16439 14795 16445
rect 14737 16405 14749 16439
rect 14783 16436 14795 16439
rect 15304 16436 15332 16467
rect 20438 16464 20444 16476
rect 20496 16464 20502 16516
rect 20714 16464 20720 16516
rect 20772 16504 20778 16516
rect 20993 16507 21051 16513
rect 20993 16504 21005 16507
rect 20772 16476 21005 16504
rect 20772 16464 20778 16476
rect 20993 16473 21005 16476
rect 21039 16473 21051 16507
rect 20993 16467 21051 16473
rect 21085 16507 21143 16513
rect 21085 16473 21097 16507
rect 21131 16473 21143 16507
rect 23952 16504 23980 16612
rect 27706 16600 27712 16612
rect 27764 16600 27770 16652
rect 28350 16600 28356 16652
rect 28408 16640 28414 16652
rect 30834 16640 30840 16652
rect 28408 16612 28453 16640
rect 30795 16612 30840 16640
rect 28408 16600 28414 16612
rect 30834 16600 30840 16612
rect 30892 16600 30898 16652
rect 31386 16640 31392 16652
rect 31347 16612 31392 16640
rect 31386 16600 31392 16612
rect 31444 16600 31450 16652
rect 32490 16600 32496 16652
rect 32548 16640 32554 16652
rect 33229 16643 33287 16649
rect 33229 16640 33241 16643
rect 32548 16612 33241 16640
rect 32548 16600 32554 16612
rect 33229 16609 33241 16612
rect 33275 16609 33287 16643
rect 33229 16603 33287 16609
rect 33778 16600 33784 16652
rect 33836 16640 33842 16652
rect 34701 16643 34759 16649
rect 34701 16640 34713 16643
rect 33836 16612 34713 16640
rect 33836 16600 33842 16612
rect 34701 16609 34713 16612
rect 34747 16609 34759 16643
rect 35250 16640 35256 16652
rect 35211 16612 35256 16640
rect 34701 16603 34759 16609
rect 35250 16600 35256 16612
rect 35308 16600 35314 16652
rect 36188 16649 36216 16680
rect 36173 16643 36231 16649
rect 36173 16609 36185 16643
rect 36219 16609 36231 16643
rect 36173 16603 36231 16609
rect 37093 16643 37151 16649
rect 37093 16609 37105 16643
rect 37139 16640 37151 16643
rect 38488 16640 38516 16748
rect 45922 16736 45928 16748
rect 45980 16736 45986 16788
rect 46293 16779 46351 16785
rect 46293 16745 46305 16779
rect 46339 16776 46351 16779
rect 48130 16776 48136 16788
rect 46339 16748 48136 16776
rect 46339 16745 46351 16748
rect 46293 16739 46351 16745
rect 48130 16736 48136 16748
rect 48188 16736 48194 16788
rect 50154 16776 50160 16788
rect 50115 16748 50160 16776
rect 50154 16736 50160 16748
rect 50212 16776 50218 16788
rect 50798 16776 50804 16788
rect 50212 16748 50804 16776
rect 50212 16736 50218 16748
rect 50798 16736 50804 16748
rect 50856 16776 50862 16788
rect 51077 16779 51135 16785
rect 51077 16776 51089 16779
rect 50856 16748 51089 16776
rect 50856 16736 50862 16748
rect 51077 16745 51089 16748
rect 51123 16745 51135 16779
rect 51077 16739 51135 16745
rect 52181 16779 52239 16785
rect 52181 16745 52193 16779
rect 52227 16776 52239 16779
rect 53466 16776 53472 16788
rect 52227 16748 53472 16776
rect 52227 16745 52239 16748
rect 52181 16739 52239 16745
rect 53466 16736 53472 16748
rect 53524 16736 53530 16788
rect 53650 16776 53656 16788
rect 53611 16748 53656 16776
rect 53650 16736 53656 16748
rect 53708 16736 53714 16788
rect 53742 16736 53748 16788
rect 53800 16776 53806 16788
rect 54113 16779 54171 16785
rect 54113 16776 54125 16779
rect 53800 16748 54125 16776
rect 53800 16736 53806 16748
rect 54113 16745 54125 16748
rect 54159 16745 54171 16779
rect 54113 16739 54171 16745
rect 54297 16779 54355 16785
rect 54297 16745 54309 16779
rect 54343 16745 54355 16779
rect 54297 16739 54355 16745
rect 39025 16711 39083 16717
rect 39025 16677 39037 16711
rect 39071 16708 39083 16711
rect 43990 16708 43996 16720
rect 39071 16680 41414 16708
rect 43951 16680 43996 16708
rect 39071 16677 39083 16680
rect 39025 16671 39083 16677
rect 38746 16640 38752 16652
rect 37139 16612 38516 16640
rect 38707 16612 38752 16640
rect 37139 16609 37151 16612
rect 37093 16603 37151 16609
rect 38746 16600 38752 16612
rect 38804 16600 38810 16652
rect 41386 16640 41414 16680
rect 43990 16668 43996 16680
rect 44048 16668 44054 16720
rect 47121 16711 47179 16717
rect 46032 16680 46980 16708
rect 46032 16649 46060 16680
rect 46017 16643 46075 16649
rect 46017 16640 46029 16643
rect 41386 16612 46029 16640
rect 46017 16609 46029 16612
rect 46063 16609 46075 16643
rect 46017 16603 46075 16609
rect 24118 16532 24124 16584
rect 24176 16572 24182 16584
rect 24397 16575 24455 16581
rect 24397 16572 24409 16575
rect 24176 16544 24409 16572
rect 24176 16532 24182 16544
rect 24397 16541 24409 16544
rect 24443 16541 24455 16575
rect 24397 16535 24455 16541
rect 24486 16532 24492 16584
rect 24544 16572 24550 16584
rect 24673 16575 24731 16581
rect 24544 16544 24589 16572
rect 24544 16532 24550 16544
rect 24673 16541 24685 16575
rect 24719 16541 24731 16575
rect 26418 16572 26424 16584
rect 26379 16544 26424 16572
rect 24673 16535 24731 16541
rect 24688 16504 24716 16535
rect 26418 16532 26424 16544
rect 26476 16532 26482 16584
rect 26510 16532 26516 16584
rect 26568 16572 26574 16584
rect 26786 16572 26792 16584
rect 26568 16544 26613 16572
rect 26747 16544 26792 16572
rect 26568 16532 26574 16544
rect 26786 16532 26792 16544
rect 26844 16532 26850 16584
rect 26927 16575 26985 16581
rect 26927 16541 26939 16575
rect 26973 16572 26985 16575
rect 28074 16572 28080 16584
rect 26973 16544 27936 16572
rect 28035 16544 28080 16572
rect 26973 16541 26985 16544
rect 26927 16535 26985 16541
rect 26697 16507 26755 16513
rect 26697 16504 26709 16507
rect 23952 16476 24716 16504
rect 25884 16476 26709 16504
rect 21085 16467 21143 16473
rect 14783 16408 15332 16436
rect 14783 16405 14795 16408
rect 14737 16399 14795 16405
rect 15838 16396 15844 16448
rect 15896 16436 15902 16448
rect 16298 16436 16304 16448
rect 15896 16408 16304 16436
rect 15896 16396 15902 16408
rect 16298 16396 16304 16408
rect 16356 16396 16362 16448
rect 20070 16396 20076 16448
rect 20128 16436 20134 16448
rect 21100 16436 21128 16467
rect 20128 16408 21128 16436
rect 20128 16396 20134 16408
rect 23382 16396 23388 16448
rect 23440 16436 23446 16448
rect 23661 16439 23719 16445
rect 23661 16436 23673 16439
rect 23440 16408 23673 16436
rect 23440 16396 23446 16408
rect 23661 16405 23673 16408
rect 23707 16405 23719 16439
rect 23661 16399 23719 16405
rect 25130 16396 25136 16448
rect 25188 16436 25194 16448
rect 25884 16445 25912 16476
rect 26697 16473 26709 16476
rect 26743 16473 26755 16507
rect 27908 16504 27936 16544
rect 28074 16532 28080 16544
rect 28132 16532 28138 16584
rect 28626 16532 28632 16584
rect 28684 16572 28690 16584
rect 31021 16575 31079 16581
rect 31021 16572 31033 16575
rect 28684 16544 31033 16572
rect 28684 16532 28690 16544
rect 31021 16541 31033 16544
rect 31067 16541 31079 16575
rect 32950 16572 32956 16584
rect 32911 16544 32956 16572
rect 31021 16535 31079 16541
rect 32950 16532 32956 16544
rect 33008 16532 33014 16584
rect 33962 16532 33968 16584
rect 34020 16572 34026 16584
rect 35069 16575 35127 16581
rect 35069 16572 35081 16575
rect 34020 16544 35081 16572
rect 34020 16532 34026 16544
rect 35069 16541 35081 16544
rect 35115 16541 35127 16575
rect 35069 16535 35127 16541
rect 36078 16532 36084 16584
rect 36136 16572 36142 16584
rect 36265 16575 36323 16581
rect 36265 16572 36277 16575
rect 36136 16544 36277 16572
rect 36136 16532 36142 16544
rect 36265 16541 36277 16544
rect 36311 16541 36323 16575
rect 36265 16535 36323 16541
rect 37182 16532 37188 16584
rect 37240 16572 37246 16584
rect 38654 16572 38660 16584
rect 37240 16544 38660 16572
rect 37240 16532 37246 16544
rect 38654 16532 38660 16544
rect 38712 16532 38718 16584
rect 43165 16575 43223 16581
rect 43165 16541 43177 16575
rect 43211 16572 43223 16575
rect 43254 16572 43260 16584
rect 43211 16544 43260 16572
rect 43211 16541 43223 16544
rect 43165 16535 43223 16541
rect 43254 16532 43260 16544
rect 43312 16532 43318 16584
rect 43717 16575 43775 16581
rect 43717 16541 43729 16575
rect 43763 16541 43775 16575
rect 43717 16535 43775 16541
rect 28442 16504 28448 16516
rect 27908 16476 28448 16504
rect 26697 16467 26755 16473
rect 28442 16464 28448 16476
rect 28500 16464 28506 16516
rect 31297 16507 31355 16513
rect 28552 16476 29960 16504
rect 25869 16439 25927 16445
rect 25869 16436 25881 16439
rect 25188 16408 25881 16436
rect 25188 16396 25194 16408
rect 25869 16405 25881 16408
rect 25915 16405 25927 16439
rect 25869 16399 25927 16405
rect 26878 16396 26884 16448
rect 26936 16436 26942 16448
rect 28552 16436 28580 16476
rect 26936 16408 28580 16436
rect 29733 16439 29791 16445
rect 26936 16396 26942 16408
rect 29733 16405 29745 16439
rect 29779 16436 29791 16439
rect 29822 16436 29828 16448
rect 29779 16408 29828 16436
rect 29779 16405 29791 16408
rect 29733 16399 29791 16405
rect 29822 16396 29828 16408
rect 29880 16396 29886 16448
rect 29932 16436 29960 16476
rect 31297 16473 31309 16507
rect 31343 16504 31355 16507
rect 42518 16504 42524 16516
rect 31343 16476 42524 16504
rect 31343 16473 31355 16476
rect 31297 16467 31355 16473
rect 42518 16464 42524 16476
rect 42576 16504 42582 16516
rect 42889 16507 42947 16513
rect 42889 16504 42901 16507
rect 42576 16476 42901 16504
rect 42576 16464 42582 16476
rect 42889 16473 42901 16476
rect 42935 16473 42947 16507
rect 42889 16467 42947 16473
rect 43073 16507 43131 16513
rect 43073 16473 43085 16507
rect 43119 16473 43131 16507
rect 43732 16504 43760 16535
rect 43898 16532 43904 16584
rect 43956 16572 43962 16584
rect 43993 16575 44051 16581
rect 43993 16572 44005 16575
rect 43956 16544 44005 16572
rect 43956 16532 43962 16544
rect 43993 16541 44005 16544
rect 44039 16541 44051 16575
rect 45922 16572 45928 16584
rect 45835 16544 45928 16572
rect 43993 16535 44051 16541
rect 45922 16532 45928 16544
rect 45980 16572 45986 16584
rect 46952 16581 46980 16680
rect 47121 16677 47133 16711
rect 47167 16708 47179 16711
rect 50246 16708 50252 16720
rect 47167 16680 50252 16708
rect 47167 16677 47179 16680
rect 47121 16671 47179 16677
rect 50246 16668 50252 16680
rect 50304 16668 50310 16720
rect 53098 16668 53104 16720
rect 53156 16708 53162 16720
rect 54312 16708 54340 16739
rect 53156 16680 54340 16708
rect 53156 16668 53162 16680
rect 51166 16600 51172 16652
rect 51224 16640 51230 16652
rect 51224 16612 51580 16640
rect 51224 16600 51230 16612
rect 46753 16575 46811 16581
rect 46753 16572 46765 16575
rect 45980 16544 46765 16572
rect 45980 16532 45986 16544
rect 46753 16541 46765 16544
rect 46799 16541 46811 16575
rect 46753 16535 46811 16541
rect 46937 16575 46995 16581
rect 46937 16541 46949 16575
rect 46983 16541 46995 16575
rect 51552 16572 51580 16612
rect 51626 16600 51632 16652
rect 51684 16640 51690 16652
rect 51684 16612 52040 16640
rect 51684 16600 51690 16612
rect 51810 16572 51816 16584
rect 51552 16544 51816 16572
rect 46937 16535 46995 16541
rect 51810 16532 51816 16544
rect 51868 16532 51874 16584
rect 52012 16581 52040 16612
rect 52546 16600 52552 16652
rect 52604 16640 52610 16652
rect 57146 16640 57152 16652
rect 52604 16612 53512 16640
rect 57107 16612 57152 16640
rect 52604 16600 52610 16612
rect 51997 16575 52055 16581
rect 51997 16541 52009 16575
rect 52043 16574 52055 16575
rect 52043 16546 52077 16574
rect 53190 16572 53196 16584
rect 52043 16541 52055 16546
rect 53103 16544 53196 16572
rect 51997 16535 52055 16541
rect 53190 16532 53196 16544
rect 53248 16572 53254 16584
rect 53484 16581 53512 16612
rect 57146 16600 57152 16612
rect 57204 16600 57210 16652
rect 53469 16575 53527 16581
rect 53248 16544 53420 16572
rect 53248 16532 53254 16544
rect 44450 16504 44456 16516
rect 43732 16476 44456 16504
rect 43073 16467 43131 16473
rect 31849 16439 31907 16445
rect 31849 16436 31861 16439
rect 29932 16408 31861 16436
rect 31849 16405 31861 16408
rect 31895 16436 31907 16439
rect 32490 16436 32496 16448
rect 31895 16408 32496 16436
rect 31895 16405 31907 16408
rect 31849 16399 31907 16405
rect 32490 16396 32496 16408
rect 32548 16396 32554 16448
rect 32674 16396 32680 16448
rect 32732 16436 32738 16448
rect 34514 16436 34520 16448
rect 32732 16408 34520 16436
rect 32732 16396 32738 16408
rect 34514 16396 34520 16408
rect 34572 16396 34578 16448
rect 35069 16439 35127 16445
rect 35069 16405 35081 16439
rect 35115 16436 35127 16439
rect 39206 16436 39212 16448
rect 35115 16408 39212 16436
rect 35115 16405 35127 16408
rect 35069 16399 35127 16405
rect 39206 16396 39212 16408
rect 39264 16396 39270 16448
rect 41966 16396 41972 16448
rect 42024 16436 42030 16448
rect 42337 16439 42395 16445
rect 42337 16436 42349 16439
rect 42024 16408 42349 16436
rect 42024 16396 42030 16408
rect 42337 16405 42349 16408
rect 42383 16436 42395 16439
rect 43088 16436 43116 16467
rect 44450 16464 44456 16476
rect 44508 16464 44514 16516
rect 42383 16408 43116 16436
rect 43165 16439 43223 16445
rect 42383 16405 42395 16408
rect 42337 16399 42395 16405
rect 43165 16405 43177 16439
rect 43211 16436 43223 16439
rect 43806 16436 43812 16448
rect 43211 16408 43812 16436
rect 43211 16405 43223 16408
rect 43165 16399 43223 16405
rect 43806 16396 43812 16408
rect 43864 16396 43870 16448
rect 53098 16396 53104 16448
rect 53156 16436 53162 16448
rect 53285 16439 53343 16445
rect 53285 16436 53297 16439
rect 53156 16408 53297 16436
rect 53156 16396 53162 16408
rect 53285 16405 53297 16408
rect 53331 16405 53343 16439
rect 53392 16436 53420 16544
rect 53469 16541 53481 16575
rect 53515 16574 53527 16575
rect 53515 16546 53549 16574
rect 56226 16572 56232 16584
rect 53515 16541 53527 16546
rect 56187 16544 56232 16572
rect 53469 16535 53527 16541
rect 53484 16504 53512 16535
rect 56226 16532 56232 16544
rect 56284 16532 56290 16584
rect 56318 16532 56324 16584
rect 56376 16572 56382 16584
rect 56413 16575 56471 16581
rect 56413 16572 56425 16575
rect 56376 16544 56425 16572
rect 56376 16532 56382 16544
rect 56413 16541 56425 16544
rect 56459 16541 56471 16575
rect 58158 16572 58164 16584
rect 58119 16544 58164 16572
rect 56413 16535 56471 16541
rect 58158 16532 58164 16544
rect 58216 16532 58222 16584
rect 54481 16507 54539 16513
rect 54481 16504 54493 16507
rect 53484 16476 54493 16504
rect 54481 16473 54493 16476
rect 54527 16473 54539 16507
rect 57885 16507 57943 16513
rect 57885 16504 57897 16507
rect 54481 16467 54539 16473
rect 57716 16476 57897 16504
rect 57716 16448 57744 16476
rect 57885 16473 57897 16476
rect 57931 16473 57943 16507
rect 57885 16467 57943 16473
rect 54271 16439 54329 16445
rect 54271 16436 54283 16439
rect 53392 16408 54283 16436
rect 53285 16399 53343 16405
rect 54271 16405 54283 16408
rect 54317 16405 54329 16439
rect 54271 16399 54329 16405
rect 57698 16396 57704 16448
rect 57756 16396 57762 16448
rect 1104 16346 58880 16368
rect 1104 16294 19574 16346
rect 19626 16294 19638 16346
rect 19690 16294 19702 16346
rect 19754 16294 19766 16346
rect 19818 16294 19830 16346
rect 19882 16294 50294 16346
rect 50346 16294 50358 16346
rect 50410 16294 50422 16346
rect 50474 16294 50486 16346
rect 50538 16294 50550 16346
rect 50602 16294 58880 16346
rect 1104 16272 58880 16294
rect 1762 16232 1768 16244
rect 1723 16204 1768 16232
rect 1762 16192 1768 16204
rect 1820 16192 1826 16244
rect 3697 16235 3755 16241
rect 3697 16201 3709 16235
rect 3743 16232 3755 16235
rect 4154 16232 4160 16244
rect 3743 16204 4160 16232
rect 3743 16201 3755 16204
rect 3697 16195 3755 16201
rect 4154 16192 4160 16204
rect 4212 16192 4218 16244
rect 8202 16232 8208 16244
rect 8163 16204 8208 16232
rect 8202 16192 8208 16204
rect 8260 16192 8266 16244
rect 8662 16192 8668 16244
rect 8720 16232 8726 16244
rect 9125 16235 9183 16241
rect 9125 16232 9137 16235
rect 8720 16204 9137 16232
rect 8720 16192 8726 16204
rect 9125 16201 9137 16204
rect 9171 16232 9183 16235
rect 9306 16232 9312 16244
rect 9171 16204 9312 16232
rect 9171 16201 9183 16204
rect 9125 16195 9183 16201
rect 9306 16192 9312 16204
rect 9364 16232 9370 16244
rect 9582 16232 9588 16244
rect 9364 16204 9588 16232
rect 9364 16192 9370 16204
rect 9582 16192 9588 16204
rect 9640 16192 9646 16244
rect 13538 16232 13544 16244
rect 12820 16204 13544 16232
rect 1780 16096 1808 16192
rect 2682 16164 2688 16176
rect 2424 16136 2688 16164
rect 2424 16105 2452 16136
rect 2682 16124 2688 16136
rect 2740 16164 2746 16176
rect 3329 16167 3387 16173
rect 3329 16164 3341 16167
rect 2740 16136 3341 16164
rect 2740 16124 2746 16136
rect 3329 16133 3341 16136
rect 3375 16133 3387 16167
rect 8220 16164 8248 16192
rect 9493 16167 9551 16173
rect 8220 16136 9444 16164
rect 3329 16127 3387 16133
rect 2409 16099 2467 16105
rect 2409 16096 2421 16099
rect 1780 16068 2421 16096
rect 2409 16065 2421 16068
rect 2455 16065 2467 16099
rect 2774 16096 2780 16108
rect 2409 16059 2467 16065
rect 2746 16056 2780 16096
rect 2832 16096 2838 16108
rect 3237 16099 3295 16105
rect 3237 16096 3249 16099
rect 2832 16068 3249 16096
rect 2832 16056 2838 16068
rect 3237 16065 3249 16068
rect 3283 16065 3295 16099
rect 3510 16096 3516 16108
rect 3471 16068 3516 16096
rect 3237 16059 3295 16065
rect 3510 16056 3516 16068
rect 3568 16056 3574 16108
rect 7190 16096 7196 16108
rect 7151 16068 7196 16096
rect 7190 16056 7196 16068
rect 7248 16056 7254 16108
rect 7558 16096 7564 16108
rect 7519 16068 7564 16096
rect 7558 16056 7564 16068
rect 7616 16056 7622 16108
rect 8021 16099 8079 16105
rect 8021 16065 8033 16099
rect 8067 16096 8079 16099
rect 8110 16096 8116 16108
rect 8067 16068 8116 16096
rect 8067 16065 8079 16068
rect 8021 16059 8079 16065
rect 8110 16056 8116 16068
rect 8168 16056 8174 16108
rect 9030 16096 9036 16108
rect 8991 16068 9036 16096
rect 9030 16056 9036 16068
rect 9088 16056 9094 16108
rect 9214 16056 9220 16108
rect 9272 16096 9278 16108
rect 9309 16099 9367 16105
rect 9309 16096 9321 16099
rect 9272 16068 9321 16096
rect 9272 16056 9278 16068
rect 9309 16065 9321 16068
rect 9355 16065 9367 16099
rect 9416 16096 9444 16136
rect 9493 16133 9505 16167
rect 9539 16164 9551 16167
rect 12434 16164 12440 16176
rect 9539 16136 10548 16164
rect 9539 16133 9551 16136
rect 9493 16127 9551 16133
rect 9950 16096 9956 16108
rect 9416 16068 9674 16096
rect 9911 16068 9956 16096
rect 9309 16059 9367 16065
rect 2501 16031 2559 16037
rect 2501 15997 2513 16031
rect 2547 16028 2559 16031
rect 2746 16028 2774 16056
rect 2547 16000 2774 16028
rect 9646 16028 9674 16068
rect 9950 16056 9956 16068
rect 10008 16056 10014 16108
rect 10520 16105 10548 16136
rect 12406 16124 12440 16164
rect 12492 16124 12498 16176
rect 10505 16099 10563 16105
rect 10505 16065 10517 16099
rect 10551 16096 10563 16099
rect 10962 16096 10968 16108
rect 10551 16068 10968 16096
rect 10551 16065 10563 16068
rect 10505 16059 10563 16065
rect 10962 16056 10968 16068
rect 11020 16056 11026 16108
rect 10042 16028 10048 16040
rect 9646 16000 10048 16028
rect 2547 15997 2559 16000
rect 2501 15991 2559 15997
rect 10042 15988 10048 16000
rect 10100 15988 10106 16040
rect 10321 16031 10379 16037
rect 10321 15997 10333 16031
rect 10367 16028 10379 16031
rect 12406 16028 12434 16124
rect 12820 16096 12848 16204
rect 13538 16192 13544 16204
rect 13596 16192 13602 16244
rect 21266 16232 21272 16244
rect 19720 16204 21272 16232
rect 12989 16167 13047 16173
rect 12989 16133 13001 16167
rect 13035 16164 13047 16167
rect 13630 16164 13636 16176
rect 13035 16136 13636 16164
rect 13035 16133 13047 16136
rect 12989 16127 13047 16133
rect 13630 16124 13636 16136
rect 13688 16164 13694 16176
rect 14277 16167 14335 16173
rect 14277 16164 14289 16167
rect 13688 16136 14289 16164
rect 13688 16124 13694 16136
rect 14277 16133 14289 16136
rect 14323 16133 14335 16167
rect 17310 16164 17316 16176
rect 14277 16127 14335 16133
rect 14384 16136 17316 16164
rect 12887 16099 12945 16105
rect 12887 16096 12899 16099
rect 12820 16068 12899 16096
rect 12887 16065 12899 16068
rect 12933 16065 12945 16099
rect 12887 16059 12945 16065
rect 13081 16099 13139 16105
rect 13081 16065 13093 16099
rect 13127 16096 13139 16099
rect 14182 16096 14188 16108
rect 13127 16068 14188 16096
rect 13127 16065 13139 16068
rect 13081 16059 13139 16065
rect 13096 16028 13124 16059
rect 14182 16056 14188 16068
rect 14240 16056 14246 16108
rect 10367 16000 10548 16028
rect 10367 15997 10379 16000
rect 10321 15991 10379 15997
rect 10520 15972 10548 16000
rect 10612 16000 13124 16028
rect 2777 15963 2835 15969
rect 2777 15929 2789 15963
rect 2823 15960 2835 15963
rect 2866 15960 2872 15972
rect 2823 15932 2872 15960
rect 2823 15929 2835 15932
rect 2777 15923 2835 15929
rect 2866 15920 2872 15932
rect 2924 15960 2930 15972
rect 3786 15960 3792 15972
rect 2924 15932 3792 15960
rect 2924 15920 2930 15932
rect 3786 15920 3792 15932
rect 3844 15920 3850 15972
rect 6914 15920 6920 15972
rect 6972 15960 6978 15972
rect 6972 15932 10456 15960
rect 6972 15920 6978 15932
rect 10428 15892 10456 15932
rect 10502 15920 10508 15972
rect 10560 15920 10566 15972
rect 10612 15892 10640 16000
rect 13354 15988 13360 16040
rect 13412 16028 13418 16040
rect 14384 16028 14412 16136
rect 17310 16124 17316 16136
rect 17368 16124 17374 16176
rect 17954 16124 17960 16176
rect 18012 16164 18018 16176
rect 19720 16164 19748 16204
rect 21266 16192 21272 16204
rect 21324 16192 21330 16244
rect 23661 16235 23719 16241
rect 23661 16201 23673 16235
rect 23707 16232 23719 16235
rect 26234 16232 26240 16244
rect 23707 16204 26240 16232
rect 23707 16201 23719 16204
rect 23661 16195 23719 16201
rect 26234 16192 26240 16204
rect 26292 16192 26298 16244
rect 26418 16192 26424 16244
rect 26476 16232 26482 16244
rect 27157 16235 27215 16241
rect 27157 16232 27169 16235
rect 26476 16204 27169 16232
rect 26476 16192 26482 16204
rect 27157 16201 27169 16204
rect 27203 16201 27215 16235
rect 27614 16232 27620 16244
rect 27157 16195 27215 16201
rect 27356 16204 27620 16232
rect 18012 16136 19748 16164
rect 18012 16124 18018 16136
rect 15838 16056 15844 16108
rect 15896 16096 15902 16108
rect 15933 16099 15991 16105
rect 15933 16096 15945 16099
rect 15896 16068 15945 16096
rect 15896 16056 15902 16068
rect 15933 16065 15945 16068
rect 15979 16065 15991 16099
rect 16114 16096 16120 16108
rect 16075 16068 16120 16096
rect 15933 16059 15991 16065
rect 16114 16056 16120 16068
rect 16172 16056 16178 16108
rect 17129 16099 17187 16105
rect 17129 16065 17141 16099
rect 17175 16096 17187 16099
rect 19334 16096 19340 16108
rect 17175 16068 19340 16096
rect 17175 16065 17187 16068
rect 17129 16059 17187 16065
rect 19334 16056 19340 16068
rect 19392 16056 19398 16108
rect 19610 16096 19616 16108
rect 19571 16068 19616 16096
rect 19610 16056 19616 16068
rect 19668 16056 19674 16108
rect 19720 16105 19748 16136
rect 19889 16167 19947 16173
rect 19889 16133 19901 16167
rect 19935 16164 19947 16167
rect 20438 16164 20444 16176
rect 19935 16136 20444 16164
rect 19935 16133 19947 16136
rect 19889 16127 19947 16133
rect 20438 16124 20444 16136
rect 20496 16164 20502 16176
rect 20990 16164 20996 16176
rect 20496 16136 20996 16164
rect 20496 16124 20502 16136
rect 20990 16124 20996 16136
rect 21048 16124 21054 16176
rect 22370 16124 22376 16176
rect 22428 16164 22434 16176
rect 22428 16136 23525 16164
rect 22428 16124 22434 16136
rect 20162 16105 20168 16108
rect 19706 16099 19764 16105
rect 19706 16065 19718 16099
rect 19752 16065 19764 16099
rect 19706 16059 19764 16065
rect 19981 16099 20039 16105
rect 19981 16065 19993 16099
rect 20027 16065 20039 16099
rect 19981 16059 20039 16065
rect 20119 16099 20168 16105
rect 20119 16065 20131 16099
rect 20165 16065 20168 16099
rect 20119 16059 20168 16065
rect 13412 16000 14412 16028
rect 14461 16031 14519 16037
rect 13412 15988 13418 16000
rect 14461 15997 14473 16031
rect 14507 16028 14519 16031
rect 14918 16028 14924 16040
rect 14507 16000 14924 16028
rect 14507 15997 14519 16000
rect 14461 15991 14519 15997
rect 14918 15988 14924 16000
rect 14976 16028 14982 16040
rect 16132 16028 16160 16056
rect 14976 16000 16160 16028
rect 14976 15988 14982 16000
rect 11330 15920 11336 15972
rect 11388 15960 11394 15972
rect 19426 15960 19432 15972
rect 11388 15932 19432 15960
rect 11388 15920 11394 15932
rect 19426 15920 19432 15932
rect 19484 15920 19490 15972
rect 10428 15864 10640 15892
rect 15197 15895 15255 15901
rect 15197 15861 15209 15895
rect 15243 15892 15255 15895
rect 15286 15892 15292 15904
rect 15243 15864 15292 15892
rect 15243 15861 15255 15864
rect 15197 15855 15255 15861
rect 15286 15852 15292 15864
rect 15344 15852 15350 15904
rect 16117 15895 16175 15901
rect 16117 15861 16129 15895
rect 16163 15892 16175 15895
rect 16390 15892 16396 15904
rect 16163 15864 16396 15892
rect 16163 15861 16175 15864
rect 16117 15855 16175 15861
rect 16390 15852 16396 15864
rect 16448 15852 16454 15904
rect 16850 15852 16856 15904
rect 16908 15892 16914 15904
rect 17221 15895 17279 15901
rect 17221 15892 17233 15895
rect 16908 15864 17233 15892
rect 16908 15852 16914 15864
rect 17221 15861 17233 15864
rect 17267 15861 17279 15895
rect 17221 15855 17279 15861
rect 18874 15852 18880 15904
rect 18932 15892 18938 15904
rect 19058 15892 19064 15904
rect 18932 15864 19064 15892
rect 18932 15852 18938 15864
rect 19058 15852 19064 15864
rect 19116 15892 19122 15904
rect 19996 15892 20024 16059
rect 20162 16056 20168 16059
rect 20220 16096 20226 16108
rect 20622 16096 20628 16108
rect 20220 16068 20628 16096
rect 20220 16056 20226 16068
rect 20622 16056 20628 16068
rect 20680 16056 20686 16108
rect 22830 16056 22836 16108
rect 22888 16096 22894 16108
rect 23017 16099 23075 16105
rect 23017 16096 23029 16099
rect 22888 16068 23029 16096
rect 22888 16056 22894 16068
rect 23017 16065 23029 16068
rect 23063 16065 23075 16099
rect 23017 16059 23075 16065
rect 23110 16099 23168 16105
rect 23110 16065 23122 16099
rect 23156 16065 23168 16099
rect 23290 16096 23296 16108
rect 23251 16068 23296 16096
rect 23110 16059 23168 16065
rect 21726 15988 21732 16040
rect 21784 16028 21790 16040
rect 23124 16028 23152 16059
rect 23290 16056 23296 16068
rect 23348 16056 23354 16108
rect 23497 16105 23525 16136
rect 25038 16124 25044 16176
rect 25096 16164 25102 16176
rect 26329 16167 26387 16173
rect 26329 16164 26341 16167
rect 25096 16136 26341 16164
rect 25096 16124 25102 16136
rect 26329 16133 26341 16136
rect 26375 16164 26387 16167
rect 26510 16164 26516 16176
rect 26375 16136 26516 16164
rect 26375 16133 26387 16136
rect 26329 16127 26387 16133
rect 26510 16124 26516 16136
rect 26568 16164 26574 16176
rect 27246 16164 27252 16176
rect 26568 16136 27252 16164
rect 26568 16124 26574 16136
rect 27246 16124 27252 16136
rect 27304 16124 27310 16176
rect 23385 16099 23443 16105
rect 23385 16065 23397 16099
rect 23431 16065 23443 16099
rect 23385 16059 23443 16065
rect 23482 16099 23540 16105
rect 23482 16065 23494 16099
rect 23528 16065 23540 16099
rect 23482 16059 23540 16065
rect 21784 16000 23152 16028
rect 21784 15988 21790 16000
rect 23198 15988 23204 16040
rect 23256 16028 23262 16040
rect 23400 16028 23428 16059
rect 24118 16056 24124 16108
rect 24176 16096 24182 16108
rect 24213 16099 24271 16105
rect 24213 16096 24225 16099
rect 24176 16068 24225 16096
rect 24176 16056 24182 16068
rect 24213 16065 24225 16068
rect 24259 16065 24271 16099
rect 24213 16059 24271 16065
rect 24946 16056 24952 16108
rect 25004 16096 25010 16108
rect 27356 16105 27384 16204
rect 27614 16192 27620 16204
rect 27672 16192 27678 16244
rect 27706 16192 27712 16244
rect 27764 16232 27770 16244
rect 32490 16232 32496 16244
rect 27764 16204 30420 16232
rect 32451 16204 32496 16232
rect 27764 16192 27770 16204
rect 27525 16167 27583 16173
rect 27525 16133 27537 16167
rect 27571 16164 27583 16167
rect 28074 16164 28080 16176
rect 27571 16136 28080 16164
rect 27571 16133 27583 16136
rect 27525 16127 27583 16133
rect 28074 16124 28080 16136
rect 28132 16124 28138 16176
rect 28442 16164 28448 16176
rect 28403 16136 28448 16164
rect 28442 16124 28448 16136
rect 28500 16124 28506 16176
rect 29178 16164 29184 16176
rect 29139 16136 29184 16164
rect 29178 16124 29184 16136
rect 29236 16124 29242 16176
rect 27341 16099 27399 16105
rect 25004 16068 27292 16096
rect 25004 16056 25010 16068
rect 25038 16028 25044 16040
rect 23256 16000 25044 16028
rect 23256 15988 23262 16000
rect 25038 15988 25044 16000
rect 25096 15988 25102 16040
rect 27264 16028 27292 16068
rect 27341 16065 27353 16099
rect 27387 16065 27399 16099
rect 27341 16059 27399 16065
rect 27430 16056 27436 16108
rect 27488 16096 27494 16108
rect 27709 16099 27767 16105
rect 27709 16096 27721 16099
rect 27488 16068 27533 16096
rect 27632 16068 27721 16096
rect 27488 16056 27494 16068
rect 27632 16028 27660 16068
rect 27709 16065 27721 16068
rect 27755 16065 27767 16099
rect 27709 16059 27767 16065
rect 28166 16056 28172 16108
rect 28224 16096 28230 16108
rect 28261 16099 28319 16105
rect 28261 16096 28273 16099
rect 28224 16068 28273 16096
rect 28224 16056 28230 16068
rect 28261 16065 28273 16068
rect 28307 16096 28319 16099
rect 28905 16099 28963 16105
rect 28905 16096 28917 16099
rect 28307 16068 28917 16096
rect 28307 16065 28319 16068
rect 28261 16059 28319 16065
rect 28905 16065 28917 16068
rect 28951 16065 28963 16099
rect 28905 16059 28963 16065
rect 28997 16099 29055 16105
rect 28997 16065 29009 16099
rect 29043 16096 29055 16099
rect 29086 16096 29092 16108
rect 29043 16068 29092 16096
rect 29043 16065 29055 16068
rect 28997 16059 29055 16065
rect 29086 16056 29092 16068
rect 29144 16056 29150 16108
rect 29638 16056 29644 16108
rect 29696 16096 29702 16108
rect 30009 16099 30067 16105
rect 30009 16096 30021 16099
rect 29696 16068 30021 16096
rect 29696 16056 29702 16068
rect 30009 16065 30021 16068
rect 30055 16065 30067 16099
rect 30009 16059 30067 16065
rect 30285 16099 30343 16105
rect 30285 16065 30297 16099
rect 30331 16065 30343 16099
rect 30285 16059 30343 16065
rect 27264 16000 27660 16028
rect 20257 15963 20315 15969
rect 20257 15929 20269 15963
rect 20303 15929 20315 15963
rect 20257 15923 20315 15929
rect 19116 15864 20024 15892
rect 20272 15892 20300 15923
rect 20346 15920 20352 15972
rect 20404 15960 20410 15972
rect 20404 15932 22094 15960
rect 20404 15920 20410 15932
rect 20622 15892 20628 15904
rect 20272 15864 20628 15892
rect 19116 15852 19122 15864
rect 20622 15852 20628 15864
rect 20680 15852 20686 15904
rect 22066 15892 22094 15932
rect 22370 15920 22376 15972
rect 22428 15960 22434 15972
rect 22465 15963 22523 15969
rect 22465 15960 22477 15963
rect 22428 15932 22477 15960
rect 22428 15920 22434 15932
rect 22465 15929 22477 15932
rect 22511 15929 22523 15963
rect 25777 15963 25835 15969
rect 25777 15960 25789 15963
rect 22465 15923 22523 15929
rect 24412 15932 25789 15960
rect 24412 15892 24440 15932
rect 25777 15929 25789 15932
rect 25823 15929 25835 15963
rect 25777 15923 25835 15929
rect 29181 15963 29239 15969
rect 29181 15929 29193 15963
rect 29227 15960 29239 15963
rect 30300 15960 30328 16059
rect 29227 15932 30328 15960
rect 30392 15960 30420 16204
rect 32490 16192 32496 16204
rect 32548 16192 32554 16244
rect 34422 16192 34428 16244
rect 34480 16232 34486 16244
rect 34609 16235 34667 16241
rect 34609 16232 34621 16235
rect 34480 16204 34621 16232
rect 34480 16192 34486 16204
rect 34609 16201 34621 16204
rect 34655 16201 34667 16235
rect 34609 16195 34667 16201
rect 36633 16235 36691 16241
rect 36633 16201 36645 16235
rect 36679 16232 36691 16235
rect 43990 16232 43996 16244
rect 36679 16204 43996 16232
rect 36679 16201 36691 16204
rect 36633 16195 36691 16201
rect 43990 16192 43996 16204
rect 44048 16192 44054 16244
rect 53009 16235 53067 16241
rect 53009 16201 53021 16235
rect 53055 16232 53067 16235
rect 53190 16232 53196 16244
rect 53055 16204 53196 16232
rect 53055 16201 53067 16204
rect 53009 16195 53067 16201
rect 53190 16192 53196 16204
rect 53248 16192 53254 16244
rect 58158 16232 58164 16244
rect 58119 16204 58164 16232
rect 58158 16192 58164 16204
rect 58216 16192 58222 16244
rect 32508 16096 32536 16192
rect 33137 16099 33195 16105
rect 33137 16096 33149 16099
rect 32508 16068 33149 16096
rect 33137 16065 33149 16068
rect 33183 16065 33195 16099
rect 34440 16096 34468 16192
rect 35250 16124 35256 16176
rect 35308 16164 35314 16176
rect 36265 16167 36323 16173
rect 36265 16164 36277 16167
rect 35308 16136 36277 16164
rect 35308 16124 35314 16136
rect 36265 16133 36277 16136
rect 36311 16164 36323 16167
rect 38562 16164 38568 16176
rect 36311 16136 38568 16164
rect 36311 16133 36323 16136
rect 36265 16127 36323 16133
rect 38562 16124 38568 16136
rect 38620 16124 38626 16176
rect 43806 16124 43812 16176
rect 43864 16164 43870 16176
rect 43864 16136 44404 16164
rect 43864 16124 43870 16136
rect 33810 16068 34468 16096
rect 33137 16059 33195 16065
rect 34514 16056 34520 16108
rect 34572 16096 34578 16108
rect 35802 16096 35808 16108
rect 34572 16068 35808 16096
rect 34572 16056 34578 16068
rect 35802 16056 35808 16068
rect 35860 16096 35866 16108
rect 36081 16099 36139 16105
rect 36081 16096 36093 16099
rect 35860 16068 36093 16096
rect 35860 16056 35866 16068
rect 36081 16065 36093 16068
rect 36127 16065 36139 16099
rect 36354 16096 36360 16108
rect 36315 16068 36360 16096
rect 36081 16059 36139 16065
rect 36354 16056 36360 16068
rect 36412 16056 36418 16108
rect 36538 16105 36544 16108
rect 36495 16099 36544 16105
rect 36495 16065 36507 16099
rect 36541 16065 36544 16099
rect 36495 16059 36544 16065
rect 36538 16056 36544 16059
rect 36596 16056 36602 16108
rect 38654 16096 38660 16108
rect 38615 16068 38660 16096
rect 38654 16056 38660 16068
rect 38712 16056 38718 16108
rect 38930 16056 38936 16108
rect 38988 16096 38994 16108
rect 42794 16096 42800 16108
rect 38988 16068 42800 16096
rect 38988 16056 38994 16068
rect 42794 16056 42800 16068
rect 42852 16056 42858 16108
rect 43073 16099 43131 16105
rect 43073 16065 43085 16099
rect 43119 16096 43131 16099
rect 43254 16096 43260 16108
rect 43119 16068 43260 16096
rect 43119 16065 43131 16068
rect 43073 16059 43131 16065
rect 43254 16056 43260 16068
rect 43312 16056 43318 16108
rect 43898 16056 43904 16108
rect 43956 16096 43962 16108
rect 44376 16105 44404 16136
rect 56134 16124 56140 16176
rect 56192 16164 56198 16176
rect 56192 16136 56548 16164
rect 56192 16124 56198 16136
rect 44269 16099 44327 16105
rect 44269 16096 44281 16099
rect 43956 16068 44281 16096
rect 43956 16056 43962 16068
rect 44269 16065 44281 16068
rect 44315 16065 44327 16099
rect 44269 16059 44327 16065
rect 44361 16099 44419 16105
rect 44361 16065 44373 16099
rect 44407 16065 44419 16099
rect 44361 16059 44419 16065
rect 52733 16099 52791 16105
rect 52733 16065 52745 16099
rect 52779 16096 52791 16099
rect 52914 16096 52920 16108
rect 52779 16068 52920 16096
rect 52779 16065 52791 16068
rect 52733 16059 52791 16065
rect 52914 16056 52920 16068
rect 52972 16056 52978 16108
rect 56229 16099 56287 16105
rect 56229 16065 56241 16099
rect 56275 16096 56287 16099
rect 56318 16096 56324 16108
rect 56275 16068 56324 16096
rect 56275 16065 56287 16068
rect 56229 16059 56287 16065
rect 56318 16056 56324 16068
rect 56376 16056 56382 16108
rect 56520 16105 56548 16136
rect 56505 16099 56563 16105
rect 56505 16065 56517 16099
rect 56551 16065 56563 16099
rect 56505 16059 56563 16065
rect 56597 16099 56655 16105
rect 56597 16065 56609 16099
rect 56643 16096 56655 16099
rect 57146 16096 57152 16108
rect 56643 16068 57152 16096
rect 56643 16065 56655 16068
rect 56597 16059 56655 16065
rect 57146 16056 57152 16068
rect 57204 16056 57210 16108
rect 30469 16031 30527 16037
rect 30469 15997 30481 16031
rect 30515 16028 30527 16031
rect 34054 16028 34060 16040
rect 30515 16000 34060 16028
rect 30515 15997 30527 16000
rect 30469 15991 30527 15997
rect 34054 15988 34060 16000
rect 34112 15988 34118 16040
rect 34149 16031 34207 16037
rect 34149 15997 34161 16031
rect 34195 16028 34207 16031
rect 34330 16028 34336 16040
rect 34195 16000 34336 16028
rect 34195 15997 34207 16000
rect 34149 15991 34207 15997
rect 34330 15988 34336 16000
rect 34388 15988 34394 16040
rect 38565 16031 38623 16037
rect 38565 16028 38577 16031
rect 34440 16000 38577 16028
rect 30392 15932 33456 15960
rect 29227 15929 29239 15932
rect 29181 15923 29239 15929
rect 22066 15864 24440 15892
rect 24486 15852 24492 15904
rect 24544 15892 24550 15904
rect 24762 15892 24768 15904
rect 24544 15864 24768 15892
rect 24544 15852 24550 15864
rect 24762 15852 24768 15864
rect 24820 15852 24826 15904
rect 25792 15892 25820 15923
rect 26234 15892 26240 15904
rect 25792 15864 26240 15892
rect 26234 15852 26240 15864
rect 26292 15852 26298 15904
rect 29822 15852 29828 15904
rect 29880 15892 29886 15904
rect 30101 15895 30159 15901
rect 30101 15892 30113 15895
rect 29880 15864 30113 15892
rect 29880 15852 29886 15864
rect 30101 15861 30113 15864
rect 30147 15861 30159 15895
rect 33428 15892 33456 15932
rect 34440 15892 34468 16000
rect 38565 15997 38577 16000
rect 38611 15997 38623 16031
rect 38565 15991 38623 15997
rect 39485 16031 39543 16037
rect 39485 15997 39497 16031
rect 39531 16028 39543 16031
rect 39531 16000 41414 16028
rect 39531 15997 39543 16000
rect 39485 15991 39543 15997
rect 41386 15960 41414 16000
rect 44082 15988 44088 16040
rect 44140 16028 44146 16040
rect 44177 16031 44235 16037
rect 44177 16028 44189 16031
rect 44140 16000 44189 16028
rect 44140 15988 44146 16000
rect 44177 15997 44189 16000
rect 44223 15997 44235 16031
rect 44450 16028 44456 16040
rect 44411 16000 44456 16028
rect 44177 15991 44235 15997
rect 44450 15988 44456 16000
rect 44508 15988 44514 16040
rect 52822 15988 52828 16040
rect 52880 16028 52886 16040
rect 53009 16031 53067 16037
rect 53009 16028 53021 16031
rect 52880 16000 53021 16028
rect 52880 15988 52886 16000
rect 53009 15997 53021 16000
rect 53055 15997 53067 16031
rect 53009 15991 53067 15997
rect 48682 15960 48688 15972
rect 41386 15932 48688 15960
rect 48682 15920 48688 15932
rect 48740 15920 48746 15972
rect 33428 15864 34468 15892
rect 30101 15855 30159 15861
rect 39206 15852 39212 15904
rect 39264 15892 39270 15904
rect 44174 15892 44180 15904
rect 39264 15864 44180 15892
rect 39264 15852 39270 15864
rect 44174 15852 44180 15864
rect 44232 15852 44238 15904
rect 44637 15895 44695 15901
rect 44637 15861 44649 15895
rect 44683 15892 44695 15895
rect 47302 15892 47308 15904
rect 44683 15864 47308 15892
rect 44683 15861 44695 15864
rect 44637 15855 44695 15861
rect 47302 15852 47308 15864
rect 47360 15852 47366 15904
rect 52825 15895 52883 15901
rect 52825 15861 52837 15895
rect 52871 15892 52883 15895
rect 53006 15892 53012 15904
rect 52871 15864 53012 15892
rect 52871 15861 52883 15864
rect 52825 15855 52883 15861
rect 53006 15852 53012 15864
rect 53064 15852 53070 15904
rect 56318 15892 56324 15904
rect 56279 15864 56324 15892
rect 56318 15852 56324 15864
rect 56376 15852 56382 15904
rect 56778 15892 56784 15904
rect 56739 15864 56784 15892
rect 56778 15852 56784 15864
rect 56836 15852 56842 15904
rect 1104 15802 58880 15824
rect 1104 15750 4214 15802
rect 4266 15750 4278 15802
rect 4330 15750 4342 15802
rect 4394 15750 4406 15802
rect 4458 15750 4470 15802
rect 4522 15750 34934 15802
rect 34986 15750 34998 15802
rect 35050 15750 35062 15802
rect 35114 15750 35126 15802
rect 35178 15750 35190 15802
rect 35242 15750 58880 15802
rect 1104 15728 58880 15750
rect 2682 15648 2688 15700
rect 2740 15688 2746 15700
rect 3053 15691 3111 15697
rect 3053 15688 3065 15691
rect 2740 15660 3065 15688
rect 2740 15648 2746 15660
rect 3053 15657 3065 15660
rect 3099 15657 3111 15691
rect 3053 15651 3111 15657
rect 9030 15648 9036 15700
rect 9088 15688 9094 15700
rect 10045 15691 10103 15697
rect 9088 15660 9996 15688
rect 9088 15648 9094 15660
rect 7837 15623 7895 15629
rect 7837 15589 7849 15623
rect 7883 15620 7895 15623
rect 9674 15620 9680 15632
rect 7883 15592 9680 15620
rect 7883 15589 7895 15592
rect 7837 15583 7895 15589
rect 9674 15580 9680 15592
rect 9732 15580 9738 15632
rect 9214 15512 9220 15564
rect 9272 15552 9278 15564
rect 9272 15524 9628 15552
rect 9272 15512 9278 15524
rect 3786 15484 3792 15496
rect 3747 15456 3792 15484
rect 3786 15444 3792 15456
rect 3844 15444 3850 15496
rect 3973 15487 4031 15493
rect 3973 15453 3985 15487
rect 4019 15484 4031 15487
rect 4614 15484 4620 15496
rect 4019 15456 4620 15484
rect 4019 15453 4031 15456
rect 3973 15447 4031 15453
rect 4614 15444 4620 15456
rect 4672 15444 4678 15496
rect 6914 15484 6920 15496
rect 6875 15456 6920 15484
rect 6914 15444 6920 15456
rect 6972 15444 6978 15496
rect 7377 15487 7435 15493
rect 7377 15453 7389 15487
rect 7423 15453 7435 15487
rect 7742 15484 7748 15496
rect 7703 15456 7748 15484
rect 7377 15447 7435 15453
rect 7392 15416 7420 15447
rect 7742 15444 7748 15456
rect 7800 15444 7806 15496
rect 9600 15493 9628 15524
rect 9493 15487 9551 15493
rect 9493 15453 9505 15487
rect 9539 15453 9551 15487
rect 9493 15447 9551 15453
rect 9585 15487 9643 15493
rect 9585 15453 9597 15487
rect 9631 15453 9643 15487
rect 9585 15447 9643 15453
rect 9508 15416 9536 15447
rect 9674 15444 9680 15496
rect 9732 15478 9738 15496
rect 9769 15487 9827 15493
rect 9769 15478 9781 15487
rect 9732 15453 9781 15478
rect 9815 15453 9827 15487
rect 9732 15450 9827 15453
rect 9732 15444 9738 15450
rect 9769 15447 9827 15450
rect 9861 15487 9919 15493
rect 9861 15453 9873 15487
rect 9907 15484 9919 15487
rect 9968 15484 9996 15660
rect 10045 15657 10057 15691
rect 10091 15688 10103 15691
rect 13722 15688 13728 15700
rect 10091 15660 13728 15688
rect 10091 15657 10103 15660
rect 10045 15651 10103 15657
rect 13722 15648 13728 15660
rect 13780 15648 13786 15700
rect 14461 15691 14519 15697
rect 14461 15657 14473 15691
rect 14507 15688 14519 15691
rect 14550 15688 14556 15700
rect 14507 15660 14556 15688
rect 14507 15657 14519 15660
rect 14461 15651 14519 15657
rect 14550 15648 14556 15660
rect 14608 15648 14614 15700
rect 14642 15648 14648 15700
rect 14700 15688 14706 15700
rect 14700 15660 19334 15688
rect 14700 15648 14706 15660
rect 10594 15580 10600 15632
rect 10652 15620 10658 15632
rect 13354 15620 13360 15632
rect 10652 15592 13360 15620
rect 10652 15580 10658 15592
rect 13354 15580 13360 15592
rect 13412 15580 13418 15632
rect 13538 15620 13544 15632
rect 13499 15592 13544 15620
rect 13538 15580 13544 15592
rect 13596 15580 13602 15632
rect 11330 15552 11336 15564
rect 10612 15524 11336 15552
rect 9907 15456 9996 15484
rect 9907 15453 9919 15456
rect 9861 15447 9919 15453
rect 10042 15444 10048 15496
rect 10100 15484 10106 15496
rect 10612 15493 10640 15524
rect 11330 15512 11336 15524
rect 11388 15512 11394 15564
rect 11885 15555 11943 15561
rect 11885 15521 11897 15555
rect 11931 15552 11943 15555
rect 14642 15552 14648 15564
rect 11931 15524 14648 15552
rect 11931 15521 11943 15524
rect 11885 15515 11943 15521
rect 10597 15487 10655 15493
rect 10597 15484 10609 15487
rect 10100 15456 10609 15484
rect 10100 15444 10106 15456
rect 10597 15453 10609 15456
rect 10643 15453 10655 15487
rect 10597 15447 10655 15453
rect 10778 15444 10784 15496
rect 10836 15484 10842 15496
rect 11900 15484 11928 15515
rect 14642 15512 14648 15524
rect 14700 15512 14706 15564
rect 19306 15552 19334 15660
rect 19610 15648 19616 15700
rect 19668 15688 19674 15700
rect 19797 15691 19855 15697
rect 19797 15688 19809 15691
rect 19668 15660 19809 15688
rect 19668 15648 19674 15660
rect 19797 15657 19809 15660
rect 19843 15657 19855 15691
rect 22830 15688 22836 15700
rect 22791 15660 22836 15688
rect 19797 15651 19855 15657
rect 22830 15648 22836 15660
rect 22888 15648 22894 15700
rect 26789 15691 26847 15697
rect 26789 15657 26801 15691
rect 26835 15688 26847 15691
rect 26878 15688 26884 15700
rect 26835 15660 26884 15688
rect 26835 15657 26847 15660
rect 26789 15651 26847 15657
rect 26878 15648 26884 15660
rect 26936 15648 26942 15700
rect 27430 15648 27436 15700
rect 27488 15688 27494 15700
rect 29086 15688 29092 15700
rect 27488 15660 29092 15688
rect 27488 15648 27494 15660
rect 29086 15648 29092 15660
rect 29144 15648 29150 15700
rect 29638 15648 29644 15700
rect 29696 15688 29702 15700
rect 29825 15691 29883 15697
rect 29825 15688 29837 15691
rect 29696 15660 29837 15688
rect 29696 15648 29702 15660
rect 29825 15657 29837 15660
rect 29871 15657 29883 15691
rect 31018 15688 31024 15700
rect 30979 15660 31024 15688
rect 29825 15651 29883 15657
rect 31018 15648 31024 15660
rect 31076 15688 31082 15700
rect 32030 15688 32036 15700
rect 31076 15660 32036 15688
rect 31076 15648 31082 15660
rect 32030 15648 32036 15660
rect 32088 15688 32094 15700
rect 32398 15688 32404 15700
rect 32088 15660 32404 15688
rect 32088 15648 32094 15660
rect 32398 15648 32404 15660
rect 32456 15648 32462 15700
rect 39850 15688 39856 15700
rect 39811 15660 39856 15688
rect 39850 15648 39856 15660
rect 39908 15648 39914 15700
rect 43806 15648 43812 15700
rect 43864 15688 43870 15700
rect 44085 15691 44143 15697
rect 44085 15688 44097 15691
rect 43864 15660 44097 15688
rect 43864 15648 43870 15660
rect 44085 15657 44097 15660
rect 44131 15657 44143 15691
rect 44085 15651 44143 15657
rect 46569 15691 46627 15697
rect 46569 15657 46581 15691
rect 46615 15657 46627 15691
rect 46569 15651 46627 15657
rect 46753 15691 46811 15697
rect 46753 15657 46765 15691
rect 46799 15688 46811 15691
rect 52546 15688 52552 15700
rect 46799 15660 52552 15688
rect 46799 15657 46811 15660
rect 46753 15651 46811 15657
rect 19426 15580 19432 15632
rect 19484 15620 19490 15632
rect 20070 15620 20076 15632
rect 19484 15592 20076 15620
rect 19484 15580 19490 15592
rect 20070 15580 20076 15592
rect 20128 15580 20134 15632
rect 20438 15580 20444 15632
rect 20496 15620 20502 15632
rect 20898 15620 20904 15632
rect 20496 15592 20904 15620
rect 20496 15580 20502 15592
rect 20898 15580 20904 15592
rect 20956 15580 20962 15632
rect 23750 15620 23756 15632
rect 23032 15592 23756 15620
rect 20346 15552 20352 15564
rect 19306 15524 20352 15552
rect 20346 15512 20352 15524
rect 20404 15512 20410 15564
rect 14182 15484 14188 15496
rect 10836 15456 11928 15484
rect 14143 15456 14188 15484
rect 10836 15444 10842 15456
rect 14182 15444 14188 15456
rect 14240 15444 14246 15496
rect 14277 15487 14335 15493
rect 14277 15453 14289 15487
rect 14323 15453 14335 15487
rect 14277 15447 14335 15453
rect 10410 15416 10416 15428
rect 7392 15388 8984 15416
rect 9508 15388 10416 15416
rect 8956 15360 8984 15388
rect 10410 15376 10416 15388
rect 10468 15376 10474 15428
rect 13538 15376 13544 15428
rect 13596 15416 13602 15428
rect 14292 15416 14320 15447
rect 14458 15444 14464 15496
rect 14516 15484 14522 15496
rect 15102 15484 15108 15496
rect 14516 15456 15108 15484
rect 14516 15444 14522 15456
rect 15102 15444 15108 15456
rect 15160 15444 15166 15496
rect 15381 15487 15439 15493
rect 15381 15453 15393 15487
rect 15427 15484 15439 15487
rect 15470 15484 15476 15496
rect 15427 15456 15476 15484
rect 15427 15453 15439 15456
rect 15381 15447 15439 15453
rect 15470 15444 15476 15456
rect 15528 15484 15534 15496
rect 15746 15484 15752 15496
rect 15528 15456 15752 15484
rect 15528 15444 15534 15456
rect 15746 15444 15752 15456
rect 15804 15444 15810 15496
rect 16390 15484 16396 15496
rect 16351 15456 16396 15484
rect 16390 15444 16396 15456
rect 16448 15444 16454 15496
rect 16574 15493 16580 15496
rect 16541 15487 16580 15493
rect 16541 15453 16553 15487
rect 16541 15447 16580 15453
rect 16574 15444 16580 15447
rect 16632 15444 16638 15496
rect 16942 15493 16948 15496
rect 16899 15487 16948 15493
rect 16899 15453 16911 15487
rect 16945 15453 16948 15487
rect 16899 15447 16948 15453
rect 16942 15444 16948 15447
rect 17000 15444 17006 15496
rect 19245 15487 19303 15493
rect 19245 15453 19257 15487
rect 19291 15484 19303 15487
rect 19334 15484 19340 15496
rect 19291 15456 19340 15484
rect 19291 15453 19303 15456
rect 19245 15447 19303 15453
rect 19334 15444 19340 15456
rect 19392 15444 19398 15496
rect 19426 15444 19432 15496
rect 19484 15484 19490 15496
rect 19613 15487 19671 15493
rect 19484 15456 19529 15484
rect 19484 15444 19490 15456
rect 19613 15453 19625 15487
rect 19659 15484 19671 15487
rect 20254 15484 20260 15496
rect 19659 15456 20260 15484
rect 19659 15453 19671 15456
rect 19613 15447 19671 15453
rect 20254 15444 20260 15456
rect 20312 15484 20318 15496
rect 20441 15487 20499 15493
rect 20441 15484 20453 15487
rect 20312 15456 20453 15484
rect 20312 15444 20318 15456
rect 20441 15453 20453 15456
rect 20487 15453 20499 15487
rect 20441 15447 20499 15453
rect 21361 15487 21419 15493
rect 21361 15453 21373 15487
rect 21407 15484 21419 15487
rect 21726 15484 21732 15496
rect 21407 15456 21732 15484
rect 21407 15453 21419 15456
rect 21361 15447 21419 15453
rect 13596 15388 14320 15416
rect 15764 15416 15792 15444
rect 16669 15419 16727 15425
rect 16669 15416 16681 15419
rect 15764 15388 16681 15416
rect 13596 15376 13602 15388
rect 16669 15385 16681 15388
rect 16715 15385 16727 15419
rect 16669 15379 16727 15385
rect 16758 15376 16764 15428
rect 16816 15416 16822 15428
rect 19521 15419 19579 15425
rect 16816 15388 16861 15416
rect 16816 15376 16822 15388
rect 19521 15385 19533 15419
rect 19567 15416 19579 15419
rect 21376 15416 21404 15447
rect 21726 15444 21732 15456
rect 21784 15444 21790 15496
rect 23032 15493 23060 15592
rect 23750 15580 23756 15592
rect 23808 15620 23814 15632
rect 24302 15620 24308 15632
rect 23808 15592 24308 15620
rect 23808 15580 23814 15592
rect 24302 15580 24308 15592
rect 24360 15580 24366 15632
rect 24397 15623 24455 15629
rect 24397 15589 24409 15623
rect 24443 15620 24455 15623
rect 24762 15620 24768 15632
rect 24443 15592 24768 15620
rect 24443 15589 24455 15592
rect 24397 15583 24455 15589
rect 24762 15580 24768 15592
rect 24820 15580 24826 15632
rect 30834 15580 30840 15632
rect 30892 15620 30898 15632
rect 36354 15620 36360 15632
rect 30892 15592 36360 15620
rect 30892 15580 30898 15592
rect 36354 15580 36360 15592
rect 36412 15620 36418 15632
rect 37366 15620 37372 15632
rect 36412 15592 37372 15620
rect 36412 15580 36418 15592
rect 37366 15580 37372 15592
rect 37424 15580 37430 15632
rect 23474 15552 23480 15564
rect 23308 15524 23480 15552
rect 23017 15487 23075 15493
rect 23017 15453 23029 15487
rect 23063 15453 23075 15487
rect 23017 15447 23075 15453
rect 23106 15416 23112 15428
rect 19567 15388 21404 15416
rect 23067 15388 23112 15416
rect 19567 15385 19579 15388
rect 19521 15379 19579 15385
rect 23106 15376 23112 15388
rect 23164 15376 23170 15428
rect 23201 15419 23259 15425
rect 23201 15385 23213 15419
rect 23247 15416 23259 15419
rect 23308 15416 23336 15524
rect 23474 15512 23480 15524
rect 23532 15552 23538 15564
rect 24670 15552 24676 15564
rect 23532 15524 24676 15552
rect 23532 15512 23538 15524
rect 24670 15512 24676 15524
rect 24728 15552 24734 15564
rect 24728 15524 24808 15552
rect 24728 15512 24734 15524
rect 23382 15444 23388 15496
rect 23440 15484 23446 15496
rect 23440 15456 23533 15484
rect 23440 15444 23446 15456
rect 24394 15444 24400 15496
rect 24452 15484 24458 15496
rect 24780 15493 24808 15524
rect 26234 15512 26240 15564
rect 26292 15512 26298 15564
rect 28534 15512 28540 15564
rect 28592 15552 28598 15564
rect 32674 15552 32680 15564
rect 28592 15524 32680 15552
rect 28592 15512 28598 15524
rect 32674 15512 32680 15524
rect 32732 15512 32738 15564
rect 39868 15552 39896 15648
rect 40957 15623 41015 15629
rect 40957 15589 40969 15623
rect 41003 15620 41015 15623
rect 46584 15620 46612 15651
rect 52546 15648 52552 15660
rect 52604 15648 52610 15700
rect 52917 15691 52975 15697
rect 52917 15657 52929 15691
rect 52963 15657 52975 15691
rect 53098 15688 53104 15700
rect 53059 15660 53104 15688
rect 52917 15651 52975 15657
rect 50433 15623 50491 15629
rect 41003 15592 45554 15620
rect 46584 15592 46888 15620
rect 41003 15589 41015 15592
rect 40957 15583 41015 15589
rect 40497 15555 40555 15561
rect 40497 15552 40509 15555
rect 39868 15524 40509 15552
rect 40497 15521 40509 15524
rect 40543 15521 40555 15555
rect 45526 15552 45554 15592
rect 45526 15524 46796 15552
rect 40497 15515 40555 15521
rect 24581 15487 24639 15493
rect 24581 15484 24593 15487
rect 24452 15456 24593 15484
rect 24452 15444 24458 15456
rect 24581 15453 24593 15456
rect 24627 15453 24639 15487
rect 24581 15447 24639 15453
rect 24765 15487 24823 15493
rect 24765 15453 24777 15487
rect 24811 15453 24823 15487
rect 24765 15447 24823 15453
rect 24949 15487 25007 15493
rect 24949 15453 24961 15487
rect 24995 15484 25007 15487
rect 25222 15484 25228 15496
rect 24995 15456 25228 15484
rect 24995 15453 25007 15456
rect 24949 15447 25007 15453
rect 25222 15444 25228 15456
rect 25280 15444 25286 15496
rect 26053 15487 26111 15493
rect 26053 15453 26065 15487
rect 26099 15484 26111 15487
rect 26252 15484 26280 15512
rect 32125 15487 32183 15493
rect 32125 15484 32137 15487
rect 26099 15456 26280 15484
rect 31588 15456 32137 15484
rect 26099 15453 26111 15456
rect 26053 15447 26111 15453
rect 23247 15388 23336 15416
rect 23247 15385 23259 15388
rect 23201 15379 23259 15385
rect 3786 15308 3792 15360
rect 3844 15348 3850 15360
rect 3881 15351 3939 15357
rect 3881 15348 3893 15351
rect 3844 15320 3893 15348
rect 3844 15308 3850 15320
rect 3881 15317 3893 15320
rect 3927 15317 3939 15351
rect 8938 15348 8944 15360
rect 8899 15320 8944 15348
rect 3881 15311 3939 15317
rect 8938 15308 8944 15320
rect 8996 15308 9002 15360
rect 10686 15348 10692 15360
rect 10647 15320 10692 15348
rect 10686 15308 10692 15320
rect 10744 15308 10750 15360
rect 14274 15308 14280 15360
rect 14332 15348 14338 15360
rect 15838 15348 15844 15360
rect 14332 15320 15844 15348
rect 14332 15308 14338 15320
rect 15838 15308 15844 15320
rect 15896 15308 15902 15360
rect 17037 15351 17095 15357
rect 17037 15317 17049 15351
rect 17083 15348 17095 15351
rect 17586 15348 17592 15360
rect 17083 15320 17592 15348
rect 17083 15317 17095 15320
rect 17037 15311 17095 15317
rect 17586 15308 17592 15320
rect 17644 15308 17650 15360
rect 20254 15308 20260 15360
rect 20312 15348 20318 15360
rect 20349 15351 20407 15357
rect 20349 15348 20361 15351
rect 20312 15320 20361 15348
rect 20312 15308 20318 15320
rect 20349 15317 20361 15320
rect 20395 15317 20407 15351
rect 20349 15311 20407 15317
rect 21269 15351 21327 15357
rect 21269 15317 21281 15351
rect 21315 15348 21327 15351
rect 21910 15348 21916 15360
rect 21315 15320 21916 15348
rect 21315 15317 21327 15320
rect 21269 15311 21327 15317
rect 21910 15308 21916 15320
rect 21968 15308 21974 15360
rect 22278 15308 22284 15360
rect 22336 15348 22342 15360
rect 23400 15348 23428 15444
rect 24673 15419 24731 15425
rect 24673 15385 24685 15419
rect 24719 15416 24731 15419
rect 24854 15416 24860 15428
rect 24719 15388 24860 15416
rect 24719 15385 24731 15388
rect 24673 15379 24731 15385
rect 24854 15376 24860 15388
rect 24912 15376 24918 15428
rect 26237 15419 26295 15425
rect 26237 15385 26249 15419
rect 26283 15416 26295 15419
rect 26878 15416 26884 15428
rect 26283 15388 26884 15416
rect 26283 15385 26295 15388
rect 26237 15379 26295 15385
rect 26878 15376 26884 15388
rect 26936 15376 26942 15428
rect 25866 15348 25872 15360
rect 22336 15320 23428 15348
rect 25827 15320 25872 15348
rect 22336 15308 22342 15320
rect 25866 15308 25872 15320
rect 25924 15308 25930 15360
rect 31386 15308 31392 15360
rect 31444 15348 31450 15360
rect 31588 15357 31616 15456
rect 32125 15453 32137 15456
rect 32171 15484 32183 15487
rect 32306 15484 32312 15496
rect 32171 15456 32312 15484
rect 32171 15453 32183 15456
rect 32125 15447 32183 15453
rect 32306 15444 32312 15456
rect 32364 15444 32370 15496
rect 32493 15487 32551 15493
rect 32493 15453 32505 15487
rect 32539 15484 32551 15487
rect 33134 15484 33140 15496
rect 32539 15456 33140 15484
rect 32539 15453 32551 15456
rect 32493 15447 32551 15453
rect 33134 15444 33140 15456
rect 33192 15444 33198 15496
rect 40586 15484 40592 15496
rect 40547 15456 40592 15484
rect 40586 15444 40592 15456
rect 40644 15444 40650 15496
rect 41966 15484 41972 15496
rect 41927 15456 41972 15484
rect 41966 15444 41972 15456
rect 42024 15444 42030 15496
rect 42518 15484 42524 15496
rect 42479 15456 42524 15484
rect 42518 15444 42524 15456
rect 42576 15444 42582 15496
rect 42794 15484 42800 15496
rect 42755 15456 42800 15484
rect 42794 15444 42800 15456
rect 42852 15444 42858 15496
rect 46293 15487 46351 15493
rect 46293 15484 46305 15487
rect 45526 15456 46305 15484
rect 34057 15419 34115 15425
rect 34057 15416 34069 15419
rect 33336 15388 34069 15416
rect 33336 15360 33364 15388
rect 34057 15385 34069 15388
rect 34103 15385 34115 15419
rect 41984 15416 42012 15444
rect 42613 15419 42671 15425
rect 42613 15416 42625 15419
rect 41984 15388 42625 15416
rect 34057 15379 34115 15385
rect 42613 15385 42625 15388
rect 42659 15385 42671 15419
rect 43898 15416 43904 15428
rect 43859 15388 43904 15416
rect 42613 15379 42671 15385
rect 43898 15376 43904 15388
rect 43956 15376 43962 15428
rect 44450 15416 44456 15428
rect 44192 15388 44456 15416
rect 31573 15351 31631 15357
rect 31573 15348 31585 15351
rect 31444 15320 31585 15348
rect 31444 15308 31450 15320
rect 31573 15317 31585 15320
rect 31619 15317 31631 15351
rect 32122 15348 32128 15360
rect 32083 15320 32128 15348
rect 31573 15311 31631 15317
rect 32122 15308 32128 15320
rect 32180 15308 32186 15360
rect 32214 15308 32220 15360
rect 32272 15348 32278 15360
rect 32309 15351 32367 15357
rect 32309 15348 32321 15351
rect 32272 15320 32321 15348
rect 32272 15308 32278 15320
rect 32309 15317 32321 15320
rect 32355 15317 32367 15351
rect 32309 15311 32367 15317
rect 32398 15308 32404 15360
rect 32456 15348 32462 15360
rect 32953 15351 33011 15357
rect 32953 15348 32965 15351
rect 32456 15320 32965 15348
rect 32456 15308 32462 15320
rect 32953 15317 32965 15320
rect 32999 15348 33011 15351
rect 33318 15348 33324 15360
rect 32999 15320 33324 15348
rect 32999 15317 33011 15320
rect 32953 15311 33011 15317
rect 33318 15308 33324 15320
rect 33376 15308 33382 15360
rect 33502 15348 33508 15360
rect 33463 15320 33508 15348
rect 33502 15308 33508 15320
rect 33560 15308 33566 15360
rect 42981 15351 43039 15357
rect 42981 15317 42993 15351
rect 43027 15348 43039 15351
rect 44101 15351 44159 15357
rect 44101 15348 44113 15351
rect 43027 15320 44113 15348
rect 43027 15317 43039 15320
rect 42981 15311 43039 15317
rect 44101 15317 44113 15320
rect 44147 15348 44159 15351
rect 44192 15348 44220 15388
rect 44450 15376 44456 15388
rect 44508 15376 44514 15428
rect 44147 15320 44220 15348
rect 44269 15351 44327 15357
rect 44147 15317 44159 15320
rect 44101 15311 44159 15317
rect 44269 15317 44281 15351
rect 44315 15348 44327 15351
rect 45278 15348 45284 15360
rect 44315 15320 45284 15348
rect 44315 15317 44327 15320
rect 44269 15311 44327 15317
rect 45278 15308 45284 15320
rect 45336 15348 45342 15360
rect 45526 15348 45554 15456
rect 46293 15453 46305 15456
rect 46339 15453 46351 15487
rect 46293 15447 46351 15453
rect 46768 15416 46796 15524
rect 46860 15496 46888 15592
rect 50433 15589 50445 15623
rect 50479 15620 50491 15623
rect 52270 15620 52276 15632
rect 50479 15592 52276 15620
rect 50479 15589 50491 15592
rect 50433 15583 50491 15589
rect 52270 15580 52276 15592
rect 52328 15580 52334 15632
rect 52932 15620 52960 15651
rect 53098 15648 53104 15660
rect 53156 15648 53162 15700
rect 53006 15620 53012 15632
rect 52932 15592 53012 15620
rect 53006 15580 53012 15592
rect 53064 15580 53070 15632
rect 47302 15552 47308 15564
rect 47263 15524 47308 15552
rect 47302 15512 47308 15524
rect 47360 15512 47366 15564
rect 47765 15555 47823 15561
rect 47765 15521 47777 15555
rect 47811 15552 47823 15555
rect 52822 15552 52828 15564
rect 47811 15524 52828 15552
rect 47811 15521 47823 15524
rect 47765 15515 47823 15521
rect 46842 15444 46848 15496
rect 46900 15484 46906 15496
rect 47397 15487 47455 15493
rect 47397 15484 47409 15487
rect 46900 15456 47409 15484
rect 46900 15444 46906 15456
rect 47397 15453 47409 15456
rect 47443 15453 47455 15487
rect 49970 15484 49976 15496
rect 47397 15447 47455 15453
rect 49620 15456 49976 15484
rect 49620 15416 49648 15456
rect 49970 15444 49976 15456
rect 50028 15444 50034 15496
rect 50062 15444 50068 15496
rect 50120 15484 50126 15496
rect 52748 15493 52776 15524
rect 52822 15512 52828 15524
rect 52880 15512 52886 15564
rect 53558 15552 53564 15564
rect 53519 15524 53564 15552
rect 53558 15512 53564 15524
rect 53616 15512 53622 15564
rect 56778 15552 56784 15564
rect 56739 15524 56784 15552
rect 56778 15512 56784 15524
rect 56836 15512 56842 15564
rect 57701 15555 57759 15561
rect 57701 15521 57713 15555
rect 57747 15552 57759 15555
rect 57882 15552 57888 15564
rect 57747 15524 57888 15552
rect 57747 15521 57759 15524
rect 57701 15515 57759 15521
rect 57882 15512 57888 15524
rect 57940 15512 57946 15564
rect 50157 15487 50215 15493
rect 50157 15484 50169 15487
rect 50120 15456 50169 15484
rect 50120 15444 50126 15456
rect 50157 15453 50169 15456
rect 50203 15453 50215 15487
rect 50157 15447 50215 15453
rect 52733 15487 52791 15493
rect 52733 15453 52745 15487
rect 52779 15453 52791 15487
rect 52914 15484 52920 15496
rect 52875 15456 52920 15484
rect 52733 15447 52791 15453
rect 52914 15444 52920 15456
rect 52972 15444 52978 15496
rect 57054 15484 57060 15496
rect 57015 15456 57060 15484
rect 57054 15444 57060 15456
rect 57112 15444 57118 15496
rect 50433 15419 50491 15425
rect 50433 15416 50445 15419
rect 46768 15388 49648 15416
rect 49712 15388 50445 15416
rect 49712 15360 49740 15388
rect 50433 15385 50445 15388
rect 50479 15385 50491 15419
rect 50433 15379 50491 15385
rect 45336 15320 45554 15348
rect 45336 15308 45342 15320
rect 48682 15308 48688 15360
rect 48740 15348 48746 15360
rect 49694 15348 49700 15360
rect 48740 15320 49700 15348
rect 48740 15308 48746 15320
rect 49694 15308 49700 15320
rect 49752 15308 49758 15360
rect 50154 15308 50160 15360
rect 50212 15348 50218 15360
rect 50249 15351 50307 15357
rect 50249 15348 50261 15351
rect 50212 15320 50261 15348
rect 50212 15308 50218 15320
rect 50249 15317 50261 15320
rect 50295 15317 50307 15351
rect 50249 15311 50307 15317
rect 1104 15258 58880 15280
rect 1104 15206 19574 15258
rect 19626 15206 19638 15258
rect 19690 15206 19702 15258
rect 19754 15206 19766 15258
rect 19818 15206 19830 15258
rect 19882 15206 50294 15258
rect 50346 15206 50358 15258
rect 50410 15206 50422 15258
rect 50474 15206 50486 15258
rect 50538 15206 50550 15258
rect 50602 15206 58880 15258
rect 1104 15184 58880 15206
rect 2593 15147 2651 15153
rect 2593 15113 2605 15147
rect 2639 15144 2651 15147
rect 7561 15147 7619 15153
rect 2639 15116 4016 15144
rect 2639 15113 2651 15116
rect 2593 15107 2651 15113
rect 2133 15079 2191 15085
rect 2133 15045 2145 15079
rect 2179 15076 2191 15079
rect 2682 15076 2688 15088
rect 2179 15048 2688 15076
rect 2179 15045 2191 15048
rect 2133 15039 2191 15045
rect 2682 15036 2688 15048
rect 2740 15076 2746 15088
rect 2869 15079 2927 15085
rect 2869 15076 2881 15079
rect 2740 15048 2881 15076
rect 2740 15036 2746 15048
rect 2869 15045 2881 15048
rect 2915 15045 2927 15079
rect 2869 15039 2927 15045
rect 2961 15079 3019 15085
rect 2961 15045 2973 15079
rect 3007 15076 3019 15079
rect 3510 15076 3516 15088
rect 3007 15048 3516 15076
rect 3007 15045 3019 15048
rect 2961 15039 3019 15045
rect 3510 15036 3516 15048
rect 3568 15036 3574 15088
rect 3786 15076 3792 15088
rect 3747 15048 3792 15076
rect 3786 15036 3792 15048
rect 3844 15036 3850 15088
rect 2774 14968 2780 15020
rect 2832 15008 2838 15020
rect 3145 15011 3203 15017
rect 2832 14980 2877 15008
rect 2832 14968 2838 14980
rect 3145 14977 3157 15011
rect 3191 15008 3203 15011
rect 3191 14980 3372 15008
rect 3191 14977 3203 14980
rect 3145 14971 3203 14977
rect 3344 14804 3372 14980
rect 3418 14968 3424 15020
rect 3476 15008 3482 15020
rect 3605 15011 3663 15017
rect 3605 15008 3617 15011
rect 3476 14980 3617 15008
rect 3476 14968 3482 14980
rect 3605 14977 3617 14980
rect 3651 14977 3663 15011
rect 3878 15008 3884 15020
rect 3839 14980 3884 15008
rect 3605 14971 3663 14977
rect 3878 14968 3884 14980
rect 3936 14968 3942 15020
rect 3988 15017 4016 15116
rect 7561 15113 7573 15147
rect 7607 15144 7619 15147
rect 7742 15144 7748 15156
rect 7607 15116 7748 15144
rect 7607 15113 7619 15116
rect 7561 15107 7619 15113
rect 7742 15104 7748 15116
rect 7800 15104 7806 15156
rect 9214 15144 9220 15156
rect 9175 15116 9220 15144
rect 9214 15104 9220 15116
rect 9272 15104 9278 15156
rect 10873 15147 10931 15153
rect 10873 15113 10885 15147
rect 10919 15144 10931 15147
rect 12342 15144 12348 15156
rect 10919 15116 12348 15144
rect 10919 15113 10931 15116
rect 10873 15107 10931 15113
rect 12342 15104 12348 15116
rect 12400 15104 12406 15156
rect 14182 15104 14188 15156
rect 14240 15144 14246 15156
rect 14619 15147 14677 15153
rect 14619 15144 14631 15147
rect 14240 15116 14631 15144
rect 14240 15104 14246 15116
rect 14619 15113 14631 15116
rect 14665 15113 14677 15147
rect 19334 15144 19340 15156
rect 14619 15107 14677 15113
rect 14752 15116 19340 15144
rect 6638 15036 6644 15088
rect 6696 15076 6702 15088
rect 10042 15076 10048 15088
rect 6696 15048 7696 15076
rect 10003 15048 10048 15076
rect 6696 15036 6702 15048
rect 3978 15011 4036 15017
rect 3978 14977 3990 15011
rect 4024 14977 4036 15011
rect 5810 15008 5816 15020
rect 5723 14980 5816 15008
rect 3978 14971 4036 14977
rect 5810 14968 5816 14980
rect 5868 15008 5874 15020
rect 6549 15011 6607 15017
rect 6549 15008 6561 15011
rect 5868 14980 6561 15008
rect 5868 14968 5874 14980
rect 6549 14977 6561 14980
rect 6595 14977 6607 15011
rect 7190 15008 7196 15020
rect 6549 14971 6607 14977
rect 6932 14980 7196 15008
rect 4157 14875 4215 14881
rect 4157 14841 4169 14875
rect 4203 14872 4215 14875
rect 4982 14872 4988 14884
rect 4203 14844 4988 14872
rect 4203 14841 4215 14844
rect 4157 14835 4215 14841
rect 4982 14832 4988 14844
rect 5040 14832 5046 14884
rect 4706 14804 4712 14816
rect 3344 14776 4712 14804
rect 4706 14764 4712 14776
rect 4764 14764 4770 14816
rect 6564 14804 6592 14971
rect 6932 14949 6960 14980
rect 7190 14968 7196 14980
rect 7248 15008 7254 15020
rect 7668 15017 7696 15048
rect 10042 15036 10048 15048
rect 10100 15036 10106 15088
rect 11517 15079 11575 15085
rect 11517 15045 11529 15079
rect 11563 15045 11575 15079
rect 11733 15079 11791 15085
rect 11733 15076 11745 15079
rect 11517 15039 11575 15045
rect 11624 15048 11745 15076
rect 7377 15011 7435 15017
rect 7377 15008 7389 15011
rect 7248 14980 7389 15008
rect 7248 14968 7254 14980
rect 7377 14977 7389 14980
rect 7423 14977 7435 15011
rect 7377 14971 7435 14977
rect 7653 15011 7711 15017
rect 7653 14977 7665 15011
rect 7699 14977 7711 15011
rect 7653 14971 7711 14977
rect 7837 15011 7895 15017
rect 7837 14977 7849 15011
rect 7883 15008 7895 15011
rect 9217 15011 9275 15017
rect 7883 14980 8432 15008
rect 7883 14977 7895 14980
rect 7837 14971 7895 14977
rect 6641 14943 6699 14949
rect 6641 14909 6653 14943
rect 6687 14909 6699 14943
rect 6641 14903 6699 14909
rect 6917 14943 6975 14949
rect 6917 14909 6929 14943
rect 6963 14909 6975 14943
rect 6917 14903 6975 14909
rect 6656 14872 6684 14903
rect 7852 14872 7880 14971
rect 8404 14881 8432 14980
rect 9217 14977 9229 15011
rect 9263 14977 9275 15011
rect 9217 14971 9275 14977
rect 9401 15011 9459 15017
rect 9401 14977 9413 15011
rect 9447 15008 9459 15011
rect 9861 15011 9919 15017
rect 9861 15008 9873 15011
rect 9447 14980 9873 15008
rect 9447 14977 9459 14980
rect 9401 14971 9459 14977
rect 9861 14977 9873 14980
rect 9907 14977 9919 15011
rect 9861 14971 9919 14977
rect 9232 14940 9260 14971
rect 10134 14968 10140 15020
rect 10192 15008 10198 15020
rect 10229 15011 10287 15017
rect 10229 15008 10241 15011
rect 10192 14980 10241 15008
rect 10192 14968 10198 14980
rect 10229 14977 10241 14980
rect 10275 14977 10287 15011
rect 10686 15008 10692 15020
rect 10599 14980 10692 15008
rect 10229 14971 10287 14977
rect 10686 14968 10692 14980
rect 10744 15008 10750 15020
rect 11532 15008 11560 15039
rect 10744 14980 11560 15008
rect 10744 14968 10750 14980
rect 10704 14940 10732 14968
rect 9232 14912 10732 14940
rect 6656 14844 7880 14872
rect 8389 14875 8447 14881
rect 8389 14841 8401 14875
rect 8435 14872 8447 14875
rect 8938 14872 8944 14884
rect 8435 14844 8944 14872
rect 8435 14841 8447 14844
rect 8389 14835 8447 14841
rect 8938 14832 8944 14844
rect 8996 14832 9002 14884
rect 10410 14832 10416 14884
rect 10468 14872 10474 14884
rect 11624 14872 11652 15048
rect 11733 15045 11745 15048
rect 11779 15076 11791 15079
rect 12066 15076 12072 15088
rect 11779 15048 12072 15076
rect 11779 15045 11791 15048
rect 11733 15039 11791 15045
rect 12066 15036 12072 15048
rect 12124 15036 12130 15088
rect 14752 15076 14780 15116
rect 19334 15104 19340 15116
rect 19392 15104 19398 15156
rect 20530 15144 20536 15156
rect 20272 15116 20536 15144
rect 12452 15048 14780 15076
rect 14829 15079 14887 15085
rect 12452 15020 12480 15048
rect 14829 15045 14841 15079
rect 14875 15076 14887 15079
rect 15010 15076 15016 15088
rect 14875 15048 15016 15076
rect 14875 15045 14887 15048
rect 14829 15039 14887 15045
rect 15010 15036 15016 15048
rect 15068 15036 15074 15088
rect 15749 15079 15807 15085
rect 15749 15076 15761 15079
rect 15672 15048 15761 15076
rect 11882 14968 11888 15020
rect 11940 15008 11946 15020
rect 12345 15011 12403 15017
rect 12345 15008 12357 15011
rect 11940 14980 12357 15008
rect 11940 14968 11946 14980
rect 12345 14977 12357 14980
rect 12391 14977 12403 15011
rect 12345 14971 12403 14977
rect 12434 14968 12440 15020
rect 12492 15008 12498 15020
rect 12492 14980 12585 15008
rect 12492 14968 12498 14980
rect 12618 14968 12624 15020
rect 12676 15008 12682 15020
rect 13265 15011 13323 15017
rect 12676 14980 12721 15008
rect 12676 14968 12682 14980
rect 13265 14977 13277 15011
rect 13311 14977 13323 15011
rect 13265 14971 13323 14977
rect 13280 14940 13308 14971
rect 13446 14968 13452 15020
rect 13504 15008 13510 15020
rect 13541 15011 13599 15017
rect 13541 15008 13553 15011
rect 13504 14980 13553 15008
rect 13504 14968 13510 14980
rect 13541 14977 13553 14980
rect 13587 14977 13599 15011
rect 13541 14971 13599 14977
rect 14001 15011 14059 15017
rect 14001 14977 14013 15011
rect 14047 15008 14059 15011
rect 15194 15008 15200 15020
rect 14047 14980 15200 15008
rect 14047 14977 14059 14980
rect 14001 14971 14059 14977
rect 15194 14968 15200 14980
rect 15252 14968 15258 15020
rect 15562 15008 15568 15020
rect 15523 14980 15568 15008
rect 15562 14968 15568 14980
rect 15620 14968 15626 15020
rect 12636 14912 13308 14940
rect 10468 14844 11652 14872
rect 10468 14832 10474 14844
rect 12526 14832 12532 14884
rect 12584 14872 12590 14884
rect 12636 14881 12664 14912
rect 15470 14900 15476 14952
rect 15528 14940 15534 14952
rect 15672 14940 15700 15048
rect 15749 15045 15761 15048
rect 15795 15045 15807 15079
rect 15749 15039 15807 15045
rect 15838 15036 15844 15088
rect 15896 15076 15902 15088
rect 17954 15076 17960 15088
rect 15896 15048 15941 15076
rect 17144 15048 17960 15076
rect 15896 15036 15902 15048
rect 17144 15017 17172 15048
rect 17954 15036 17960 15048
rect 18012 15036 18018 15088
rect 15957 15011 16015 15017
rect 15957 15008 15969 15011
rect 15948 14977 15969 15008
rect 16003 14977 16015 15011
rect 15948 14971 16015 14977
rect 17129 15011 17187 15017
rect 17129 14977 17141 15011
rect 17175 14977 17187 15011
rect 17586 15008 17592 15020
rect 17547 14980 17592 15008
rect 17129 14971 17187 14977
rect 15948 14940 15976 14971
rect 17586 14968 17592 14980
rect 17644 14968 17650 15020
rect 20070 15008 20076 15020
rect 20031 14980 20076 15008
rect 20070 14968 20076 14980
rect 20128 14968 20134 15020
rect 20166 15011 20224 15017
rect 20166 14977 20178 15011
rect 20212 15008 20224 15011
rect 20272 15008 20300 15116
rect 20530 15104 20536 15116
rect 20588 15104 20594 15156
rect 20714 15144 20720 15156
rect 20675 15116 20720 15144
rect 20714 15104 20720 15116
rect 20772 15104 20778 15156
rect 23566 15104 23572 15156
rect 23624 15144 23630 15156
rect 24210 15144 24216 15156
rect 23624 15116 24216 15144
rect 23624 15104 23630 15116
rect 24210 15104 24216 15116
rect 24268 15144 24274 15156
rect 24268 15116 24532 15144
rect 24268 15104 24274 15116
rect 20349 15079 20407 15085
rect 20349 15045 20361 15079
rect 20395 15076 20407 15079
rect 20990 15076 20996 15088
rect 20395 15048 20996 15076
rect 20395 15045 20407 15048
rect 20349 15039 20407 15045
rect 20990 15036 20996 15048
rect 21048 15036 21054 15088
rect 22094 15036 22100 15088
rect 22152 15076 22158 15088
rect 23106 15076 23112 15088
rect 22152 15048 23112 15076
rect 22152 15036 22158 15048
rect 23106 15036 23112 15048
rect 23164 15076 23170 15088
rect 24504 15085 24532 15116
rect 27614 15104 27620 15156
rect 27672 15144 27678 15156
rect 28810 15144 28816 15156
rect 27672 15116 28816 15144
rect 27672 15104 27678 15116
rect 28810 15104 28816 15116
rect 28868 15144 28874 15156
rect 29917 15147 29975 15153
rect 28868 15116 28948 15144
rect 28868 15104 28874 15116
rect 24397 15079 24455 15085
rect 24397 15076 24409 15079
rect 23164 15048 24409 15076
rect 23164 15036 23170 15048
rect 24397 15045 24409 15048
rect 24443 15045 24455 15079
rect 24397 15039 24455 15045
rect 24489 15079 24547 15085
rect 24489 15045 24501 15079
rect 24535 15045 24547 15079
rect 25038 15076 25044 15088
rect 24489 15039 24547 15045
rect 24688 15048 25044 15076
rect 20441 15011 20499 15017
rect 20441 15008 20453 15011
rect 20212 14980 20300 15008
rect 20364 14980 20453 15008
rect 20212 14977 20224 14980
rect 20166 14971 20224 14977
rect 15528 14912 15700 14940
rect 15856 14912 15976 14940
rect 16761 14943 16819 14949
rect 15528 14900 15534 14912
rect 15856 14884 15884 14912
rect 16761 14909 16773 14943
rect 16807 14909 16819 14943
rect 16761 14903 16819 14909
rect 12621 14875 12679 14881
rect 12621 14872 12633 14875
rect 12584 14844 12633 14872
rect 12584 14832 12590 14844
rect 12621 14841 12633 14844
rect 12667 14841 12679 14875
rect 13354 14872 13360 14884
rect 13315 14844 13360 14872
rect 12621 14835 12679 14841
rect 13354 14832 13360 14844
rect 13412 14832 13418 14884
rect 14458 14872 14464 14884
rect 14419 14844 14464 14872
rect 14458 14832 14464 14844
rect 14516 14832 14522 14884
rect 15838 14832 15844 14884
rect 15896 14832 15902 14884
rect 15930 14832 15936 14884
rect 15988 14872 15994 14884
rect 16776 14872 16804 14903
rect 16850 14900 16856 14952
rect 16908 14940 16914 14952
rect 17402 14940 17408 14952
rect 16908 14912 17408 14940
rect 16908 14900 16914 14912
rect 17402 14900 17408 14912
rect 17460 14940 17466 14952
rect 20181 14940 20209 14971
rect 20364 14952 20392 14980
rect 20441 14977 20453 14980
rect 20487 14977 20499 15011
rect 20441 14971 20499 14977
rect 20530 14968 20536 15020
rect 20588 15017 20594 15020
rect 20588 15011 20615 15017
rect 20603 14977 20615 15011
rect 20588 14971 20615 14977
rect 20588 14968 20594 14971
rect 23290 14968 23296 15020
rect 23348 15008 23354 15020
rect 24688 15017 24716 15048
rect 25038 15036 25044 15048
rect 25096 15036 25102 15088
rect 26234 15036 26240 15088
rect 26292 15076 26298 15088
rect 26292 15048 27200 15076
rect 26292 15036 26298 15048
rect 24300 15011 24358 15017
rect 24300 15008 24312 15011
rect 23348 14980 24312 15008
rect 23348 14968 23354 14980
rect 24300 14977 24312 14980
rect 24346 14977 24358 15011
rect 24300 14971 24358 14977
rect 24672 15011 24730 15017
rect 24672 14977 24684 15011
rect 24718 14977 24730 15011
rect 24672 14971 24730 14977
rect 17460 14912 20209 14940
rect 17460 14900 17466 14912
rect 20346 14900 20352 14952
rect 20404 14900 20410 14952
rect 24315 14940 24343 14971
rect 24762 14968 24768 15020
rect 24820 15008 24826 15020
rect 25866 15008 25872 15020
rect 24820 14980 24865 15008
rect 25827 14980 25872 15008
rect 24820 14968 24826 14980
rect 25866 14968 25872 14980
rect 25924 14968 25930 15020
rect 26145 15011 26203 15017
rect 26145 14977 26157 15011
rect 26191 14977 26203 15011
rect 26145 14971 26203 14977
rect 25590 14940 25596 14952
rect 24315 14912 25596 14940
rect 25590 14900 25596 14912
rect 25648 14900 25654 14952
rect 26160 14940 26188 14971
rect 26878 14968 26884 15020
rect 26936 15008 26942 15020
rect 27172 15017 27200 15048
rect 28074 15036 28080 15088
rect 28132 15076 28138 15088
rect 28721 15079 28779 15085
rect 28721 15076 28733 15079
rect 28132 15048 28733 15076
rect 28132 15036 28138 15048
rect 28721 15045 28733 15048
rect 28767 15045 28779 15079
rect 28721 15039 28779 15045
rect 28920 15076 28948 15116
rect 29917 15113 29929 15147
rect 29963 15144 29975 15147
rect 38378 15144 38384 15156
rect 29963 15116 37504 15144
rect 38339 15116 38384 15144
rect 29963 15113 29975 15116
rect 29917 15107 29975 15113
rect 30926 15076 30932 15088
rect 28920 15048 30788 15076
rect 30887 15048 30932 15076
rect 26973 15011 27031 15017
rect 26973 15008 26985 15011
rect 26936 14980 26985 15008
rect 26936 14968 26942 14980
rect 26973 14977 26985 14980
rect 27019 14977 27031 15011
rect 26973 14971 27031 14977
rect 27157 15011 27215 15017
rect 27157 14977 27169 15011
rect 27203 15008 27215 15011
rect 27617 15011 27675 15017
rect 27617 15008 27629 15011
rect 27203 14980 27629 15008
rect 27203 14977 27215 14980
rect 27157 14971 27215 14977
rect 27617 14977 27629 14980
rect 27663 14977 27675 15011
rect 27617 14971 27675 14977
rect 28537 15011 28595 15017
rect 28537 14977 28549 15011
rect 28583 14977 28595 15011
rect 28537 14971 28595 14977
rect 28552 14940 28580 14971
rect 28626 14968 28632 15020
rect 28684 15008 28690 15020
rect 28920 15017 28948 15048
rect 28813 15011 28871 15017
rect 28813 15008 28825 15011
rect 28684 14980 28825 15008
rect 28684 14968 28690 14980
rect 28813 14977 28825 14980
rect 28859 14977 28871 15011
rect 28813 14971 28871 14977
rect 28905 15011 28963 15017
rect 28905 14977 28917 15011
rect 28951 14977 28963 15011
rect 28905 14971 28963 14977
rect 29917 15011 29975 15017
rect 29917 14977 29929 15011
rect 29963 15008 29975 15011
rect 30006 15008 30012 15020
rect 29963 14980 30012 15008
rect 29963 14977 29975 14980
rect 29917 14971 29975 14977
rect 30006 14968 30012 14980
rect 30064 14968 30070 15020
rect 30760 15017 30788 15048
rect 30926 15036 30932 15048
rect 30984 15036 30990 15088
rect 32214 15076 32220 15088
rect 31312 15048 32220 15076
rect 30745 15011 30803 15017
rect 30745 14977 30757 15011
rect 30791 14977 30803 15011
rect 30745 14971 30803 14977
rect 30834 14968 30840 15020
rect 30892 15008 30898 15020
rect 31110 15008 31116 15020
rect 30892 14980 30937 15008
rect 31071 14980 31116 15008
rect 30892 14968 30898 14980
rect 31110 14968 31116 14980
rect 31168 14968 31174 15020
rect 28994 14940 29000 14952
rect 26160 14912 27108 14940
rect 28552 14912 29000 14940
rect 17678 14872 17684 14884
rect 15988 14844 16804 14872
rect 17639 14844 17684 14872
rect 15988 14832 15994 14844
rect 17678 14832 17684 14844
rect 17736 14832 17742 14884
rect 19518 14872 19524 14884
rect 19431 14844 19524 14872
rect 19518 14832 19524 14844
rect 19576 14872 19582 14884
rect 20364 14872 20392 14900
rect 19576 14844 20392 14872
rect 19576 14832 19582 14844
rect 20714 14832 20720 14884
rect 20772 14872 20778 14884
rect 27080 14881 27108 14912
rect 28994 14900 29000 14912
rect 29052 14900 29058 14952
rect 29549 14943 29607 14949
rect 29549 14909 29561 14943
rect 29595 14909 29607 14943
rect 29549 14903 29607 14909
rect 25961 14875 26019 14881
rect 25961 14872 25973 14875
rect 20772 14844 25973 14872
rect 20772 14832 20778 14844
rect 25961 14841 25973 14844
rect 26007 14841 26019 14875
rect 25961 14835 26019 14841
rect 27065 14875 27123 14881
rect 27065 14841 27077 14875
rect 27111 14872 27123 14875
rect 29089 14875 29147 14881
rect 27111 14844 28304 14872
rect 27111 14841 27123 14844
rect 27065 14835 27123 14841
rect 10594 14804 10600 14816
rect 6564 14776 10600 14804
rect 10594 14764 10600 14776
rect 10652 14764 10658 14816
rect 10962 14764 10968 14816
rect 11020 14804 11026 14816
rect 11701 14807 11759 14813
rect 11701 14804 11713 14807
rect 11020 14776 11713 14804
rect 11020 14764 11026 14776
rect 11701 14773 11713 14776
rect 11747 14804 11759 14807
rect 11790 14804 11796 14816
rect 11747 14776 11796 14804
rect 11747 14773 11759 14776
rect 11701 14767 11759 14773
rect 11790 14764 11796 14776
rect 11848 14764 11854 14816
rect 11885 14807 11943 14813
rect 11885 14773 11897 14807
rect 11931 14804 11943 14807
rect 13372 14804 13400 14832
rect 14642 14804 14648 14816
rect 11931 14776 13400 14804
rect 14555 14776 14648 14804
rect 11931 14773 11943 14776
rect 11885 14767 11943 14773
rect 14642 14764 14648 14776
rect 14700 14804 14706 14816
rect 15286 14804 15292 14816
rect 14700 14776 15292 14804
rect 14700 14764 14706 14776
rect 15286 14764 15292 14776
rect 15344 14764 15350 14816
rect 16117 14807 16175 14813
rect 16117 14773 16129 14807
rect 16163 14804 16175 14807
rect 17218 14804 17224 14816
rect 16163 14776 17224 14804
rect 16163 14773 16175 14776
rect 16117 14767 16175 14773
rect 17218 14764 17224 14776
rect 17276 14764 17282 14816
rect 20162 14764 20168 14816
rect 20220 14804 20226 14816
rect 20530 14804 20536 14816
rect 20220 14776 20536 14804
rect 20220 14764 20226 14776
rect 20530 14764 20536 14776
rect 20588 14764 20594 14816
rect 23566 14804 23572 14816
rect 23527 14776 23572 14804
rect 23566 14764 23572 14776
rect 23624 14764 23630 14816
rect 24118 14804 24124 14816
rect 24079 14776 24124 14804
rect 24118 14764 24124 14776
rect 24176 14764 24182 14816
rect 28276 14804 28304 14844
rect 29089 14841 29101 14875
rect 29135 14872 29147 14875
rect 29564 14872 29592 14903
rect 30098 14900 30104 14952
rect 30156 14940 30162 14952
rect 31312 14940 31340 15048
rect 32214 15036 32220 15048
rect 32272 15076 32278 15088
rect 33134 15076 33140 15088
rect 32272 15048 32444 15076
rect 32272 15036 32278 15048
rect 32030 14968 32036 15020
rect 32088 15008 32094 15020
rect 32416 15017 32444 15048
rect 32600 15048 33140 15076
rect 32600 15017 32628 15048
rect 33134 15036 33140 15048
rect 33192 15076 33198 15088
rect 33192 15048 34376 15076
rect 33192 15036 33198 15048
rect 34348 15020 34376 15048
rect 37476 15020 37504 15116
rect 38378 15104 38384 15116
rect 38436 15144 38442 15156
rect 38933 15147 38991 15153
rect 38933 15144 38945 15147
rect 38436 15116 38945 15144
rect 38436 15104 38442 15116
rect 38933 15113 38945 15116
rect 38979 15113 38991 15147
rect 50154 15144 50160 15156
rect 38933 15107 38991 15113
rect 46400 15116 50160 15144
rect 32310 15011 32368 15017
rect 32088 15006 32168 15008
rect 32310 15006 32322 15011
rect 32088 14980 32322 15006
rect 32088 14968 32094 14980
rect 32140 14978 32322 14980
rect 32310 14977 32322 14978
rect 32356 14977 32368 15011
rect 32310 14971 32368 14977
rect 32401 15011 32459 15017
rect 32401 14977 32413 15011
rect 32447 14977 32459 15011
rect 32401 14971 32459 14977
rect 32585 15011 32643 15017
rect 32585 14977 32597 15011
rect 32631 14977 32643 15011
rect 33502 15008 33508 15020
rect 32585 14971 32643 14977
rect 32692 14980 33508 15008
rect 30156 14912 30201 14940
rect 30484 14912 31340 14940
rect 32493 14943 32551 14949
rect 30156 14900 30162 14912
rect 29135 14844 29592 14872
rect 29135 14841 29147 14844
rect 29089 14835 29147 14841
rect 30484 14804 30512 14912
rect 32493 14909 32505 14943
rect 32539 14940 32551 14943
rect 32692 14940 32720 14980
rect 33502 14968 33508 14980
rect 33560 14968 33566 15020
rect 34330 15008 34336 15020
rect 34291 14980 34336 15008
rect 34330 14968 34336 14980
rect 34388 14968 34394 15020
rect 37458 15008 37464 15020
rect 37371 14980 37464 15008
rect 37458 14968 37464 14980
rect 37516 14968 37522 15020
rect 37553 15011 37611 15017
rect 37553 14977 37565 15011
rect 37599 14977 37611 15011
rect 37553 14971 37611 14977
rect 37737 15011 37795 15017
rect 37737 14977 37749 15011
rect 37783 15008 37795 15011
rect 38396 15008 38424 15104
rect 43254 15036 43260 15088
rect 43312 15076 43318 15088
rect 44082 15076 44088 15088
rect 43312 15048 44088 15076
rect 43312 15036 43318 15048
rect 44082 15036 44088 15048
rect 44140 15076 44146 15088
rect 44140 15048 45508 15076
rect 44140 15036 44146 15048
rect 37783 14980 38424 15008
rect 37783 14977 37795 14980
rect 37737 14971 37795 14977
rect 33318 14940 33324 14952
rect 32539 14912 32720 14940
rect 33279 14912 33324 14940
rect 32539 14909 32551 14912
rect 32493 14903 32551 14909
rect 32306 14832 32312 14884
rect 32364 14872 32370 14884
rect 32508 14872 32536 14903
rect 33318 14900 33324 14912
rect 33376 14900 33382 14952
rect 33870 14940 33876 14952
rect 33831 14912 33876 14940
rect 33870 14900 33876 14912
rect 33928 14900 33934 14952
rect 37568 14940 37596 14971
rect 40586 14968 40592 15020
rect 40644 15008 40650 15020
rect 40957 15011 41015 15017
rect 40957 15008 40969 15011
rect 40644 14980 40969 15008
rect 40644 14968 40650 14980
rect 40957 14977 40969 14980
rect 41003 14977 41015 15011
rect 40957 14971 41015 14977
rect 44174 14968 44180 15020
rect 44232 15008 44238 15020
rect 44269 15011 44327 15017
rect 44269 15008 44281 15011
rect 44232 14980 44281 15008
rect 44232 14968 44238 14980
rect 44269 14977 44281 14980
rect 44315 14977 44327 15011
rect 44269 14971 44327 14977
rect 38010 14940 38016 14952
rect 37568 14912 38016 14940
rect 38010 14900 38016 14912
rect 38068 14900 38074 14952
rect 44284 14940 44312 14971
rect 44358 14968 44364 15020
rect 44416 15008 44422 15020
rect 44560 15017 44588 15048
rect 44545 15011 44603 15017
rect 44416 14980 44461 15008
rect 44416 14968 44422 14980
rect 44545 14977 44557 15011
rect 44591 14977 44603 15011
rect 45189 15011 45247 15017
rect 45189 15008 45201 15011
rect 44545 14971 44603 14977
rect 44652 14980 45201 15008
rect 44652 14940 44680 14980
rect 45189 14977 45201 14980
rect 45235 14977 45247 15011
rect 45370 15008 45376 15020
rect 45331 14980 45376 15008
rect 45189 14971 45247 14977
rect 45370 14968 45376 14980
rect 45428 14968 45434 15020
rect 45480 15017 45508 15048
rect 45465 15011 45523 15017
rect 45465 14977 45477 15011
rect 45511 14977 45523 15011
rect 45465 14971 45523 14977
rect 44284 14912 44680 14940
rect 44729 14943 44787 14949
rect 44729 14909 44741 14943
rect 44775 14940 44787 14943
rect 45922 14940 45928 14952
rect 44775 14912 45928 14940
rect 44775 14909 44787 14912
rect 44729 14903 44787 14909
rect 45922 14900 45928 14912
rect 45980 14940 45986 14952
rect 46293 14943 46351 14949
rect 46293 14940 46305 14943
rect 45980 14912 46305 14940
rect 45980 14900 45986 14912
rect 46293 14909 46305 14912
rect 46339 14909 46351 14943
rect 46293 14903 46351 14909
rect 33778 14872 33784 14884
rect 32364 14844 32536 14872
rect 33739 14844 33784 14872
rect 32364 14832 32370 14844
rect 33778 14832 33784 14844
rect 33836 14832 33842 14884
rect 37921 14875 37979 14881
rect 37921 14841 37933 14875
rect 37967 14872 37979 14875
rect 46400 14872 46428 15116
rect 46477 15011 46535 15017
rect 46477 14977 46489 15011
rect 46523 14977 46535 15011
rect 48682 15008 48688 15020
rect 48643 14980 48688 15008
rect 46477 14971 46535 14977
rect 37967 14844 46428 14872
rect 37967 14841 37979 14844
rect 37921 14835 37979 14841
rect 28276 14776 30512 14804
rect 30561 14807 30619 14813
rect 30561 14773 30573 14807
rect 30607 14804 30619 14807
rect 30834 14804 30840 14816
rect 30607 14776 30840 14804
rect 30607 14773 30619 14776
rect 30561 14767 30619 14773
rect 30834 14764 30840 14776
rect 30892 14764 30898 14816
rect 32030 14764 32036 14816
rect 32088 14804 32094 14816
rect 32125 14807 32183 14813
rect 32125 14804 32137 14807
rect 32088 14776 32137 14804
rect 32088 14764 32094 14776
rect 32125 14773 32137 14776
rect 32171 14773 32183 14807
rect 32125 14767 32183 14773
rect 34425 14807 34483 14813
rect 34425 14773 34437 14807
rect 34471 14804 34483 14807
rect 34514 14804 34520 14816
rect 34471 14776 34520 14804
rect 34471 14773 34483 14776
rect 34425 14767 34483 14773
rect 34514 14764 34520 14776
rect 34572 14764 34578 14816
rect 34606 14764 34612 14816
rect 34664 14804 34670 14816
rect 35069 14807 35127 14813
rect 35069 14804 35081 14807
rect 34664 14776 35081 14804
rect 34664 14764 34670 14776
rect 35069 14773 35081 14776
rect 35115 14804 35127 14807
rect 36354 14804 36360 14816
rect 35115 14776 36360 14804
rect 35115 14773 35127 14776
rect 35069 14767 35127 14773
rect 36354 14764 36360 14776
rect 36412 14764 36418 14816
rect 40770 14804 40776 14816
rect 40731 14776 40776 14804
rect 40770 14764 40776 14776
rect 40828 14764 40834 14816
rect 44358 14764 44364 14816
rect 44416 14804 44422 14816
rect 45370 14804 45376 14816
rect 44416 14776 45376 14804
rect 44416 14764 44422 14776
rect 45370 14764 45376 14776
rect 45428 14764 45434 14816
rect 45465 14807 45523 14813
rect 45465 14773 45477 14807
rect 45511 14804 45523 14807
rect 45830 14804 45836 14816
rect 45511 14776 45836 14804
rect 45511 14773 45523 14776
rect 45465 14767 45523 14773
rect 45830 14764 45836 14776
rect 45888 14804 45894 14816
rect 46492 14804 46520 14971
rect 48682 14968 48688 14980
rect 48740 14968 48746 15020
rect 48774 14968 48780 15020
rect 48832 15008 48838 15020
rect 48869 15011 48927 15017
rect 48869 15008 48881 15011
rect 48832 14980 48881 15008
rect 48832 14968 48838 14980
rect 48869 14977 48881 14980
rect 48915 14977 48927 15011
rect 48869 14971 48927 14977
rect 48961 15011 49019 15017
rect 48961 14977 48973 15011
rect 49007 15006 49019 15011
rect 49068 15006 49096 15116
rect 49528 15085 49556 15116
rect 50154 15104 50160 15116
rect 50212 15104 50218 15156
rect 50709 15147 50767 15153
rect 50709 15113 50721 15147
rect 50755 15113 50767 15147
rect 50709 15107 50767 15113
rect 49513 15079 49571 15085
rect 49513 15045 49525 15079
rect 49559 15045 49571 15079
rect 49513 15039 49571 15045
rect 49881 15079 49939 15085
rect 49881 15045 49893 15079
rect 49927 15076 49939 15079
rect 50246 15076 50252 15088
rect 49927 15048 50252 15076
rect 49927 15045 49939 15048
rect 49881 15039 49939 15045
rect 50246 15036 50252 15048
rect 50304 15076 50310 15088
rect 50341 15079 50399 15085
rect 50341 15076 50353 15079
rect 50304 15048 50353 15076
rect 50304 15036 50310 15048
rect 50341 15045 50353 15048
rect 50387 15045 50399 15079
rect 50541 15079 50599 15085
rect 50541 15076 50553 15079
rect 50341 15039 50399 15045
rect 50448 15048 50553 15076
rect 50448 15020 50476 15048
rect 50541 15045 50553 15048
rect 50587 15045 50599 15079
rect 50724 15076 50752 15107
rect 56686 15104 56692 15156
rect 56744 15144 56750 15156
rect 56873 15147 56931 15153
rect 56873 15144 56885 15147
rect 56744 15116 56885 15144
rect 56744 15104 56750 15116
rect 56873 15113 56885 15116
rect 56919 15144 56931 15147
rect 57422 15144 57428 15156
rect 56919 15116 57428 15144
rect 56919 15113 56931 15116
rect 56873 15107 56931 15113
rect 57422 15104 57428 15116
rect 57480 15104 57486 15156
rect 52914 15076 52920 15088
rect 50724 15048 52920 15076
rect 50541 15039 50599 15045
rect 52914 15036 52920 15048
rect 52972 15076 52978 15088
rect 52972 15048 53144 15076
rect 52972 15036 52978 15048
rect 49694 15008 49700 15020
rect 49007 14978 49096 15006
rect 49437 15001 49495 15007
rect 49007 14977 49019 14978
rect 48961 14971 49019 14977
rect 49437 14967 49449 15001
rect 49483 14998 49495 15001
rect 49483 14970 49556 14998
rect 49655 14980 49700 15008
rect 49483 14967 49495 14970
rect 49437 14961 49495 14967
rect 48774 14832 48780 14884
rect 48832 14872 48838 14884
rect 49528 14872 49556 14970
rect 49694 14968 49700 14980
rect 49752 14968 49758 15020
rect 49970 14968 49976 15020
rect 50028 15008 50034 15020
rect 50430 15008 50436 15020
rect 50028 14980 50436 15008
rect 50028 14968 50034 14980
rect 50430 14968 50436 14980
rect 50488 14968 50494 15020
rect 52546 14968 52552 15020
rect 52604 15008 52610 15020
rect 53116 15017 53144 15048
rect 53558 15036 53564 15088
rect 53616 15076 53622 15088
rect 54297 15079 54355 15085
rect 54297 15076 54309 15079
rect 53616 15048 54309 15076
rect 53616 15036 53622 15048
rect 54297 15045 54309 15048
rect 54343 15045 54355 15079
rect 54297 15039 54355 15045
rect 52825 15011 52883 15017
rect 52825 15008 52837 15011
rect 52604 14980 52837 15008
rect 52604 14968 52610 14980
rect 52825 14977 52837 14980
rect 52871 14977 52883 15011
rect 52825 14971 52883 14977
rect 53101 15011 53159 15017
rect 53101 14977 53113 15011
rect 53147 15008 53159 15011
rect 53374 15008 53380 15020
rect 53147 14980 53380 15008
rect 53147 14977 53159 14980
rect 53101 14971 53159 14977
rect 53374 14968 53380 14980
rect 53432 15008 53438 15020
rect 53929 15011 53987 15017
rect 53929 15008 53941 15011
rect 53432 14980 53941 15008
rect 53432 14968 53438 14980
rect 53929 14977 53941 14980
rect 53975 14977 53987 15011
rect 56778 15008 56784 15020
rect 56739 14980 56784 15008
rect 53929 14971 53987 14977
rect 56778 14968 56784 14980
rect 56836 14968 56842 15020
rect 56965 15011 57023 15017
rect 56965 14977 56977 15011
rect 57011 15008 57023 15011
rect 57054 15008 57060 15020
rect 57011 14980 57060 15008
rect 57011 14977 57023 14980
rect 56965 14971 57023 14977
rect 57054 14968 57060 14980
rect 57112 15008 57118 15020
rect 57882 15008 57888 15020
rect 57112 14980 57888 15008
rect 57112 14968 57118 14980
rect 57882 14968 57888 14980
rect 57940 14968 57946 15020
rect 52270 14900 52276 14952
rect 52328 14940 52334 14952
rect 53745 14943 53803 14949
rect 53745 14940 53757 14943
rect 52328 14912 53757 14940
rect 52328 14900 52334 14912
rect 53745 14909 53757 14912
rect 53791 14909 53803 14943
rect 53745 14903 53803 14909
rect 50062 14872 50068 14884
rect 48832 14844 50068 14872
rect 48832 14832 48838 14844
rect 50062 14832 50068 14844
rect 50120 14832 50126 14884
rect 52822 14832 52828 14884
rect 52880 14872 52886 14884
rect 52917 14875 52975 14881
rect 52917 14872 52929 14875
rect 52880 14844 52929 14872
rect 52880 14832 52886 14844
rect 52917 14841 52929 14844
rect 52963 14841 52975 14875
rect 52917 14835 52975 14841
rect 53006 14832 53012 14884
rect 53064 14872 53070 14884
rect 53064 14844 53109 14872
rect 53064 14832 53070 14844
rect 45888 14776 46520 14804
rect 46661 14807 46719 14813
rect 45888 14764 45894 14776
rect 46661 14773 46673 14807
rect 46707 14804 46719 14807
rect 46842 14804 46848 14816
rect 46707 14776 46848 14804
rect 46707 14773 46719 14776
rect 46661 14767 46719 14773
rect 46842 14764 46848 14776
rect 46900 14764 46906 14816
rect 48961 14807 49019 14813
rect 48961 14773 48973 14807
rect 49007 14804 49019 14807
rect 50154 14804 50160 14816
rect 49007 14776 50160 14804
rect 49007 14773 49019 14776
rect 48961 14767 49019 14773
rect 50154 14764 50160 14776
rect 50212 14804 50218 14816
rect 50525 14807 50583 14813
rect 50525 14804 50537 14807
rect 50212 14776 50537 14804
rect 50212 14764 50218 14776
rect 50525 14773 50537 14776
rect 50571 14773 50583 14807
rect 50525 14767 50583 14773
rect 53190 14764 53196 14816
rect 53248 14804 53254 14816
rect 53285 14807 53343 14813
rect 53285 14804 53297 14807
rect 53248 14776 53297 14804
rect 53248 14764 53254 14776
rect 53285 14773 53297 14776
rect 53331 14773 53343 14807
rect 53285 14767 53343 14773
rect 54205 14807 54263 14813
rect 54205 14773 54217 14807
rect 54251 14804 54263 14807
rect 54478 14804 54484 14816
rect 54251 14776 54484 14804
rect 54251 14773 54263 14776
rect 54205 14767 54263 14773
rect 54478 14764 54484 14776
rect 54536 14764 54542 14816
rect 1104 14714 58880 14736
rect 1104 14662 4214 14714
rect 4266 14662 4278 14714
rect 4330 14662 4342 14714
rect 4394 14662 4406 14714
rect 4458 14662 4470 14714
rect 4522 14662 34934 14714
rect 34986 14662 34998 14714
rect 35050 14662 35062 14714
rect 35114 14662 35126 14714
rect 35178 14662 35190 14714
rect 35242 14662 58880 14714
rect 1104 14640 58880 14662
rect 1486 14560 1492 14612
rect 1544 14600 1550 14612
rect 1581 14603 1639 14609
rect 1581 14600 1593 14603
rect 1544 14572 1593 14600
rect 1544 14560 1550 14572
rect 1581 14569 1593 14572
rect 1627 14569 1639 14603
rect 1581 14563 1639 14569
rect 3878 14560 3884 14612
rect 3936 14600 3942 14612
rect 4157 14603 4215 14609
rect 4157 14600 4169 14603
rect 3936 14572 4169 14600
rect 3936 14560 3942 14572
rect 4157 14569 4169 14572
rect 4203 14569 4215 14603
rect 6914 14600 6920 14612
rect 6875 14572 6920 14600
rect 4157 14563 4215 14569
rect 6914 14560 6920 14572
rect 6972 14560 6978 14612
rect 9769 14603 9827 14609
rect 9769 14569 9781 14603
rect 9815 14600 9827 14603
rect 10042 14600 10048 14612
rect 9815 14572 10048 14600
rect 9815 14569 9827 14572
rect 9769 14563 9827 14569
rect 10042 14560 10048 14572
rect 10100 14560 10106 14612
rect 10597 14603 10655 14609
rect 10597 14569 10609 14603
rect 10643 14600 10655 14603
rect 10778 14600 10784 14612
rect 10643 14572 10784 14600
rect 10643 14569 10655 14572
rect 10597 14563 10655 14569
rect 10778 14560 10784 14572
rect 10836 14560 10842 14612
rect 12253 14603 12311 14609
rect 12253 14569 12265 14603
rect 12299 14600 12311 14603
rect 12342 14600 12348 14612
rect 12299 14572 12348 14600
rect 12299 14569 12311 14572
rect 12253 14563 12311 14569
rect 12342 14560 12348 14572
rect 12400 14560 12406 14612
rect 13173 14603 13231 14609
rect 13173 14569 13185 14603
rect 13219 14600 13231 14603
rect 13446 14600 13452 14612
rect 13219 14572 13452 14600
rect 13219 14569 13231 14572
rect 13173 14563 13231 14569
rect 13446 14560 13452 14572
rect 13504 14560 13510 14612
rect 14550 14560 14556 14612
rect 14608 14600 14614 14612
rect 15838 14600 15844 14612
rect 14608 14572 15844 14600
rect 14608 14560 14614 14572
rect 15838 14560 15844 14572
rect 15896 14600 15902 14612
rect 16206 14600 16212 14612
rect 15896 14572 16212 14600
rect 15896 14560 15902 14572
rect 16206 14560 16212 14572
rect 16264 14560 16270 14612
rect 20070 14560 20076 14612
rect 20128 14600 20134 14612
rect 20441 14603 20499 14609
rect 20441 14600 20453 14603
rect 20128 14572 20453 14600
rect 20128 14560 20134 14572
rect 20441 14569 20453 14572
rect 20487 14569 20499 14603
rect 20441 14563 20499 14569
rect 20530 14560 20536 14612
rect 20588 14600 20594 14612
rect 22278 14600 22284 14612
rect 20588 14572 22284 14600
rect 20588 14560 20594 14572
rect 22278 14560 22284 14572
rect 22336 14560 22342 14612
rect 26878 14560 26884 14612
rect 26936 14600 26942 14612
rect 27249 14603 27307 14609
rect 27249 14600 27261 14603
rect 26936 14572 27261 14600
rect 26936 14560 26942 14572
rect 27249 14569 27261 14572
rect 27295 14569 27307 14603
rect 27249 14563 27307 14569
rect 28442 14560 28448 14612
rect 28500 14600 28506 14612
rect 30098 14600 30104 14612
rect 28500 14572 30104 14600
rect 28500 14560 28506 14572
rect 30098 14560 30104 14572
rect 30156 14560 30162 14612
rect 31018 14600 31024 14612
rect 30979 14572 31024 14600
rect 31018 14560 31024 14572
rect 31076 14560 31082 14612
rect 32214 14560 32220 14612
rect 32272 14600 32278 14612
rect 33229 14603 33287 14609
rect 33229 14600 33241 14603
rect 32272 14572 33241 14600
rect 32272 14560 32278 14572
rect 33229 14569 33241 14572
rect 33275 14569 33287 14603
rect 40034 14600 40040 14612
rect 39995 14572 40040 14600
rect 33229 14563 33287 14569
rect 40034 14560 40040 14572
rect 40092 14560 40098 14612
rect 43993 14603 44051 14609
rect 43993 14569 44005 14603
rect 44039 14569 44051 14603
rect 43993 14563 44051 14569
rect 50433 14603 50491 14609
rect 50433 14569 50445 14603
rect 50479 14600 50491 14603
rect 53006 14600 53012 14612
rect 50479 14572 53012 14600
rect 50479 14569 50491 14572
rect 50433 14563 50491 14569
rect 14366 14492 14372 14544
rect 14424 14532 14430 14544
rect 18414 14532 18420 14544
rect 14424 14504 18420 14532
rect 14424 14492 14430 14504
rect 18414 14492 18420 14504
rect 18472 14492 18478 14544
rect 21818 14532 21824 14544
rect 20088 14504 21824 14532
rect 7561 14467 7619 14473
rect 7561 14433 7573 14467
rect 7607 14464 7619 14467
rect 8938 14464 8944 14476
rect 7607 14436 8944 14464
rect 7607 14433 7619 14436
rect 7561 14427 7619 14433
rect 8938 14424 8944 14436
rect 8996 14464 9002 14476
rect 14090 14464 14096 14476
rect 8996 14436 14096 14464
rect 8996 14424 9002 14436
rect 14090 14424 14096 14436
rect 14148 14464 14154 14476
rect 14642 14464 14648 14476
rect 14148 14436 14648 14464
rect 14148 14424 14154 14436
rect 14642 14424 14648 14436
rect 14700 14424 14706 14476
rect 15764 14436 17816 14464
rect 1394 14396 1400 14408
rect 1355 14368 1400 14396
rect 1394 14356 1400 14368
rect 1452 14396 1458 14408
rect 2041 14399 2099 14405
rect 2041 14396 2053 14399
rect 1452 14368 2053 14396
rect 1452 14356 1458 14368
rect 2041 14365 2053 14368
rect 2087 14365 2099 14399
rect 2041 14359 2099 14365
rect 10318 14356 10324 14408
rect 10376 14396 10382 14408
rect 10413 14399 10471 14405
rect 10413 14396 10425 14399
rect 10376 14368 10425 14396
rect 10376 14356 10382 14368
rect 10413 14365 10425 14368
rect 10459 14365 10471 14399
rect 10413 14359 10471 14365
rect 15562 14356 15568 14408
rect 15620 14396 15626 14408
rect 15764 14405 15792 14436
rect 17788 14408 17816 14436
rect 15749 14399 15807 14405
rect 15749 14396 15761 14399
rect 15620 14368 15761 14396
rect 15620 14356 15626 14368
rect 15749 14365 15761 14368
rect 15795 14365 15807 14399
rect 15930 14396 15936 14408
rect 15891 14368 15936 14396
rect 15749 14359 15807 14365
rect 15930 14356 15936 14368
rect 15988 14356 15994 14408
rect 16117 14399 16175 14405
rect 16117 14365 16129 14399
rect 16163 14396 16175 14399
rect 16666 14396 16672 14408
rect 16163 14368 16672 14396
rect 16163 14365 16175 14368
rect 16117 14359 16175 14365
rect 16666 14356 16672 14368
rect 16724 14356 16730 14408
rect 16761 14399 16819 14405
rect 16761 14365 16773 14399
rect 16807 14365 16819 14399
rect 17218 14396 17224 14408
rect 17179 14368 17224 14396
rect 16761 14359 16819 14365
rect 3510 14288 3516 14340
rect 3568 14328 3574 14340
rect 3789 14331 3847 14337
rect 3789 14328 3801 14331
rect 3568 14300 3801 14328
rect 3568 14288 3574 14300
rect 3789 14297 3801 14300
rect 3835 14297 3847 14331
rect 3789 14291 3847 14297
rect 3973 14331 4031 14337
rect 3973 14297 3985 14331
rect 4019 14297 4031 14331
rect 3973 14291 4031 14297
rect 3988 14260 4016 14291
rect 6638 14288 6644 14340
rect 6696 14328 6702 14340
rect 6825 14331 6883 14337
rect 6825 14328 6837 14331
rect 6696 14300 6837 14328
rect 6696 14288 6702 14300
rect 6825 14297 6837 14300
rect 6871 14297 6883 14331
rect 16022 14328 16028 14340
rect 15983 14300 16028 14328
rect 6825 14291 6883 14297
rect 16022 14288 16028 14300
rect 16080 14288 16086 14340
rect 4154 14260 4160 14272
rect 3988 14232 4160 14260
rect 4154 14220 4160 14232
rect 4212 14260 4218 14272
rect 4706 14260 4712 14272
rect 4212 14232 4712 14260
rect 4212 14220 4218 14232
rect 4706 14220 4712 14232
rect 4764 14260 4770 14272
rect 5350 14260 5356 14272
rect 4764 14232 5356 14260
rect 4764 14220 4770 14232
rect 5350 14220 5356 14232
rect 5408 14220 5414 14272
rect 15010 14260 15016 14272
rect 14971 14232 15016 14260
rect 15010 14220 15016 14232
rect 15068 14220 15074 14272
rect 16301 14263 16359 14269
rect 16301 14229 16313 14263
rect 16347 14260 16359 14263
rect 16776 14260 16804 14359
rect 17218 14356 17224 14368
rect 17276 14356 17282 14408
rect 17770 14356 17776 14408
rect 17828 14396 17834 14408
rect 19889 14399 19947 14405
rect 19889 14396 19901 14399
rect 17828 14368 19901 14396
rect 17828 14356 17834 14368
rect 19889 14365 19901 14368
rect 19935 14396 19947 14399
rect 20088 14396 20116 14504
rect 21818 14492 21824 14504
rect 21876 14492 21882 14544
rect 31110 14532 31116 14544
rect 29932 14504 31116 14532
rect 20530 14464 20536 14476
rect 20180 14436 20536 14464
rect 20180 14405 20208 14436
rect 20530 14424 20536 14436
rect 20588 14424 20594 14476
rect 20806 14424 20812 14476
rect 20864 14464 20870 14476
rect 27982 14464 27988 14476
rect 20864 14436 21957 14464
rect 20864 14424 20870 14436
rect 19935 14368 20116 14396
rect 20165 14399 20223 14405
rect 19935 14365 19947 14368
rect 19889 14359 19947 14365
rect 20165 14365 20177 14399
rect 20211 14365 20223 14399
rect 20165 14359 20223 14365
rect 20254 14356 20260 14408
rect 20312 14396 20318 14408
rect 20990 14396 20996 14408
rect 20312 14368 20357 14396
rect 20951 14368 20996 14396
rect 20312 14356 20318 14368
rect 20990 14356 20996 14368
rect 21048 14356 21054 14408
rect 21174 14396 21180 14408
rect 21087 14368 21180 14396
rect 21174 14356 21180 14368
rect 21232 14396 21238 14408
rect 21634 14396 21640 14408
rect 21232 14368 21640 14396
rect 21232 14356 21238 14368
rect 21634 14356 21640 14368
rect 21692 14356 21698 14408
rect 17494 14328 17500 14340
rect 17455 14300 17500 14328
rect 17494 14288 17500 14300
rect 17552 14288 17558 14340
rect 19426 14288 19432 14340
rect 19484 14328 19490 14340
rect 20073 14331 20131 14337
rect 20073 14328 20085 14331
rect 19484 14300 20085 14328
rect 19484 14288 19490 14300
rect 20073 14297 20085 14300
rect 20119 14297 20131 14331
rect 21729 14331 21787 14337
rect 21729 14328 21741 14331
rect 20073 14291 20131 14297
rect 21100 14300 21741 14328
rect 16347 14232 16804 14260
rect 20088 14260 20116 14291
rect 21100 14260 21128 14300
rect 21729 14297 21741 14300
rect 21775 14297 21787 14331
rect 21929 14328 21957 14436
rect 22020 14436 27988 14464
rect 22020 14408 22048 14436
rect 27982 14424 27988 14436
rect 28040 14424 28046 14476
rect 28184 14436 28764 14464
rect 22002 14356 22008 14408
rect 22060 14356 22066 14408
rect 24946 14396 24952 14408
rect 24907 14368 24952 14396
rect 24946 14356 24952 14368
rect 25004 14356 25010 14408
rect 28074 14356 28080 14408
rect 28132 14396 28138 14408
rect 28184 14405 28212 14436
rect 28169 14399 28227 14405
rect 28169 14396 28181 14399
rect 28132 14368 28181 14396
rect 28132 14356 28138 14368
rect 28169 14365 28181 14368
rect 28215 14365 28227 14399
rect 28169 14359 28227 14365
rect 28534 14356 28540 14408
rect 28592 14396 28598 14408
rect 28592 14368 28637 14396
rect 28592 14356 28598 14368
rect 22370 14328 22376 14340
rect 21929 14300 22376 14328
rect 21729 14291 21787 14297
rect 22370 14288 22376 14300
rect 22428 14288 22434 14340
rect 24486 14288 24492 14340
rect 24544 14328 24550 14340
rect 24765 14331 24823 14337
rect 24765 14328 24777 14331
rect 24544 14300 24777 14328
rect 24544 14288 24550 14300
rect 24765 14297 24777 14300
rect 24811 14328 24823 14331
rect 26326 14328 26332 14340
rect 24811 14300 26332 14328
rect 24811 14297 24823 14300
rect 24765 14291 24823 14297
rect 26326 14288 26332 14300
rect 26384 14288 26390 14340
rect 28258 14328 28264 14340
rect 28219 14300 28264 14328
rect 28258 14288 28264 14300
rect 28316 14288 28322 14340
rect 28350 14288 28356 14340
rect 28408 14328 28414 14340
rect 28736 14328 28764 14436
rect 28810 14356 28816 14408
rect 28868 14396 28874 14408
rect 29932 14405 29960 14504
rect 31110 14492 31116 14504
rect 31168 14532 31174 14544
rect 33870 14532 33876 14544
rect 31168 14504 33876 14532
rect 31168 14492 31174 14504
rect 33870 14492 33876 14504
rect 33928 14532 33934 14544
rect 36541 14535 36599 14541
rect 33928 14504 35204 14532
rect 33928 14492 33934 14504
rect 33410 14464 33416 14476
rect 32405 14436 33416 14464
rect 29825 14399 29883 14405
rect 29825 14396 29837 14399
rect 28868 14368 29837 14396
rect 28868 14356 28874 14368
rect 29825 14365 29837 14368
rect 29871 14365 29883 14399
rect 29825 14359 29883 14365
rect 29917 14399 29975 14405
rect 29917 14365 29929 14399
rect 29963 14365 29975 14399
rect 29917 14359 29975 14365
rect 30193 14399 30251 14405
rect 30193 14365 30205 14399
rect 30239 14396 30251 14399
rect 30558 14396 30564 14408
rect 30239 14368 30564 14396
rect 30239 14365 30251 14368
rect 30193 14359 30251 14365
rect 30558 14356 30564 14368
rect 30616 14396 30622 14408
rect 31478 14396 31484 14408
rect 30616 14368 31484 14396
rect 30616 14356 30622 14368
rect 31478 14356 31484 14368
rect 31536 14356 31542 14408
rect 32030 14396 32036 14408
rect 31991 14368 32036 14396
rect 32030 14356 32036 14368
rect 32088 14356 32094 14408
rect 32122 14356 32128 14408
rect 32180 14396 32186 14408
rect 32180 14368 32225 14396
rect 32180 14356 32186 14368
rect 32306 14356 32312 14408
rect 32364 14396 32370 14408
rect 32405 14396 32433 14436
rect 33410 14424 33416 14436
rect 33468 14464 33474 14476
rect 34606 14464 34612 14476
rect 33468 14436 34612 14464
rect 33468 14424 33474 14436
rect 34606 14424 34612 14436
rect 34664 14424 34670 14476
rect 33505 14399 33563 14405
rect 32364 14368 32457 14396
rect 32364 14356 32370 14368
rect 33505 14365 33517 14399
rect 33551 14396 33563 14399
rect 34974 14396 34980 14408
rect 33551 14368 34980 14396
rect 33551 14365 33563 14368
rect 33505 14359 33563 14365
rect 34974 14356 34980 14368
rect 35032 14356 35038 14408
rect 35176 14405 35204 14504
rect 36541 14501 36553 14535
rect 36587 14532 36599 14535
rect 43898 14532 43904 14544
rect 36587 14504 43904 14532
rect 36587 14501 36599 14504
rect 36541 14495 36599 14501
rect 43898 14492 43904 14504
rect 43956 14532 43962 14544
rect 44008 14532 44036 14563
rect 53006 14560 53012 14572
rect 53064 14560 53070 14612
rect 53374 14600 53380 14612
rect 53335 14572 53380 14600
rect 53374 14560 53380 14572
rect 53432 14560 53438 14612
rect 43956 14504 44036 14532
rect 52917 14535 52975 14541
rect 43956 14492 43962 14504
rect 52917 14501 52929 14535
rect 52963 14532 52975 14535
rect 53558 14532 53564 14544
rect 52963 14504 53564 14532
rect 52963 14501 52975 14504
rect 52917 14495 52975 14501
rect 53558 14492 53564 14504
rect 53616 14492 53622 14544
rect 53745 14535 53803 14541
rect 53745 14501 53757 14535
rect 53791 14501 53803 14535
rect 53745 14495 53803 14501
rect 38289 14467 38347 14473
rect 38289 14433 38301 14467
rect 38335 14464 38347 14467
rect 38335 14436 39804 14464
rect 38335 14433 38347 14436
rect 38289 14427 38347 14433
rect 35161 14399 35219 14405
rect 35161 14365 35173 14399
rect 35207 14365 35219 14399
rect 35161 14359 35219 14365
rect 35621 14399 35679 14405
rect 35621 14365 35633 14399
rect 35667 14365 35679 14399
rect 35989 14399 36047 14405
rect 35989 14396 36001 14399
rect 35621 14359 35679 14365
rect 35728 14368 36001 14396
rect 30009 14331 30067 14337
rect 30009 14328 30021 14331
rect 28408 14300 28453 14328
rect 28736 14300 30021 14328
rect 28408 14288 28414 14300
rect 30009 14297 30021 14300
rect 30055 14328 30067 14331
rect 30926 14328 30932 14340
rect 30055 14300 30932 14328
rect 30055 14297 30067 14300
rect 30009 14291 30067 14297
rect 30926 14288 30932 14300
rect 30984 14288 30990 14340
rect 33045 14331 33103 14337
rect 33045 14328 33057 14331
rect 32405 14300 33057 14328
rect 21818 14260 21824 14272
rect 20088 14232 21128 14260
rect 21779 14232 21824 14260
rect 16347 14229 16359 14232
rect 16301 14223 16359 14229
rect 21818 14220 21824 14232
rect 21876 14220 21882 14272
rect 23658 14260 23664 14272
rect 23619 14232 23664 14260
rect 23658 14220 23664 14232
rect 23716 14220 23722 14272
rect 27982 14260 27988 14272
rect 27943 14232 27988 14260
rect 27982 14220 27988 14232
rect 28040 14220 28046 14272
rect 29638 14260 29644 14272
rect 29599 14232 29644 14260
rect 29638 14220 29644 14232
rect 29696 14220 29702 14272
rect 31386 14220 31392 14272
rect 31444 14260 31450 14272
rect 31481 14263 31539 14269
rect 31481 14260 31493 14263
rect 31444 14232 31493 14260
rect 31444 14220 31450 14232
rect 31481 14229 31493 14232
rect 31527 14260 31539 14263
rect 32405 14260 32433 14300
rect 33045 14297 33057 14300
rect 33091 14328 33103 14331
rect 33965 14331 34023 14337
rect 33965 14328 33977 14331
rect 33091 14300 33977 14328
rect 33091 14297 33103 14300
rect 33045 14291 33103 14297
rect 33965 14297 33977 14300
rect 34011 14297 34023 14331
rect 33965 14291 34023 14297
rect 34514 14288 34520 14340
rect 34572 14328 34578 14340
rect 35636 14328 35664 14359
rect 34572 14300 35664 14328
rect 34572 14288 34578 14300
rect 31527 14232 32433 14260
rect 32493 14263 32551 14269
rect 31527 14229 31539 14232
rect 31481 14223 31539 14229
rect 32493 14229 32505 14263
rect 32539 14260 32551 14263
rect 32950 14260 32956 14272
rect 32539 14232 32956 14260
rect 32539 14229 32551 14232
rect 32493 14223 32551 14229
rect 32950 14220 32956 14232
rect 33008 14220 33014 14272
rect 33229 14263 33287 14269
rect 33229 14229 33241 14263
rect 33275 14260 33287 14263
rect 33318 14260 33324 14272
rect 33275 14232 33324 14260
rect 33275 14229 33287 14232
rect 33229 14223 33287 14229
rect 33318 14220 33324 14232
rect 33376 14220 33382 14272
rect 33778 14220 33784 14272
rect 33836 14260 33842 14272
rect 35728 14260 35756 14368
rect 35989 14365 36001 14368
rect 36035 14365 36047 14399
rect 36354 14396 36360 14408
rect 36315 14368 36360 14396
rect 35989 14359 36047 14365
rect 36354 14356 36360 14368
rect 36412 14356 36418 14408
rect 37458 14356 37464 14408
rect 37516 14396 37522 14408
rect 37737 14399 37795 14405
rect 37737 14396 37749 14399
rect 37516 14368 37749 14396
rect 37516 14356 37522 14368
rect 37737 14365 37749 14368
rect 37783 14365 37795 14399
rect 38010 14396 38016 14408
rect 37971 14368 38016 14396
rect 37737 14359 37795 14365
rect 38010 14356 38016 14368
rect 38068 14356 38074 14408
rect 38381 14399 38439 14405
rect 38381 14365 38393 14399
rect 38427 14396 38439 14399
rect 38427 14368 38792 14396
rect 38427 14365 38439 14368
rect 38381 14359 38439 14365
rect 38764 14340 38792 14368
rect 38746 14288 38752 14340
rect 38804 14328 38810 14340
rect 38841 14331 38899 14337
rect 38841 14328 38853 14331
rect 38804 14300 38853 14328
rect 38804 14288 38810 14300
rect 38841 14297 38853 14300
rect 38887 14297 38899 14331
rect 38841 14291 38899 14297
rect 39025 14331 39083 14337
rect 39025 14297 39037 14331
rect 39071 14297 39083 14331
rect 39776 14328 39804 14436
rect 40034 14424 40040 14476
rect 40092 14464 40098 14476
rect 40681 14467 40739 14473
rect 40681 14464 40693 14467
rect 40092 14436 40693 14464
rect 40092 14424 40098 14436
rect 40681 14433 40693 14436
rect 40727 14433 40739 14467
rect 44082 14464 44088 14476
rect 44043 14436 44088 14464
rect 40681 14427 40739 14433
rect 44082 14424 44088 14436
rect 44140 14424 44146 14476
rect 44266 14424 44272 14476
rect 44324 14464 44330 14476
rect 45278 14464 45284 14476
rect 44324 14436 45284 14464
rect 44324 14424 44330 14436
rect 45278 14424 45284 14436
rect 45336 14464 45342 14476
rect 45336 14436 46152 14464
rect 45336 14424 45342 14436
rect 40770 14396 40776 14408
rect 40731 14368 40776 14396
rect 40770 14356 40776 14368
rect 40828 14356 40834 14408
rect 43990 14396 43996 14408
rect 43951 14368 43996 14396
rect 43990 14356 43996 14368
rect 44048 14356 44054 14408
rect 45830 14396 45836 14408
rect 45791 14368 45836 14396
rect 45830 14356 45836 14368
rect 45888 14356 45894 14408
rect 45922 14356 45928 14408
rect 45980 14396 45986 14408
rect 46124 14405 46152 14436
rect 52270 14424 52276 14476
rect 52328 14464 52334 14476
rect 53469 14467 53527 14473
rect 53469 14464 53481 14467
rect 52328 14436 53481 14464
rect 52328 14424 52334 14436
rect 53469 14433 53481 14436
rect 53515 14433 53527 14467
rect 53469 14427 53527 14433
rect 46109 14399 46167 14405
rect 45980 14368 46025 14396
rect 45980 14356 45986 14368
rect 46109 14365 46121 14399
rect 46155 14365 46167 14399
rect 50154 14396 50160 14408
rect 50115 14368 50160 14396
rect 46109 14359 46167 14365
rect 50154 14356 50160 14368
rect 50212 14356 50218 14408
rect 50246 14356 50252 14408
rect 50304 14396 50310 14408
rect 50304 14368 50349 14396
rect 50304 14356 50310 14368
rect 50430 14356 50436 14408
rect 50488 14396 50494 14408
rect 53377 14399 53435 14405
rect 50488 14368 50533 14396
rect 50488 14356 50494 14368
rect 53377 14365 53389 14399
rect 53423 14396 53435 14399
rect 53576 14396 53604 14492
rect 53760 14464 53788 14495
rect 53760 14436 54616 14464
rect 54478 14396 54484 14408
rect 53423 14368 53604 14396
rect 54439 14368 54484 14396
rect 53423 14365 53435 14368
rect 53377 14359 53435 14365
rect 54478 14356 54484 14368
rect 54536 14356 54542 14408
rect 54588 14405 54616 14436
rect 56318 14424 56324 14476
rect 56376 14464 56382 14476
rect 56689 14467 56747 14473
rect 56689 14464 56701 14467
rect 56376 14436 56701 14464
rect 56376 14424 56382 14436
rect 56689 14433 56701 14436
rect 56735 14433 56747 14467
rect 56689 14427 56747 14433
rect 54573 14399 54631 14405
rect 54573 14365 54585 14399
rect 54619 14365 54631 14399
rect 54573 14359 54631 14365
rect 54757 14399 54815 14405
rect 54757 14365 54769 14399
rect 54803 14396 54815 14399
rect 55490 14396 55496 14408
rect 54803 14368 55496 14396
rect 54803 14365 54815 14368
rect 54757 14359 54815 14365
rect 55490 14356 55496 14368
rect 55548 14396 55554 14408
rect 55769 14399 55827 14405
rect 55769 14396 55781 14399
rect 55548 14368 55781 14396
rect 55548 14356 55554 14368
rect 55769 14365 55781 14368
rect 55815 14365 55827 14399
rect 55769 14359 55827 14365
rect 55953 14399 56011 14405
rect 55953 14365 55965 14399
rect 55999 14365 56011 14399
rect 55953 14359 56011 14365
rect 48774 14328 48780 14340
rect 39776 14300 48780 14328
rect 39025 14291 39083 14297
rect 33836 14232 35756 14260
rect 33836 14220 33842 14232
rect 38378 14220 38384 14272
rect 38436 14260 38442 14272
rect 39040 14260 39068 14291
rect 48774 14288 48780 14300
rect 48832 14288 48838 14340
rect 55122 14288 55128 14340
rect 55180 14328 55186 14340
rect 55968 14328 55996 14359
rect 57330 14356 57336 14408
rect 57388 14396 57394 14408
rect 57885 14399 57943 14405
rect 57885 14396 57897 14399
rect 57388 14368 57897 14396
rect 57388 14356 57394 14368
rect 57885 14365 57897 14368
rect 57931 14365 57943 14399
rect 57885 14359 57943 14365
rect 55180 14300 55996 14328
rect 55180 14288 55186 14300
rect 38436 14232 39068 14260
rect 41141 14263 41199 14269
rect 38436 14220 38442 14232
rect 41141 14229 41153 14263
rect 41187 14260 41199 14263
rect 42334 14260 42340 14272
rect 41187 14232 42340 14260
rect 41187 14229 41199 14232
rect 41141 14223 41199 14229
rect 42334 14220 42340 14232
rect 42392 14220 42398 14272
rect 44361 14263 44419 14269
rect 44361 14229 44373 14263
rect 44407 14260 44419 14263
rect 45002 14260 45008 14272
rect 44407 14232 45008 14260
rect 44407 14229 44419 14232
rect 44361 14223 44419 14229
rect 45002 14220 45008 14232
rect 45060 14220 45066 14272
rect 46293 14263 46351 14269
rect 46293 14229 46305 14263
rect 46339 14260 46351 14263
rect 46934 14260 46940 14272
rect 46339 14232 46940 14260
rect 46339 14229 46351 14232
rect 46293 14223 46351 14229
rect 46934 14220 46940 14232
rect 46992 14220 46998 14272
rect 58066 14260 58072 14272
rect 58027 14232 58072 14260
rect 58066 14220 58072 14232
rect 58124 14220 58130 14272
rect 1104 14170 58880 14192
rect 1104 14118 19574 14170
rect 19626 14118 19638 14170
rect 19690 14118 19702 14170
rect 19754 14118 19766 14170
rect 19818 14118 19830 14170
rect 19882 14118 50294 14170
rect 50346 14118 50358 14170
rect 50410 14118 50422 14170
rect 50474 14118 50486 14170
rect 50538 14118 50550 14170
rect 50602 14118 58880 14170
rect 1104 14096 58880 14118
rect 13725 14059 13783 14065
rect 13725 14025 13737 14059
rect 13771 14056 13783 14059
rect 16482 14056 16488 14068
rect 13771 14028 16488 14056
rect 13771 14025 13783 14028
rect 13725 14019 13783 14025
rect 16482 14016 16488 14028
rect 16540 14016 16546 14068
rect 22094 14056 22100 14068
rect 21560 14028 22100 14056
rect 4154 13988 4160 14000
rect 3436 13960 4160 13988
rect 3436 13929 3464 13960
rect 4154 13948 4160 13960
rect 4212 13948 4218 14000
rect 12526 13988 12532 14000
rect 9600 13960 11008 13988
rect 12487 13960 12532 13988
rect 3421 13923 3479 13929
rect 3421 13889 3433 13923
rect 3467 13889 3479 13923
rect 3421 13883 3479 13889
rect 3510 13880 3516 13932
rect 3568 13920 3574 13932
rect 9600 13929 9628 13960
rect 3973 13923 4031 13929
rect 3973 13920 3985 13923
rect 3568 13892 3985 13920
rect 3568 13880 3574 13892
rect 3973 13889 3985 13892
rect 4019 13889 4031 13923
rect 3973 13883 4031 13889
rect 9585 13923 9643 13929
rect 9585 13889 9597 13923
rect 9631 13889 9643 13923
rect 9585 13883 9643 13889
rect 9674 13880 9680 13932
rect 9732 13920 9738 13932
rect 10229 13923 10287 13929
rect 10229 13920 10241 13923
rect 9732 13892 10241 13920
rect 9732 13880 9738 13892
rect 10229 13889 10241 13892
rect 10275 13889 10287 13923
rect 10229 13883 10287 13889
rect 10980 13864 11008 13960
rect 12526 13948 12532 13960
rect 12584 13988 12590 14000
rect 14366 13988 14372 14000
rect 12584 13960 13400 13988
rect 12584 13948 12590 13960
rect 13372 13929 13400 13960
rect 13556 13960 14372 13988
rect 13556 13929 13584 13960
rect 14366 13948 14372 13960
rect 14424 13948 14430 14000
rect 15746 13988 15752 14000
rect 15707 13960 15752 13988
rect 15746 13948 15752 13960
rect 15804 13948 15810 14000
rect 16206 13988 16212 14000
rect 16040 13960 16212 13988
rect 16040 13954 16068 13960
rect 12713 13923 12771 13929
rect 12713 13889 12725 13923
rect 12759 13920 12771 13923
rect 13357 13923 13415 13929
rect 12759 13892 12848 13920
rect 12759 13889 12771 13892
rect 12713 13883 12771 13889
rect 5350 13852 5356 13864
rect 5311 13824 5356 13852
rect 5350 13812 5356 13824
rect 5408 13812 5414 13864
rect 7374 13812 7380 13864
rect 7432 13852 7438 13864
rect 8021 13855 8079 13861
rect 8021 13852 8033 13855
rect 7432 13824 8033 13852
rect 7432 13812 7438 13824
rect 8021 13821 8033 13824
rect 8067 13821 8079 13855
rect 8021 13815 8079 13821
rect 10962 13812 10968 13864
rect 11020 13852 11026 13864
rect 11517 13855 11575 13861
rect 11517 13852 11529 13855
rect 11020 13824 11529 13852
rect 11020 13812 11026 13824
rect 11517 13821 11529 13824
rect 11563 13821 11575 13855
rect 11517 13815 11575 13821
rect 4614 13784 4620 13796
rect 4575 13756 4620 13784
rect 4614 13744 4620 13756
rect 4672 13744 4678 13796
rect 8757 13787 8815 13793
rect 8757 13753 8769 13787
rect 8803 13784 8815 13787
rect 8846 13784 8852 13796
rect 8803 13756 8852 13784
rect 8803 13753 8815 13756
rect 8757 13747 8815 13753
rect 8846 13744 8852 13756
rect 8904 13744 8910 13796
rect 12820 13716 12848 13892
rect 13357 13889 13369 13923
rect 13403 13889 13415 13923
rect 13357 13883 13415 13889
rect 13541 13923 13599 13929
rect 13541 13889 13553 13923
rect 13587 13889 13599 13923
rect 13541 13883 13599 13889
rect 14274 13880 14280 13932
rect 14332 13920 14338 13932
rect 15013 13923 15071 13929
rect 15013 13920 15025 13923
rect 14332 13892 15025 13920
rect 14332 13880 14338 13892
rect 15013 13889 15025 13892
rect 15059 13889 15071 13923
rect 15562 13920 15568 13932
rect 15523 13892 15568 13920
rect 15013 13883 15071 13889
rect 15562 13880 15568 13892
rect 15620 13880 15626 13932
rect 15838 13920 15844 13932
rect 15799 13892 15844 13920
rect 15838 13880 15844 13892
rect 15896 13880 15902 13932
rect 15948 13926 16068 13954
rect 16206 13948 16212 13960
rect 16264 13948 16270 14000
rect 16298 13948 16304 14000
rect 16356 13988 16362 14000
rect 20806 13988 20812 14000
rect 16356 13960 20812 13988
rect 16356 13948 16362 13960
rect 20806 13948 20812 13960
rect 20864 13948 20870 14000
rect 21560 13988 21588 14028
rect 22094 14016 22100 14028
rect 22152 14016 22158 14068
rect 22370 14016 22376 14068
rect 22428 14016 22434 14068
rect 23382 14016 23388 14068
rect 23440 14056 23446 14068
rect 25777 14059 25835 14065
rect 25777 14056 25789 14059
rect 23440 14028 25789 14056
rect 23440 14016 23446 14028
rect 25777 14025 25789 14028
rect 25823 14056 25835 14059
rect 26234 14056 26240 14068
rect 25823 14028 26240 14056
rect 25823 14025 25835 14028
rect 25777 14019 25835 14025
rect 26234 14016 26240 14028
rect 26292 14016 26298 14068
rect 26326 14016 26332 14068
rect 26384 14056 26390 14068
rect 28626 14056 28632 14068
rect 26384 14028 28632 14056
rect 26384 14016 26390 14028
rect 28626 14016 28632 14028
rect 28684 14056 28690 14068
rect 29914 14056 29920 14068
rect 28684 14028 29920 14056
rect 28684 14016 28690 14028
rect 29914 14016 29920 14028
rect 29972 14016 29978 14068
rect 31021 14059 31079 14065
rect 31021 14025 31033 14059
rect 31067 14056 31079 14059
rect 32306 14056 32312 14068
rect 31067 14028 32312 14056
rect 31067 14025 31079 14028
rect 31021 14019 31079 14025
rect 32306 14016 32312 14028
rect 32364 14016 32370 14068
rect 32861 14059 32919 14065
rect 32861 14025 32873 14059
rect 32907 14056 32919 14059
rect 38010 14056 38016 14068
rect 32907 14028 38016 14056
rect 32907 14025 32919 14028
rect 32861 14019 32919 14025
rect 38010 14016 38016 14028
rect 38068 14016 38074 14068
rect 49786 14016 49792 14068
rect 49844 14056 49850 14068
rect 50433 14059 50491 14065
rect 50433 14056 50445 14059
rect 49844 14028 50445 14056
rect 49844 14016 49850 14028
rect 50433 14025 50445 14028
rect 50479 14056 50491 14059
rect 50706 14056 50712 14068
rect 50479 14028 50712 14056
rect 50479 14025 50491 14028
rect 50433 14019 50491 14025
rect 50706 14016 50712 14028
rect 50764 14016 50770 14068
rect 57882 14056 57888 14068
rect 57843 14028 57888 14056
rect 57882 14016 57888 14028
rect 57940 14016 57946 14068
rect 21008 13960 21588 13988
rect 15948 13923 16015 13926
rect 15948 13892 15969 13923
rect 15957 13889 15969 13892
rect 16003 13889 16015 13923
rect 16666 13920 16672 13932
rect 16627 13892 16672 13920
rect 15957 13883 16015 13889
rect 16666 13880 16672 13892
rect 16724 13880 16730 13932
rect 20162 13920 20168 13932
rect 20123 13892 20168 13920
rect 20162 13880 20168 13892
rect 20220 13880 20226 13932
rect 20346 13880 20352 13932
rect 20404 13920 20410 13932
rect 20717 13923 20775 13929
rect 20717 13920 20729 13923
rect 20404 13892 20729 13920
rect 20404 13880 20410 13892
rect 20717 13889 20729 13892
rect 20763 13889 20775 13923
rect 20898 13920 20904 13932
rect 20859 13892 20904 13920
rect 20717 13883 20775 13889
rect 20898 13880 20904 13892
rect 20956 13880 20962 13932
rect 21008 13929 21036 13960
rect 21634 13948 21640 14000
rect 21692 13988 21698 14000
rect 22189 13991 22247 13997
rect 21692 13960 22140 13988
rect 21692 13948 21698 13960
rect 20993 13923 21051 13929
rect 20993 13889 21005 13923
rect 21039 13889 21051 13923
rect 20993 13883 21051 13889
rect 21085 13923 21143 13929
rect 21085 13889 21097 13923
rect 21131 13918 21143 13923
rect 21821 13923 21879 13929
rect 21821 13920 21833 13923
rect 21131 13890 21220 13918
rect 21131 13889 21143 13890
rect 21085 13883 21143 13889
rect 12897 13855 12955 13861
rect 12897 13821 12909 13855
rect 12943 13852 12955 13855
rect 16942 13852 16948 13864
rect 12943 13824 15700 13852
rect 16855 13824 16948 13852
rect 12943 13821 12955 13824
rect 12897 13815 12955 13821
rect 13354 13716 13360 13728
rect 12820 13688 13360 13716
rect 13354 13676 13360 13688
rect 13412 13676 13418 13728
rect 15672 13716 15700 13824
rect 16942 13812 16948 13824
rect 17000 13852 17006 13864
rect 17862 13852 17868 13864
rect 17000 13824 17868 13852
rect 17000 13812 17006 13824
rect 17862 13812 17868 13824
rect 17920 13812 17926 13864
rect 20254 13812 20260 13864
rect 20312 13852 20318 13864
rect 21192 13852 21220 13890
rect 20312 13824 21220 13852
rect 21284 13892 21833 13920
rect 20312 13812 20318 13824
rect 21008 13796 21036 13824
rect 19981 13787 20039 13793
rect 15948 13756 17448 13784
rect 15948 13716 15976 13756
rect 16114 13716 16120 13728
rect 15672 13688 15976 13716
rect 16075 13688 16120 13716
rect 16114 13676 16120 13688
rect 16172 13676 16178 13728
rect 17420 13716 17448 13756
rect 19981 13753 19993 13787
rect 20027 13784 20039 13787
rect 20162 13784 20168 13796
rect 20027 13756 20168 13784
rect 20027 13753 20039 13756
rect 19981 13747 20039 13753
rect 20162 13744 20168 13756
rect 20220 13744 20226 13796
rect 20990 13744 20996 13796
rect 21048 13744 21054 13796
rect 21284 13793 21312 13892
rect 21821 13889 21833 13892
rect 21867 13889 21879 13923
rect 21821 13883 21879 13889
rect 21910 13880 21916 13932
rect 21968 13920 21974 13932
rect 22112 13929 22140 13960
rect 22189 13957 22201 13991
rect 22235 13988 22247 13991
rect 22388 13988 22416 14016
rect 23658 13988 23664 14000
rect 22235 13960 22416 13988
rect 23492 13960 23664 13988
rect 22235 13957 22247 13960
rect 22189 13951 22247 13957
rect 22097 13923 22155 13929
rect 21968 13892 22013 13920
rect 21968 13880 21974 13892
rect 22097 13889 22109 13923
rect 22143 13889 22155 13923
rect 22097 13883 22155 13889
rect 22327 13923 22385 13929
rect 22327 13889 22339 13923
rect 22373 13920 22385 13923
rect 22830 13920 22836 13932
rect 22373 13892 22836 13920
rect 22373 13889 22385 13892
rect 22327 13883 22385 13889
rect 22830 13880 22836 13892
rect 22888 13880 22894 13932
rect 22922 13880 22928 13932
rect 22980 13920 22986 13932
rect 23492 13929 23520 13960
rect 23658 13948 23664 13960
rect 23716 13988 23722 14000
rect 27338 13988 27344 14000
rect 23716 13960 27344 13988
rect 23716 13948 23722 13960
rect 27338 13948 27344 13960
rect 27396 13948 27402 14000
rect 28169 13991 28227 13997
rect 28169 13957 28181 13991
rect 28215 13988 28227 13991
rect 28994 13988 29000 14000
rect 28215 13960 29000 13988
rect 28215 13957 28227 13960
rect 28169 13951 28227 13957
rect 28994 13948 29000 13960
rect 29052 13948 29058 14000
rect 29730 13948 29736 14000
rect 29788 13988 29794 14000
rect 31110 13988 31116 14000
rect 29788 13960 31116 13988
rect 29788 13948 29794 13960
rect 31110 13948 31116 13960
rect 31168 13988 31174 14000
rect 31481 13991 31539 13997
rect 31481 13988 31493 13991
rect 31168 13960 31493 13988
rect 31168 13948 31174 13960
rect 31481 13957 31493 13960
rect 31527 13988 31539 13991
rect 31527 13960 32628 13988
rect 31527 13957 31539 13960
rect 31481 13951 31539 13957
rect 32600 13932 32628 13960
rect 33226 13948 33232 14000
rect 33284 13988 33290 14000
rect 33321 13991 33379 13997
rect 33321 13988 33333 13991
rect 33284 13960 33333 13988
rect 33284 13948 33290 13960
rect 33321 13957 33333 13960
rect 33367 13957 33379 13991
rect 37277 13991 37335 13997
rect 37277 13988 37289 13991
rect 33321 13951 33379 13957
rect 33704 13960 37289 13988
rect 23293 13923 23351 13929
rect 23293 13920 23305 13923
rect 22980 13892 23305 13920
rect 22980 13880 22986 13892
rect 23293 13889 23305 13892
rect 23339 13889 23351 13923
rect 23293 13883 23351 13889
rect 23477 13923 23535 13929
rect 23477 13889 23489 13923
rect 23523 13889 23535 13923
rect 23477 13883 23535 13889
rect 21269 13787 21327 13793
rect 21269 13753 21281 13787
rect 21315 13753 21327 13787
rect 21269 13747 21327 13753
rect 21358 13744 21364 13796
rect 21416 13784 21422 13796
rect 23492 13784 23520 13883
rect 24394 13880 24400 13932
rect 24452 13920 24458 13932
rect 24489 13923 24547 13929
rect 24489 13920 24501 13923
rect 24452 13892 24501 13920
rect 24452 13880 24458 13892
rect 24489 13889 24501 13892
rect 24535 13889 24547 13923
rect 24489 13883 24547 13889
rect 24762 13880 24768 13932
rect 24820 13920 24826 13932
rect 27985 13923 28043 13929
rect 27985 13920 27997 13923
rect 24820 13892 27997 13920
rect 24820 13880 24826 13892
rect 27985 13889 27997 13892
rect 28031 13920 28043 13923
rect 30098 13920 30104 13932
rect 28031 13892 30104 13920
rect 28031 13889 28043 13892
rect 27985 13883 28043 13889
rect 30098 13880 30104 13892
rect 30156 13880 30162 13932
rect 32490 13920 32496 13932
rect 32451 13892 32496 13920
rect 32490 13880 32496 13892
rect 32548 13880 32554 13932
rect 32582 13880 32588 13932
rect 32640 13920 32646 13932
rect 32640 13892 32733 13920
rect 32640 13880 32646 13892
rect 24673 13855 24731 13861
rect 24673 13821 24685 13855
rect 24719 13852 24731 13855
rect 24946 13852 24952 13864
rect 24719 13824 24952 13852
rect 24719 13821 24731 13824
rect 24673 13815 24731 13821
rect 24946 13812 24952 13824
rect 25004 13812 25010 13864
rect 28258 13812 28264 13864
rect 28316 13852 28322 13864
rect 33704 13852 33732 13960
rect 37277 13957 37289 13960
rect 37323 13988 37335 13991
rect 39114 13988 39120 14000
rect 37323 13960 39120 13988
rect 37323 13957 37335 13960
rect 37277 13951 37335 13957
rect 39114 13948 39120 13960
rect 39172 13948 39178 14000
rect 44177 13991 44235 13997
rect 44177 13957 44189 13991
rect 44223 13988 44235 13991
rect 45094 13988 45100 14000
rect 44223 13960 45100 13988
rect 44223 13957 44235 13960
rect 44177 13951 44235 13957
rect 45094 13948 45100 13960
rect 45152 13948 45158 14000
rect 56873 13991 56931 13997
rect 56873 13957 56885 13991
rect 56919 13988 56931 13991
rect 56919 13960 58112 13988
rect 56919 13957 56931 13960
rect 56873 13951 56931 13957
rect 33778 13880 33784 13932
rect 33836 13920 33842 13932
rect 34425 13923 34483 13929
rect 34425 13920 34437 13923
rect 33836 13892 34437 13920
rect 33836 13880 33842 13892
rect 34425 13889 34437 13892
rect 34471 13889 34483 13923
rect 34974 13920 34980 13932
rect 34935 13892 34980 13920
rect 34425 13883 34483 13889
rect 34974 13880 34980 13892
rect 35032 13880 35038 13932
rect 35253 13923 35311 13929
rect 35253 13889 35265 13923
rect 35299 13920 35311 13923
rect 35802 13920 35808 13932
rect 35299 13892 35808 13920
rect 35299 13889 35311 13892
rect 35253 13883 35311 13889
rect 35802 13880 35808 13892
rect 35860 13880 35866 13932
rect 36449 13923 36507 13929
rect 36449 13889 36461 13923
rect 36495 13920 36507 13923
rect 37182 13920 37188 13932
rect 36495 13892 37188 13920
rect 36495 13889 36507 13892
rect 36449 13883 36507 13889
rect 37182 13880 37188 13892
rect 37240 13880 37246 13932
rect 37366 13880 37372 13932
rect 37424 13920 37430 13932
rect 37461 13923 37519 13929
rect 37461 13920 37473 13923
rect 37424 13892 37473 13920
rect 37424 13880 37430 13892
rect 37461 13889 37473 13892
rect 37507 13889 37519 13923
rect 37461 13883 37519 13889
rect 38197 13923 38255 13929
rect 38197 13889 38209 13923
rect 38243 13920 38255 13923
rect 38746 13920 38752 13932
rect 38243 13892 38752 13920
rect 38243 13889 38255 13892
rect 38197 13883 38255 13889
rect 38746 13880 38752 13892
rect 38804 13880 38810 13932
rect 43898 13920 43904 13932
rect 43859 13892 43904 13920
rect 43898 13880 43904 13892
rect 43956 13880 43962 13932
rect 43990 13880 43996 13932
rect 44048 13920 44054 13932
rect 53190 13920 53196 13932
rect 44048 13892 44093 13920
rect 53151 13892 53196 13920
rect 44048 13880 44054 13892
rect 53190 13880 53196 13892
rect 53248 13880 53254 13932
rect 53837 13923 53895 13929
rect 53837 13889 53849 13923
rect 53883 13920 53895 13923
rect 55122 13920 55128 13932
rect 53883 13892 55128 13920
rect 53883 13889 53895 13892
rect 53837 13883 53895 13889
rect 55122 13880 55128 13892
rect 55180 13920 55186 13932
rect 55309 13923 55367 13929
rect 55309 13920 55321 13923
rect 55180 13892 55321 13920
rect 55180 13880 55186 13892
rect 55309 13889 55321 13892
rect 55355 13889 55367 13923
rect 55490 13920 55496 13932
rect 55451 13892 55496 13920
rect 55309 13883 55367 13889
rect 55490 13880 55496 13892
rect 55548 13880 55554 13932
rect 56594 13920 56600 13932
rect 56555 13892 56600 13920
rect 56594 13880 56600 13892
rect 56652 13880 56658 13932
rect 57882 13920 57888 13932
rect 57843 13892 57888 13920
rect 57882 13880 57888 13892
rect 57940 13880 57946 13932
rect 58084 13929 58112 13960
rect 58069 13923 58127 13929
rect 58069 13889 58081 13923
rect 58115 13889 58127 13923
rect 58069 13883 58127 13889
rect 28316 13824 33732 13852
rect 28316 13812 28322 13824
rect 34514 13812 34520 13864
rect 34572 13812 34578 13864
rect 38105 13855 38163 13861
rect 38105 13852 38117 13855
rect 34992 13824 38117 13852
rect 21416 13756 23520 13784
rect 21416 13744 21422 13756
rect 27798 13744 27804 13796
rect 27856 13784 27862 13796
rect 34241 13787 34299 13793
rect 34241 13784 34253 13787
rect 27856 13756 34253 13784
rect 27856 13744 27862 13756
rect 34241 13753 34253 13756
rect 34287 13753 34299 13787
rect 34241 13747 34299 13753
rect 22278 13716 22284 13728
rect 17420 13688 22284 13716
rect 22278 13676 22284 13688
rect 22336 13676 22342 13728
rect 22462 13716 22468 13728
rect 22423 13688 22468 13716
rect 22462 13676 22468 13688
rect 22520 13676 22526 13728
rect 23106 13716 23112 13728
rect 23067 13688 23112 13716
rect 23106 13676 23112 13688
rect 23164 13676 23170 13728
rect 25130 13716 25136 13728
rect 25091 13688 25136 13716
rect 25130 13676 25136 13688
rect 25188 13676 25194 13728
rect 32674 13716 32680 13728
rect 32587 13688 32680 13716
rect 32674 13676 32680 13688
rect 32732 13716 32738 13728
rect 33226 13716 33232 13728
rect 32732 13688 33232 13716
rect 32732 13676 32738 13688
rect 33226 13676 33232 13688
rect 33284 13676 33290 13728
rect 34054 13676 34060 13728
rect 34112 13716 34118 13728
rect 34992 13716 35020 13824
rect 38105 13821 38117 13824
rect 38151 13821 38163 13855
rect 38105 13815 38163 13821
rect 44082 13812 44088 13864
rect 44140 13852 44146 13864
rect 44177 13855 44235 13861
rect 44177 13852 44189 13855
rect 44140 13824 44189 13852
rect 44140 13812 44146 13824
rect 44177 13821 44189 13824
rect 44223 13821 44235 13855
rect 53006 13852 53012 13864
rect 52967 13824 53012 13852
rect 44177 13815 44235 13821
rect 53006 13812 53012 13824
rect 53064 13812 53070 13864
rect 54478 13812 54484 13864
rect 54536 13852 54542 13864
rect 56870 13852 56876 13864
rect 54536 13824 56876 13852
rect 54536 13812 54542 13824
rect 56870 13812 56876 13824
rect 56928 13812 56934 13864
rect 36170 13716 36176 13728
rect 34112 13688 35020 13716
rect 36131 13688 36176 13716
rect 34112 13676 34118 13688
rect 36170 13676 36176 13688
rect 36228 13676 36234 13728
rect 38473 13719 38531 13725
rect 38473 13685 38485 13719
rect 38519 13716 38531 13719
rect 40770 13716 40776 13728
rect 38519 13688 40776 13716
rect 38519 13685 38531 13688
rect 38473 13679 38531 13685
rect 40770 13676 40776 13688
rect 40828 13676 40834 13728
rect 55398 13716 55404 13728
rect 55359 13688 55404 13716
rect 55398 13676 55404 13688
rect 55456 13676 55462 13728
rect 56689 13719 56747 13725
rect 56689 13685 56701 13719
rect 56735 13716 56747 13719
rect 56778 13716 56784 13728
rect 56735 13688 56784 13716
rect 56735 13685 56747 13688
rect 56689 13679 56747 13685
rect 56778 13676 56784 13688
rect 56836 13676 56842 13728
rect 1104 13626 58880 13648
rect 1104 13574 4214 13626
rect 4266 13574 4278 13626
rect 4330 13574 4342 13626
rect 4394 13574 4406 13626
rect 4458 13574 4470 13626
rect 4522 13574 34934 13626
rect 34986 13574 34998 13626
rect 35050 13574 35062 13626
rect 35114 13574 35126 13626
rect 35178 13574 35190 13626
rect 35242 13574 58880 13626
rect 1104 13552 58880 13574
rect 7926 13512 7932 13524
rect 7887 13484 7932 13512
rect 7926 13472 7932 13484
rect 7984 13472 7990 13524
rect 9674 13512 9680 13524
rect 9635 13484 9680 13512
rect 9674 13472 9680 13484
rect 9732 13472 9738 13524
rect 15654 13512 15660 13524
rect 12820 13484 15660 13512
rect 3234 13444 3240 13456
rect 2240 13416 3240 13444
rect 2240 13385 2268 13416
rect 3234 13404 3240 13416
rect 3292 13404 3298 13456
rect 9585 13447 9643 13453
rect 9585 13413 9597 13447
rect 9631 13444 9643 13447
rect 9858 13444 9864 13456
rect 9631 13416 9864 13444
rect 9631 13413 9643 13416
rect 9585 13407 9643 13413
rect 9858 13404 9864 13416
rect 9916 13444 9922 13456
rect 10689 13447 10747 13453
rect 10689 13444 10701 13447
rect 9916 13416 10701 13444
rect 9916 13404 9922 13416
rect 10689 13413 10701 13416
rect 10735 13413 10747 13447
rect 12342 13444 12348 13456
rect 12303 13416 12348 13444
rect 10689 13407 10747 13413
rect 12342 13404 12348 13416
rect 12400 13404 12406 13456
rect 12820 13385 12848 13484
rect 15654 13472 15660 13484
rect 15712 13472 15718 13524
rect 17494 13472 17500 13524
rect 17552 13512 17558 13524
rect 17552 13484 24072 13512
rect 17552 13472 17558 13484
rect 18230 13444 18236 13456
rect 12912 13416 18236 13444
rect 2225 13379 2283 13385
rect 2225 13345 2237 13379
rect 2271 13345 2283 13379
rect 2225 13339 2283 13345
rect 12805 13379 12863 13385
rect 12805 13345 12817 13379
rect 12851 13345 12863 13379
rect 12805 13339 12863 13345
rect 2961 13311 3019 13317
rect 2961 13277 2973 13311
rect 3007 13277 3019 13311
rect 3142 13308 3148 13320
rect 3103 13280 3148 13308
rect 2961 13271 3019 13277
rect 2976 13240 3004 13271
rect 3142 13268 3148 13280
rect 3200 13268 3206 13320
rect 6362 13268 6368 13320
rect 6420 13308 6426 13320
rect 6457 13311 6515 13317
rect 6457 13308 6469 13311
rect 6420 13280 6469 13308
rect 6420 13268 6426 13280
rect 6457 13277 6469 13280
rect 6503 13277 6515 13311
rect 7374 13308 7380 13320
rect 6457 13271 6515 13277
rect 6564 13280 7380 13308
rect 3050 13240 3056 13252
rect 2976 13212 3056 13240
rect 3050 13200 3056 13212
rect 3108 13200 3114 13252
rect 6270 13200 6276 13252
rect 6328 13240 6334 13252
rect 6564 13240 6592 13280
rect 7374 13268 7380 13280
rect 7432 13268 7438 13320
rect 12912 13308 12940 13416
rect 18230 13404 18236 13416
rect 18288 13404 18294 13456
rect 20162 13404 20168 13456
rect 20220 13444 20226 13456
rect 22830 13444 22836 13456
rect 20220 13416 22836 13444
rect 20220 13404 20226 13416
rect 22830 13404 22836 13416
rect 22888 13404 22894 13456
rect 23750 13444 23756 13456
rect 23711 13416 23756 13444
rect 23750 13404 23756 13416
rect 23808 13404 23814 13456
rect 15378 13336 15384 13388
rect 15436 13376 15442 13388
rect 15565 13379 15623 13385
rect 15565 13376 15577 13379
rect 15436 13348 15577 13376
rect 15436 13336 15442 13348
rect 15565 13345 15577 13348
rect 15611 13376 15623 13379
rect 21358 13376 21364 13388
rect 15611 13348 17724 13376
rect 15611 13345 15623 13348
rect 15565 13339 15623 13345
rect 14550 13308 14556 13320
rect 12820 13280 12940 13308
rect 14511 13280 14556 13308
rect 12820 13249 12848 13280
rect 14550 13268 14556 13280
rect 14608 13268 14614 13320
rect 16022 13308 16028 13320
rect 15983 13280 16028 13308
rect 16022 13268 16028 13280
rect 16080 13268 16086 13320
rect 16393 13311 16451 13317
rect 16393 13277 16405 13311
rect 16439 13308 16451 13311
rect 16942 13308 16948 13320
rect 16439 13280 16948 13308
rect 16439 13277 16451 13280
rect 16393 13271 16451 13277
rect 16942 13268 16948 13280
rect 17000 13268 17006 13320
rect 17402 13268 17408 13320
rect 17460 13308 17466 13320
rect 17696 13317 17724 13348
rect 17972 13348 21364 13376
rect 17497 13311 17555 13317
rect 17497 13308 17509 13311
rect 17460 13280 17509 13308
rect 17460 13268 17466 13280
rect 17497 13277 17509 13280
rect 17543 13277 17555 13311
rect 17497 13271 17555 13277
rect 17681 13311 17739 13317
rect 17681 13277 17693 13311
rect 17727 13277 17739 13311
rect 17862 13308 17868 13320
rect 17823 13280 17868 13308
rect 17681 13271 17739 13277
rect 17862 13268 17868 13280
rect 17920 13268 17926 13320
rect 6328 13212 6592 13240
rect 9217 13243 9275 13249
rect 6328 13200 6334 13212
rect 9217 13209 9229 13243
rect 9263 13209 9275 13243
rect 9217 13203 9275 13209
rect 12805 13243 12863 13249
rect 12805 13209 12817 13243
rect 12851 13209 12863 13243
rect 12805 13203 12863 13209
rect 12897 13243 12955 13249
rect 12897 13209 12909 13243
rect 12943 13240 12955 13243
rect 13078 13240 13084 13252
rect 12943 13212 13084 13240
rect 12943 13209 12955 13212
rect 12897 13203 12955 13209
rect 9232 13172 9260 13203
rect 9674 13172 9680 13184
rect 9232 13144 9680 13172
rect 9674 13132 9680 13144
rect 9732 13172 9738 13184
rect 10229 13175 10287 13181
rect 10229 13172 10241 13175
rect 9732 13144 10241 13172
rect 9732 13132 9738 13144
rect 10229 13141 10241 13144
rect 10275 13172 10287 13175
rect 10870 13172 10876 13184
rect 10275 13144 10876 13172
rect 10275 13141 10287 13144
rect 10229 13135 10287 13141
rect 10870 13132 10876 13144
rect 10928 13132 10934 13184
rect 11793 13175 11851 13181
rect 11793 13141 11805 13175
rect 11839 13172 11851 13175
rect 12820 13172 12848 13203
rect 13078 13200 13084 13212
rect 13136 13200 13142 13252
rect 13170 13200 13176 13252
rect 13228 13240 13234 13252
rect 13541 13243 13599 13249
rect 13541 13240 13553 13243
rect 13228 13212 13553 13240
rect 13228 13200 13234 13212
rect 13541 13209 13553 13212
rect 13587 13240 13599 13243
rect 15381 13243 15439 13249
rect 13587 13212 15332 13240
rect 13587 13209 13599 13212
rect 13541 13203 13599 13209
rect 11839 13144 12848 13172
rect 14737 13175 14795 13181
rect 11839 13141 11851 13144
rect 11793 13135 11851 13141
rect 14737 13141 14749 13175
rect 14783 13172 14795 13175
rect 14826 13172 14832 13184
rect 14783 13144 14832 13172
rect 14783 13141 14795 13144
rect 14737 13135 14795 13141
rect 14826 13132 14832 13144
rect 14884 13132 14890 13184
rect 15304 13172 15332 13212
rect 15381 13209 15393 13243
rect 15427 13240 15439 13243
rect 15930 13240 15936 13252
rect 15427 13212 15936 13240
rect 15427 13209 15439 13212
rect 15381 13203 15439 13209
rect 15930 13200 15936 13212
rect 15988 13240 15994 13252
rect 16209 13243 16267 13249
rect 16209 13240 16221 13243
rect 15988 13212 16221 13240
rect 15988 13200 15994 13212
rect 16209 13209 16221 13212
rect 16255 13209 16267 13243
rect 16209 13203 16267 13209
rect 16298 13200 16304 13252
rect 16356 13240 16362 13252
rect 17770 13240 17776 13252
rect 16356 13212 16401 13240
rect 16500 13212 16804 13240
rect 17731 13212 17776 13240
rect 16356 13200 16362 13212
rect 16500 13172 16528 13212
rect 15304 13144 16528 13172
rect 16577 13175 16635 13181
rect 16577 13141 16589 13175
rect 16623 13172 16635 13175
rect 16666 13172 16672 13184
rect 16623 13144 16672 13172
rect 16623 13141 16635 13144
rect 16577 13135 16635 13141
rect 16666 13132 16672 13144
rect 16724 13132 16730 13184
rect 16776 13172 16804 13212
rect 17770 13200 17776 13212
rect 17828 13200 17834 13252
rect 17972 13172 18000 13348
rect 21358 13336 21364 13348
rect 21416 13336 21422 13388
rect 23106 13336 23112 13388
rect 23164 13376 23170 13388
rect 23201 13379 23259 13385
rect 23201 13376 23213 13379
rect 23164 13348 23213 13376
rect 23164 13336 23170 13348
rect 23201 13345 23213 13348
rect 23247 13345 23259 13379
rect 23201 13339 23259 13345
rect 23293 13379 23351 13385
rect 23293 13345 23305 13379
rect 23339 13345 23351 13379
rect 23293 13339 23351 13345
rect 19245 13311 19303 13317
rect 19245 13277 19257 13311
rect 19291 13277 19303 13311
rect 19245 13271 19303 13277
rect 16776 13144 18000 13172
rect 18049 13175 18107 13181
rect 18049 13141 18061 13175
rect 18095 13172 18107 13175
rect 19260 13172 19288 13271
rect 19334 13268 19340 13320
rect 19392 13308 19398 13320
rect 19705 13311 19763 13317
rect 19705 13308 19717 13311
rect 19392 13280 19717 13308
rect 19392 13268 19398 13280
rect 19705 13277 19717 13280
rect 19751 13277 19763 13311
rect 19705 13271 19763 13277
rect 20530 13268 20536 13320
rect 20588 13308 20594 13320
rect 20625 13311 20683 13317
rect 20625 13308 20637 13311
rect 20588 13280 20637 13308
rect 20588 13268 20594 13280
rect 20625 13277 20637 13280
rect 20671 13277 20683 13311
rect 22094 13308 22100 13320
rect 22055 13280 22100 13308
rect 20625 13271 20683 13277
rect 22094 13268 22100 13280
rect 22152 13268 22158 13320
rect 23014 13268 23020 13320
rect 23072 13308 23078 13320
rect 23308 13308 23336 13339
rect 23072 13280 23336 13308
rect 23072 13268 23078 13280
rect 19978 13240 19984 13252
rect 19939 13212 19984 13240
rect 19978 13200 19984 13212
rect 20036 13200 20042 13252
rect 20346 13200 20352 13252
rect 20404 13240 20410 13252
rect 20441 13243 20499 13249
rect 20441 13240 20453 13243
rect 20404 13212 20453 13240
rect 20404 13200 20410 13212
rect 20441 13209 20453 13212
rect 20487 13209 20499 13243
rect 20441 13203 20499 13209
rect 22646 13200 22652 13252
rect 22704 13240 22710 13252
rect 23290 13240 23296 13252
rect 22704 13212 23296 13240
rect 22704 13200 22710 13212
rect 23290 13200 23296 13212
rect 23348 13200 23354 13252
rect 18095 13144 19288 13172
rect 22005 13175 22063 13181
rect 18095 13141 18107 13144
rect 18049 13135 18107 13141
rect 22005 13141 22017 13175
rect 22051 13172 22063 13175
rect 22094 13172 22100 13184
rect 22051 13144 22100 13172
rect 22051 13141 22063 13144
rect 22005 13135 22063 13141
rect 22094 13132 22100 13144
rect 22152 13132 22158 13184
rect 24044 13172 24072 13484
rect 24118 13472 24124 13524
rect 24176 13512 24182 13524
rect 28077 13515 28135 13521
rect 24176 13484 26372 13512
rect 24176 13472 24182 13484
rect 25501 13447 25559 13453
rect 25501 13413 25513 13447
rect 25547 13413 25559 13447
rect 25501 13407 25559 13413
rect 25516 13376 25544 13407
rect 26145 13379 26203 13385
rect 26145 13376 26157 13379
rect 25516 13348 26157 13376
rect 26145 13345 26157 13348
rect 26191 13345 26203 13379
rect 26344 13376 26372 13484
rect 28077 13481 28089 13515
rect 28123 13512 28135 13515
rect 30926 13512 30932 13524
rect 28123 13484 30932 13512
rect 28123 13481 28135 13484
rect 28077 13475 28135 13481
rect 30926 13472 30932 13484
rect 30984 13472 30990 13524
rect 31110 13512 31116 13524
rect 31071 13484 31116 13512
rect 31110 13472 31116 13484
rect 31168 13472 31174 13524
rect 31202 13472 31208 13524
rect 31260 13512 31266 13524
rect 53190 13512 53196 13524
rect 31260 13484 35572 13512
rect 53151 13484 53196 13512
rect 31260 13472 31266 13484
rect 29825 13447 29883 13453
rect 29825 13413 29837 13447
rect 29871 13444 29883 13447
rect 35544 13444 35572 13484
rect 53190 13472 53196 13484
rect 53248 13472 53254 13524
rect 56594 13472 56600 13524
rect 56652 13512 56658 13524
rect 56781 13515 56839 13521
rect 56781 13512 56793 13515
rect 56652 13484 56793 13512
rect 56652 13472 56658 13484
rect 56781 13481 56793 13484
rect 56827 13481 56839 13515
rect 56781 13475 56839 13481
rect 57149 13515 57207 13521
rect 57149 13481 57161 13515
rect 57195 13512 57207 13515
rect 57882 13512 57888 13524
rect 57195 13484 57888 13512
rect 57195 13481 57207 13484
rect 57149 13475 57207 13481
rect 57882 13472 57888 13484
rect 57940 13472 57946 13524
rect 57790 13444 57796 13456
rect 29871 13416 35480 13444
rect 35544 13416 57796 13444
rect 29871 13413 29883 13416
rect 29825 13407 29883 13413
rect 35345 13379 35403 13385
rect 35345 13376 35357 13379
rect 26344 13348 35357 13376
rect 26145 13339 26203 13345
rect 35345 13345 35357 13348
rect 35391 13345 35403 13379
rect 35345 13339 35403 13345
rect 24854 13308 24860 13320
rect 24815 13280 24860 13308
rect 24854 13268 24860 13280
rect 24912 13268 24918 13320
rect 24950 13311 25008 13317
rect 24950 13277 24962 13311
rect 24996 13308 25008 13311
rect 25038 13308 25044 13320
rect 24996 13280 25044 13308
rect 24996 13277 25008 13280
rect 24950 13271 25008 13277
rect 25038 13268 25044 13280
rect 25096 13268 25102 13320
rect 25222 13308 25228 13320
rect 25183 13280 25228 13308
rect 25222 13268 25228 13280
rect 25280 13268 25286 13320
rect 25363 13311 25421 13317
rect 25363 13277 25375 13311
rect 25409 13308 25421 13311
rect 25590 13308 25596 13320
rect 25409 13280 25596 13308
rect 25409 13277 25421 13280
rect 25363 13271 25421 13277
rect 25590 13268 25596 13280
rect 25648 13268 25654 13320
rect 26234 13308 26240 13320
rect 26195 13280 26240 13308
rect 26234 13268 26240 13280
rect 26292 13268 26298 13320
rect 27798 13308 27804 13320
rect 27759 13280 27804 13308
rect 27798 13268 27804 13280
rect 27856 13268 27862 13320
rect 27982 13268 27988 13320
rect 28040 13308 28046 13320
rect 28077 13311 28135 13317
rect 28077 13308 28089 13311
rect 28040 13280 28089 13308
rect 28040 13268 28046 13280
rect 28077 13277 28089 13280
rect 28123 13277 28135 13311
rect 28077 13271 28135 13277
rect 29638 13268 29644 13320
rect 29696 13308 29702 13320
rect 29825 13311 29883 13317
rect 29825 13308 29837 13311
rect 29696 13280 29837 13308
rect 29696 13268 29702 13280
rect 29825 13277 29837 13280
rect 29871 13277 29883 13311
rect 29825 13271 29883 13277
rect 30006 13268 30012 13320
rect 30064 13308 30070 13320
rect 30101 13311 30159 13317
rect 30101 13308 30113 13311
rect 30064 13280 30113 13308
rect 30064 13268 30070 13280
rect 30101 13277 30113 13280
rect 30147 13308 30159 13311
rect 30190 13308 30196 13320
rect 30147 13280 30196 13308
rect 30147 13277 30159 13280
rect 30101 13271 30159 13277
rect 30190 13268 30196 13280
rect 30248 13268 30254 13320
rect 32030 13268 32036 13320
rect 32088 13308 32094 13320
rect 32217 13311 32275 13317
rect 32217 13308 32229 13311
rect 32088 13280 32229 13308
rect 32088 13268 32094 13280
rect 32217 13277 32229 13280
rect 32263 13277 32275 13311
rect 32217 13271 32275 13277
rect 32493 13311 32551 13317
rect 32493 13277 32505 13311
rect 32539 13308 32551 13311
rect 32582 13308 32588 13320
rect 32539 13280 32588 13308
rect 32539 13277 32551 13280
rect 32493 13271 32551 13277
rect 32582 13268 32588 13280
rect 32640 13268 32646 13320
rect 24118 13200 24124 13252
rect 24176 13240 24182 13252
rect 25130 13240 25136 13252
rect 24176 13212 25136 13240
rect 24176 13200 24182 13212
rect 25130 13200 25136 13212
rect 25188 13200 25194 13252
rect 28718 13240 28724 13252
rect 25240 13212 28724 13240
rect 25240 13172 25268 13212
rect 28718 13200 28724 13212
rect 28776 13200 28782 13252
rect 32122 13200 32128 13252
rect 32180 13240 32186 13252
rect 32306 13240 32312 13252
rect 32180 13212 32312 13240
rect 32180 13200 32186 13212
rect 32306 13200 32312 13212
rect 32364 13200 32370 13252
rect 35452 13240 35480 13416
rect 57790 13404 57796 13416
rect 57848 13404 57854 13456
rect 36265 13379 36323 13385
rect 36265 13345 36277 13379
rect 36311 13376 36323 13379
rect 40681 13379 40739 13385
rect 40681 13376 40693 13379
rect 36311 13348 40693 13376
rect 36311 13345 36323 13348
rect 36265 13339 36323 13345
rect 40681 13345 40693 13348
rect 40727 13376 40739 13379
rect 41138 13376 41144 13388
rect 40727 13348 41144 13376
rect 40727 13345 40739 13348
rect 40681 13339 40739 13345
rect 41138 13336 41144 13348
rect 41196 13336 41202 13388
rect 46750 13376 46756 13388
rect 46711 13348 46756 13376
rect 46750 13336 46756 13348
rect 46808 13336 46814 13388
rect 50706 13376 50712 13388
rect 50667 13348 50712 13376
rect 50706 13336 50712 13348
rect 50764 13336 50770 13388
rect 56870 13376 56876 13388
rect 56831 13348 56876 13376
rect 56870 13336 56876 13348
rect 56928 13336 56934 13388
rect 35621 13311 35679 13317
rect 35621 13277 35633 13311
rect 35667 13308 35679 13311
rect 36170 13308 36176 13320
rect 35667 13280 36176 13308
rect 35667 13277 35679 13280
rect 35621 13271 35679 13277
rect 36170 13268 36176 13280
rect 36228 13268 36234 13320
rect 40770 13308 40776 13320
rect 40731 13280 40776 13308
rect 40770 13268 40776 13280
rect 40828 13268 40834 13320
rect 42334 13308 42340 13320
rect 42295 13280 42340 13308
rect 42334 13268 42340 13280
rect 42392 13268 42398 13320
rect 42521 13311 42579 13317
rect 42521 13277 42533 13311
rect 42567 13277 42579 13311
rect 45002 13308 45008 13320
rect 44963 13280 45008 13308
rect 42521 13271 42579 13277
rect 37734 13240 37740 13252
rect 35452 13212 37740 13240
rect 37734 13200 37740 13212
rect 37792 13200 37798 13252
rect 42536 13240 42564 13271
rect 45002 13268 45008 13280
rect 45060 13268 45066 13320
rect 45094 13268 45100 13320
rect 45152 13308 45158 13320
rect 45152 13280 45197 13308
rect 45152 13268 45158 13280
rect 45278 13268 45284 13320
rect 45336 13308 45342 13320
rect 46934 13308 46940 13320
rect 45336 13280 45381 13308
rect 46895 13280 46940 13308
rect 45336 13268 45342 13280
rect 46934 13268 46940 13280
rect 46992 13268 46998 13320
rect 48314 13308 48320 13320
rect 48275 13280 48320 13308
rect 48314 13268 48320 13280
rect 48372 13268 48378 13320
rect 50798 13308 50804 13320
rect 42886 13240 42892 13252
rect 41386 13212 42892 13240
rect 27062 13172 27068 13184
rect 24044 13144 25268 13172
rect 27023 13144 27068 13172
rect 27062 13132 27068 13144
rect 27120 13132 27126 13184
rect 27246 13132 27252 13184
rect 27304 13172 27310 13184
rect 27893 13175 27951 13181
rect 27893 13172 27905 13175
rect 27304 13144 27905 13172
rect 27304 13132 27310 13144
rect 27893 13141 27905 13144
rect 27939 13172 27951 13175
rect 28537 13175 28595 13181
rect 28537 13172 28549 13175
rect 27939 13144 28549 13172
rect 27939 13141 27951 13144
rect 27893 13135 27951 13141
rect 28537 13141 28549 13144
rect 28583 13141 28595 13175
rect 28537 13135 28595 13141
rect 29362 13132 29368 13184
rect 29420 13172 29426 13184
rect 30009 13175 30067 13181
rect 30009 13172 30021 13175
rect 29420 13144 30021 13172
rect 29420 13132 29426 13144
rect 30009 13141 30021 13144
rect 30055 13141 30067 13175
rect 30009 13135 30067 13141
rect 31754 13132 31760 13184
rect 31812 13172 31818 13184
rect 32490 13172 32496 13184
rect 31812 13144 32496 13172
rect 31812 13132 31818 13144
rect 32490 13132 32496 13144
rect 32548 13132 32554 13184
rect 32677 13175 32735 13181
rect 32677 13141 32689 13175
rect 32723 13172 32735 13175
rect 34790 13172 34796 13184
rect 32723 13144 34796 13172
rect 32723 13141 32735 13144
rect 32677 13135 32735 13141
rect 34790 13132 34796 13144
rect 34848 13132 34854 13184
rect 37550 13132 37556 13184
rect 37608 13172 37614 13184
rect 38470 13172 38476 13184
rect 37608 13144 38476 13172
rect 37608 13132 37614 13144
rect 38470 13132 38476 13144
rect 38528 13132 38534 13184
rect 41141 13175 41199 13181
rect 41141 13141 41153 13175
rect 41187 13172 41199 13175
rect 41386 13172 41414 13212
rect 42886 13200 42892 13212
rect 42944 13200 42950 13252
rect 47673 13243 47731 13249
rect 47673 13209 47685 13243
rect 47719 13240 47731 13243
rect 47946 13240 47952 13252
rect 47719 13212 47952 13240
rect 47719 13209 47731 13212
rect 47673 13203 47731 13209
rect 47946 13200 47952 13212
rect 48004 13240 48010 13252
rect 48424 13240 48452 13294
rect 50759 13280 50804 13308
rect 50798 13268 50804 13280
rect 50856 13268 50862 13320
rect 53006 13308 53012 13320
rect 52919 13280 53012 13308
rect 53006 13268 53012 13280
rect 53064 13268 53070 13320
rect 56778 13308 56784 13320
rect 56739 13280 56784 13308
rect 56778 13268 56784 13280
rect 56836 13268 56842 13320
rect 48004 13212 48452 13240
rect 49329 13243 49387 13249
rect 48004 13200 48010 13212
rect 49329 13209 49341 13243
rect 49375 13240 49387 13243
rect 53024 13240 53052 13268
rect 49375 13212 53052 13240
rect 49375 13209 49387 13212
rect 49329 13203 49387 13209
rect 43346 13172 43352 13184
rect 41187 13144 41414 13172
rect 43307 13144 43352 13172
rect 41187 13141 41199 13144
rect 41141 13135 41199 13141
rect 43346 13132 43352 13144
rect 43404 13132 43410 13184
rect 45462 13172 45468 13184
rect 45423 13144 45468 13172
rect 45462 13132 45468 13144
rect 45520 13132 45526 13184
rect 51166 13172 51172 13184
rect 51127 13144 51172 13172
rect 51166 13132 51172 13144
rect 51224 13132 51230 13184
rect 53469 13175 53527 13181
rect 53469 13141 53481 13175
rect 53515 13172 53527 13175
rect 54478 13172 54484 13184
rect 53515 13144 54484 13172
rect 53515 13141 53527 13144
rect 53469 13135 53527 13141
rect 54478 13132 54484 13144
rect 54536 13132 54542 13184
rect 1104 13082 58880 13104
rect 1104 13030 19574 13082
rect 19626 13030 19638 13082
rect 19690 13030 19702 13082
rect 19754 13030 19766 13082
rect 19818 13030 19830 13082
rect 19882 13030 50294 13082
rect 50346 13030 50358 13082
rect 50410 13030 50422 13082
rect 50474 13030 50486 13082
rect 50538 13030 50550 13082
rect 50602 13030 58880 13082
rect 1104 13008 58880 13030
rect 1578 12968 1584 12980
rect 1539 12940 1584 12968
rect 1578 12928 1584 12940
rect 1636 12928 1642 12980
rect 10413 12971 10471 12977
rect 10413 12937 10425 12971
rect 10459 12968 10471 12971
rect 10962 12968 10968 12980
rect 10459 12940 10968 12968
rect 10459 12937 10471 12940
rect 10413 12931 10471 12937
rect 3050 12860 3056 12912
rect 3108 12900 3114 12912
rect 3234 12900 3240 12912
rect 3108 12872 3240 12900
rect 3108 12860 3114 12872
rect 3234 12860 3240 12872
rect 3292 12900 3298 12912
rect 6362 12900 6368 12912
rect 3292 12872 4200 12900
rect 6323 12872 6368 12900
rect 3292 12860 3298 12872
rect 1394 12832 1400 12844
rect 1355 12804 1400 12832
rect 1394 12792 1400 12804
rect 1452 12792 1458 12844
rect 2866 12792 2872 12844
rect 2924 12832 2930 12844
rect 3145 12835 3203 12841
rect 3145 12832 3157 12835
rect 2924 12804 3157 12832
rect 2924 12792 2930 12804
rect 3145 12801 3157 12804
rect 3191 12801 3203 12835
rect 3145 12795 3203 12801
rect 4065 12835 4123 12841
rect 4065 12801 4077 12835
rect 4111 12801 4123 12835
rect 4065 12795 4123 12801
rect 2590 12764 2596 12776
rect 2551 12736 2596 12764
rect 2590 12724 2596 12736
rect 2648 12724 2654 12776
rect 3050 12588 3056 12640
rect 3108 12628 3114 12640
rect 4080 12628 4108 12795
rect 4172 12764 4200 12872
rect 6362 12860 6368 12872
rect 6420 12860 6426 12912
rect 9674 12900 9680 12912
rect 9508 12872 9680 12900
rect 6546 12832 6552 12844
rect 6507 12804 6552 12832
rect 6546 12792 6552 12804
rect 6604 12792 6610 12844
rect 6733 12835 6791 12841
rect 6733 12801 6745 12835
rect 6779 12832 6791 12835
rect 7282 12832 7288 12844
rect 6779 12804 7288 12832
rect 6779 12801 6791 12804
rect 6733 12795 6791 12801
rect 7282 12792 7288 12804
rect 7340 12792 7346 12844
rect 8573 12835 8631 12841
rect 8573 12801 8585 12835
rect 8619 12832 8631 12835
rect 8662 12832 8668 12844
rect 8619 12804 8668 12832
rect 8619 12801 8631 12804
rect 8573 12795 8631 12801
rect 8662 12792 8668 12804
rect 8720 12792 8726 12844
rect 8846 12832 8852 12844
rect 8807 12804 8852 12832
rect 8846 12792 8852 12804
rect 8904 12792 8910 12844
rect 9508 12841 9536 12872
rect 9674 12860 9680 12872
rect 9732 12860 9738 12912
rect 9493 12835 9551 12841
rect 9493 12801 9505 12835
rect 9539 12801 9551 12835
rect 9493 12795 9551 12801
rect 9861 12835 9919 12841
rect 9861 12801 9873 12835
rect 9907 12832 9919 12835
rect 10428 12832 10456 12931
rect 10962 12928 10968 12940
rect 11020 12928 11026 12980
rect 13078 12968 13084 12980
rect 13039 12940 13084 12968
rect 13078 12928 13084 12940
rect 13136 12928 13142 12980
rect 14918 12968 14924 12980
rect 14879 12940 14924 12968
rect 14918 12928 14924 12940
rect 14976 12968 14982 12980
rect 15102 12968 15108 12980
rect 14976 12940 15108 12968
rect 14976 12928 14982 12940
rect 15102 12928 15108 12940
rect 15160 12928 15166 12980
rect 16945 12971 17003 12977
rect 16945 12937 16957 12971
rect 16991 12968 17003 12971
rect 19153 12971 19211 12977
rect 16991 12940 19104 12968
rect 16991 12937 17003 12940
rect 16945 12931 17003 12937
rect 13633 12903 13691 12909
rect 13633 12900 13645 12903
rect 12406 12872 13645 12900
rect 9907 12804 10456 12832
rect 9907 12801 9919 12804
rect 9861 12795 9919 12801
rect 11974 12792 11980 12844
rect 12032 12832 12038 12844
rect 12069 12835 12127 12841
rect 12069 12832 12081 12835
rect 12032 12804 12081 12832
rect 12032 12792 12038 12804
rect 12069 12801 12081 12804
rect 12115 12832 12127 12835
rect 12406 12832 12434 12872
rect 13633 12869 13645 12872
rect 13679 12869 13691 12903
rect 13633 12863 13691 12869
rect 14277 12903 14335 12909
rect 14277 12869 14289 12903
rect 14323 12900 14335 12903
rect 15654 12900 15660 12912
rect 14323 12872 15660 12900
rect 14323 12869 14335 12872
rect 14277 12863 14335 12869
rect 15654 12860 15660 12872
rect 15712 12860 15718 12912
rect 16114 12860 16120 12912
rect 16172 12900 16178 12912
rect 16172 12872 16896 12900
rect 16172 12860 16178 12872
rect 12115 12804 12434 12832
rect 12115 12801 12127 12804
rect 12069 12795 12127 12801
rect 12710 12792 12716 12844
rect 12768 12832 12774 12844
rect 12989 12835 13047 12841
rect 12989 12832 13001 12835
rect 12768 12804 13001 12832
rect 12768 12792 12774 12804
rect 12989 12801 13001 12804
rect 13035 12801 13047 12835
rect 13170 12832 13176 12844
rect 13131 12804 13176 12832
rect 12989 12795 13047 12801
rect 13170 12792 13176 12804
rect 13228 12792 13234 12844
rect 14734 12792 14740 12844
rect 14792 12832 14798 12844
rect 15473 12835 15531 12841
rect 15473 12832 15485 12835
rect 14792 12804 15485 12832
rect 14792 12792 14798 12804
rect 15473 12801 15485 12804
rect 15519 12832 15531 12835
rect 15838 12832 15844 12844
rect 15519 12804 15844 12832
rect 15519 12801 15531 12804
rect 15473 12795 15531 12801
rect 15838 12792 15844 12804
rect 15896 12792 15902 12844
rect 16666 12832 16672 12844
rect 16627 12804 16672 12832
rect 16666 12792 16672 12804
rect 16724 12792 16730 12844
rect 16868 12841 16896 12872
rect 17770 12860 17776 12912
rect 17828 12900 17834 12912
rect 18785 12903 18843 12909
rect 18785 12900 18797 12903
rect 17828 12872 18797 12900
rect 17828 12860 17834 12872
rect 18785 12869 18797 12872
rect 18831 12869 18843 12903
rect 19076 12900 19104 12940
rect 19153 12937 19165 12971
rect 19199 12968 19211 12971
rect 19334 12968 19340 12980
rect 19199 12940 19340 12968
rect 19199 12937 19211 12940
rect 19153 12931 19211 12937
rect 19334 12928 19340 12940
rect 19392 12928 19398 12980
rect 19426 12928 19432 12980
rect 19484 12968 19490 12980
rect 19705 12971 19763 12977
rect 19705 12968 19717 12971
rect 19484 12940 19717 12968
rect 19484 12928 19490 12940
rect 19705 12937 19717 12940
rect 19751 12968 19763 12971
rect 20070 12968 20076 12980
rect 19751 12940 20076 12968
rect 19751 12937 19763 12940
rect 19705 12931 19763 12937
rect 20070 12928 20076 12940
rect 20128 12928 20134 12980
rect 23290 12928 23296 12980
rect 23348 12968 23354 12980
rect 23937 12971 23995 12977
rect 23937 12968 23949 12971
rect 23348 12940 23949 12968
rect 23348 12928 23354 12940
rect 23937 12937 23949 12940
rect 23983 12937 23995 12971
rect 23937 12931 23995 12937
rect 24412 12940 24808 12968
rect 24026 12900 24032 12912
rect 19076 12872 24032 12900
rect 18785 12863 18843 12869
rect 24026 12860 24032 12872
rect 24084 12860 24090 12912
rect 16853 12835 16911 12841
rect 16853 12801 16865 12835
rect 16899 12801 16911 12835
rect 16853 12795 16911 12801
rect 17954 12792 17960 12844
rect 18012 12832 18018 12844
rect 18601 12835 18659 12841
rect 18601 12832 18613 12835
rect 18012 12804 18613 12832
rect 18012 12792 18018 12804
rect 18601 12801 18613 12804
rect 18647 12801 18659 12835
rect 18874 12832 18880 12844
rect 18835 12804 18880 12832
rect 18601 12795 18659 12801
rect 18874 12792 18880 12804
rect 18932 12792 18938 12844
rect 18969 12835 19027 12841
rect 18969 12801 18981 12835
rect 19015 12801 19027 12835
rect 18969 12795 19027 12801
rect 8389 12767 8447 12773
rect 8389 12764 8401 12767
rect 4172 12736 8401 12764
rect 8389 12733 8401 12736
rect 8435 12733 8447 12767
rect 8389 12727 8447 12733
rect 12345 12767 12403 12773
rect 12345 12733 12357 12767
rect 12391 12764 12403 12767
rect 12434 12764 12440 12776
rect 12391 12736 12440 12764
rect 12391 12733 12403 12736
rect 12345 12727 12403 12733
rect 12434 12724 12440 12736
rect 12492 12724 12498 12776
rect 16022 12724 16028 12776
rect 16080 12764 16086 12776
rect 17034 12764 17040 12776
rect 16080 12736 17040 12764
rect 16080 12724 16086 12736
rect 17034 12724 17040 12736
rect 17092 12724 17098 12776
rect 18506 12724 18512 12776
rect 18564 12764 18570 12776
rect 18984 12764 19012 12795
rect 20070 12792 20076 12844
rect 20128 12832 20134 12844
rect 24412 12832 24440 12940
rect 24670 12900 24676 12912
rect 24631 12872 24676 12900
rect 24670 12860 24676 12872
rect 24728 12860 24734 12912
rect 24780 12900 24808 12940
rect 24854 12928 24860 12980
rect 24912 12968 24918 12980
rect 25041 12971 25099 12977
rect 25041 12968 25053 12971
rect 24912 12940 25053 12968
rect 24912 12928 24918 12940
rect 25041 12937 25053 12940
rect 25087 12937 25099 12971
rect 25041 12931 25099 12937
rect 27062 12928 27068 12980
rect 27120 12968 27126 12980
rect 37182 12968 37188 12980
rect 27120 12940 37188 12968
rect 27120 12928 27126 12940
rect 37182 12928 37188 12940
rect 37240 12928 37246 12980
rect 37550 12928 37556 12980
rect 37608 12968 37614 12980
rect 37829 12971 37887 12977
rect 37829 12968 37841 12971
rect 37608 12940 37841 12968
rect 37608 12928 37614 12940
rect 37829 12937 37841 12940
rect 37875 12937 37887 12971
rect 37829 12931 37887 12937
rect 43346 12928 43352 12980
rect 43404 12968 43410 12980
rect 48314 12968 48320 12980
rect 43404 12940 48320 12968
rect 43404 12928 43410 12940
rect 38746 12900 38752 12912
rect 24780 12872 31754 12900
rect 20128 12804 24440 12832
rect 20128 12792 20134 12804
rect 24486 12792 24492 12844
rect 24544 12832 24550 12844
rect 24762 12832 24768 12844
rect 24544 12804 24589 12832
rect 24723 12804 24768 12832
rect 24544 12792 24550 12804
rect 24762 12792 24768 12804
rect 24820 12792 24826 12844
rect 24857 12835 24915 12841
rect 24857 12801 24869 12835
rect 24903 12832 24915 12835
rect 24946 12832 24952 12844
rect 24903 12804 24952 12832
rect 24903 12801 24915 12804
rect 24857 12795 24915 12801
rect 24946 12792 24952 12804
rect 25004 12792 25010 12844
rect 25590 12832 25596 12844
rect 25551 12804 25596 12832
rect 25590 12792 25596 12804
rect 25648 12792 25654 12844
rect 28534 12792 28540 12844
rect 28592 12832 28598 12844
rect 28629 12835 28687 12841
rect 28629 12832 28641 12835
rect 28592 12804 28641 12832
rect 28592 12792 28598 12804
rect 28629 12801 28641 12804
rect 28675 12801 28687 12835
rect 28629 12795 28687 12801
rect 29178 12792 29184 12844
rect 29236 12832 29242 12844
rect 29362 12832 29368 12844
rect 29236 12804 29368 12832
rect 29236 12792 29242 12804
rect 29362 12792 29368 12804
rect 29420 12792 29426 12844
rect 30558 12832 30564 12844
rect 30519 12804 30564 12832
rect 30558 12792 30564 12804
rect 30616 12792 30622 12844
rect 20346 12764 20352 12776
rect 18564 12736 19012 12764
rect 19444 12736 20352 12764
rect 18564 12724 18570 12736
rect 17052 12696 17080 12724
rect 19444 12696 19472 12736
rect 20346 12724 20352 12736
rect 20404 12724 20410 12776
rect 25038 12724 25044 12776
rect 25096 12764 25102 12776
rect 27430 12764 27436 12776
rect 25096 12736 27436 12764
rect 25096 12724 25102 12736
rect 27430 12724 27436 12736
rect 27488 12724 27494 12776
rect 28166 12724 28172 12776
rect 28224 12764 28230 12776
rect 28353 12767 28411 12773
rect 28353 12764 28365 12767
rect 28224 12736 28365 12764
rect 28224 12724 28230 12736
rect 28353 12733 28365 12736
rect 28399 12733 28411 12767
rect 28353 12727 28411 12733
rect 28810 12724 28816 12776
rect 28868 12764 28874 12776
rect 29089 12767 29147 12773
rect 29089 12764 29101 12767
rect 28868 12736 29101 12764
rect 28868 12724 28874 12736
rect 29089 12733 29101 12736
rect 29135 12733 29147 12767
rect 31726 12764 31754 12872
rect 36740 12872 38752 12900
rect 32030 12792 32036 12844
rect 32088 12832 32094 12844
rect 32125 12835 32183 12841
rect 32125 12832 32137 12835
rect 32088 12804 32137 12832
rect 32088 12792 32094 12804
rect 32125 12801 32137 12804
rect 32171 12801 32183 12835
rect 32306 12832 32312 12844
rect 32267 12804 32312 12832
rect 32125 12795 32183 12801
rect 32306 12792 32312 12804
rect 32364 12792 32370 12844
rect 36740 12841 36768 12872
rect 36725 12835 36783 12841
rect 36725 12801 36737 12835
rect 36771 12801 36783 12835
rect 37734 12832 37740 12844
rect 37695 12804 37740 12832
rect 36725 12795 36783 12801
rect 37734 12792 37740 12804
rect 37792 12792 37798 12844
rect 38028 12841 38056 12872
rect 38746 12860 38752 12872
rect 38804 12900 38810 12912
rect 42886 12900 42892 12912
rect 38804 12872 38976 12900
rect 42847 12872 42892 12900
rect 38804 12860 38810 12872
rect 38948 12841 38976 12872
rect 42886 12860 42892 12872
rect 42944 12860 42950 12912
rect 45094 12860 45100 12912
rect 45152 12900 45158 12912
rect 47872 12909 47900 12940
rect 48314 12928 48320 12940
rect 48372 12928 48378 12980
rect 50341 12971 50399 12977
rect 50341 12937 50353 12971
rect 50387 12968 50399 12971
rect 50706 12968 50712 12980
rect 50387 12940 50712 12968
rect 50387 12937 50399 12940
rect 50341 12931 50399 12937
rect 50706 12928 50712 12940
rect 50764 12928 50770 12980
rect 54478 12968 54484 12980
rect 54439 12940 54484 12968
rect 54478 12928 54484 12940
rect 54536 12928 54542 12980
rect 55030 12968 55036 12980
rect 54588 12940 55036 12968
rect 46661 12903 46719 12909
rect 45152 12872 45232 12900
rect 45152 12860 45158 12872
rect 38013 12835 38071 12841
rect 38013 12801 38025 12835
rect 38059 12801 38071 12835
rect 38013 12795 38071 12801
rect 38657 12835 38715 12841
rect 38657 12801 38669 12835
rect 38703 12801 38715 12835
rect 38841 12835 38899 12841
rect 38841 12832 38853 12835
rect 38657 12795 38715 12801
rect 38764 12804 38853 12832
rect 32490 12764 32496 12776
rect 31726 12736 32496 12764
rect 29089 12727 29147 12733
rect 32490 12724 32496 12736
rect 32548 12764 32554 12776
rect 32674 12764 32680 12776
rect 32548 12736 32680 12764
rect 32548 12724 32554 12736
rect 32674 12724 32680 12736
rect 32732 12724 32738 12776
rect 33134 12724 33140 12776
rect 33192 12764 33198 12776
rect 36449 12767 36507 12773
rect 36449 12764 36461 12767
rect 33192 12736 36461 12764
rect 33192 12724 33198 12736
rect 36449 12733 36461 12736
rect 36495 12733 36507 12767
rect 37752 12764 37780 12792
rect 38672 12764 38700 12795
rect 37752 12736 38700 12764
rect 36449 12727 36507 12733
rect 25774 12696 25780 12708
rect 17052 12668 19472 12696
rect 25735 12668 25780 12696
rect 25774 12656 25780 12668
rect 25832 12656 25838 12708
rect 29454 12656 29460 12708
rect 29512 12696 29518 12708
rect 32217 12699 32275 12705
rect 32217 12696 32229 12699
rect 29512 12668 32229 12696
rect 29512 12656 29518 12668
rect 32217 12665 32229 12668
rect 32263 12665 32275 12699
rect 32217 12659 32275 12665
rect 38470 12656 38476 12708
rect 38528 12696 38534 12708
rect 38764 12696 38792 12804
rect 38841 12801 38853 12804
rect 38887 12801 38899 12835
rect 38841 12795 38899 12801
rect 38933 12835 38991 12841
rect 38933 12801 38945 12835
rect 38979 12801 38991 12835
rect 38933 12795 38991 12801
rect 40770 12792 40776 12844
rect 40828 12832 40834 12844
rect 41325 12835 41383 12841
rect 41325 12832 41337 12835
rect 40828 12804 41337 12832
rect 40828 12792 40834 12804
rect 41325 12801 41337 12804
rect 41371 12801 41383 12835
rect 41325 12795 41383 12801
rect 41601 12835 41659 12841
rect 41601 12801 41613 12835
rect 41647 12832 41659 12835
rect 45002 12832 45008 12844
rect 41647 12804 43576 12832
rect 44963 12804 45008 12832
rect 41647 12801 41659 12804
rect 41601 12795 41659 12801
rect 41138 12764 41144 12776
rect 41099 12736 41144 12764
rect 41138 12724 41144 12736
rect 41196 12724 41202 12776
rect 41693 12767 41751 12773
rect 41693 12733 41705 12767
rect 41739 12764 41751 12767
rect 42429 12767 42487 12773
rect 42429 12764 42441 12767
rect 41739 12736 42441 12764
rect 41739 12733 41751 12736
rect 41693 12727 41751 12733
rect 42429 12733 42441 12736
rect 42475 12733 42487 12767
rect 42429 12727 42487 12733
rect 38528 12668 38792 12696
rect 38528 12656 38534 12668
rect 42334 12656 42340 12708
rect 42392 12696 42398 12708
rect 42521 12699 42579 12705
rect 42521 12696 42533 12699
rect 42392 12668 42533 12696
rect 42392 12656 42398 12668
rect 42521 12665 42533 12668
rect 42567 12665 42579 12699
rect 43548 12696 43576 12804
rect 45002 12792 45008 12804
rect 45060 12792 45066 12844
rect 45204 12841 45232 12872
rect 46661 12869 46673 12903
rect 46707 12900 46719 12903
rect 47765 12903 47823 12909
rect 47765 12900 47777 12903
rect 46707 12872 47777 12900
rect 46707 12869 46719 12872
rect 46661 12863 46719 12869
rect 47765 12869 47777 12872
rect 47811 12869 47823 12903
rect 47765 12863 47823 12869
rect 47857 12903 47915 12909
rect 47857 12869 47869 12903
rect 47903 12869 47915 12903
rect 50724 12900 50752 12928
rect 54588 12909 54616 12940
rect 55030 12928 55036 12940
rect 55088 12968 55094 12980
rect 55398 12968 55404 12980
rect 55088 12940 55404 12968
rect 55088 12928 55094 12940
rect 55398 12928 55404 12940
rect 55456 12928 55462 12980
rect 54573 12903 54631 12909
rect 50724 12872 51028 12900
rect 47857 12863 47915 12869
rect 45189 12835 45247 12841
rect 45189 12801 45201 12835
rect 45235 12801 45247 12835
rect 45189 12795 45247 12801
rect 45278 12792 45284 12844
rect 45336 12832 45342 12844
rect 46569 12835 46627 12841
rect 46569 12832 46581 12835
rect 45336 12804 46581 12832
rect 45336 12792 45342 12804
rect 46569 12801 46581 12804
rect 46615 12801 46627 12835
rect 46750 12832 46756 12844
rect 46711 12804 46756 12832
rect 46569 12795 46627 12801
rect 46750 12792 46756 12804
rect 46808 12792 46814 12844
rect 46842 12792 46848 12844
rect 46900 12832 46906 12844
rect 47581 12835 47639 12841
rect 47581 12832 47593 12835
rect 46900 12804 47593 12832
rect 46900 12792 46906 12804
rect 47581 12801 47593 12804
rect 47627 12801 47639 12835
rect 47581 12795 47639 12801
rect 47946 12792 47952 12844
rect 48004 12832 48010 12844
rect 50798 12832 50804 12844
rect 48004 12804 48049 12832
rect 50711 12804 50804 12832
rect 48004 12792 48010 12804
rect 50798 12792 50804 12804
rect 50856 12792 50862 12844
rect 51000 12841 51028 12872
rect 54573 12869 54585 12903
rect 54619 12869 54631 12903
rect 55677 12903 55735 12909
rect 54573 12863 54631 12869
rect 54680 12872 55628 12900
rect 50985 12835 51043 12841
rect 50985 12801 50997 12835
rect 51031 12801 51043 12835
rect 50985 12795 51043 12801
rect 51166 12792 51172 12844
rect 51224 12832 51230 12844
rect 51442 12832 51448 12844
rect 51224 12804 51448 12832
rect 51224 12792 51230 12804
rect 51442 12792 51448 12804
rect 51500 12832 51506 12844
rect 51905 12835 51963 12841
rect 51905 12832 51917 12835
rect 51500 12804 51917 12832
rect 51500 12792 51506 12804
rect 51905 12801 51917 12804
rect 51951 12801 51963 12835
rect 51905 12795 51963 12801
rect 54113 12835 54171 12841
rect 54113 12801 54125 12835
rect 54159 12832 54171 12835
rect 54680 12832 54708 12872
rect 54159 12804 54708 12832
rect 54159 12801 54171 12804
rect 54113 12795 54171 12801
rect 55030 12792 55036 12844
rect 55088 12832 55094 12844
rect 55217 12835 55275 12841
rect 55088 12804 55133 12832
rect 55088 12792 55094 12804
rect 55217 12801 55229 12835
rect 55263 12801 55275 12835
rect 55217 12795 55275 12801
rect 55309 12835 55367 12841
rect 55309 12801 55321 12835
rect 55355 12801 55367 12835
rect 55309 12795 55367 12801
rect 55401 12835 55459 12841
rect 55401 12801 55413 12835
rect 55447 12801 55459 12835
rect 55600 12832 55628 12872
rect 55677 12869 55689 12903
rect 55723 12900 55735 12903
rect 56778 12900 56784 12912
rect 55723 12872 56784 12900
rect 55723 12869 55735 12872
rect 55677 12863 55735 12869
rect 56321 12835 56379 12841
rect 56321 12832 56333 12835
rect 55600 12804 56333 12832
rect 55401 12795 55459 12801
rect 56321 12801 56333 12804
rect 56367 12832 56379 12835
rect 56594 12832 56600 12844
rect 56367 12804 56600 12832
rect 56367 12801 56379 12804
rect 56321 12795 56379 12801
rect 45097 12767 45155 12773
rect 45097 12733 45109 12767
rect 45143 12764 45155 12767
rect 46106 12764 46112 12776
rect 45143 12736 46112 12764
rect 45143 12733 45155 12736
rect 45097 12727 45155 12733
rect 46106 12724 46112 12736
rect 46164 12764 46170 12776
rect 46768 12764 46796 12792
rect 46164 12736 46796 12764
rect 46164 12724 46170 12736
rect 50816 12696 50844 12792
rect 51626 12764 51632 12776
rect 51587 12736 51632 12764
rect 51626 12724 51632 12736
rect 51684 12724 51690 12776
rect 52089 12767 52147 12773
rect 52089 12733 52101 12767
rect 52135 12764 52147 12767
rect 54205 12767 54263 12773
rect 54205 12764 54217 12767
rect 52135 12736 54217 12764
rect 52135 12733 52147 12736
rect 52089 12727 52147 12733
rect 54205 12733 54217 12736
rect 54251 12733 54263 12767
rect 54205 12727 54263 12733
rect 43548 12668 50844 12696
rect 51077 12699 51135 12705
rect 42521 12659 42579 12665
rect 51077 12665 51089 12699
rect 51123 12696 51135 12699
rect 52546 12696 52552 12708
rect 51123 12668 52552 12696
rect 51123 12665 51135 12668
rect 51077 12659 51135 12665
rect 52546 12656 52552 12668
rect 52604 12656 52610 12708
rect 54220 12696 54248 12727
rect 54478 12724 54484 12776
rect 54536 12764 54542 12776
rect 55232 12764 55260 12795
rect 54536 12736 55260 12764
rect 54536 12724 54542 12736
rect 55324 12696 55352 12795
rect 54220 12668 55352 12696
rect 5902 12628 5908 12640
rect 3108 12600 5908 12628
rect 3108 12588 3114 12600
rect 5902 12588 5908 12600
rect 5960 12588 5966 12640
rect 7834 12628 7840 12640
rect 7795 12600 7840 12628
rect 7834 12588 7840 12600
rect 7892 12588 7898 12640
rect 10870 12628 10876 12640
rect 10831 12600 10876 12628
rect 10870 12588 10876 12600
rect 10928 12588 10934 12640
rect 18141 12631 18199 12637
rect 18141 12597 18153 12631
rect 18187 12628 18199 12631
rect 18874 12628 18880 12640
rect 18187 12600 18880 12628
rect 18187 12597 18199 12600
rect 18141 12591 18199 12597
rect 18874 12588 18880 12600
rect 18932 12588 18938 12640
rect 23014 12628 23020 12640
rect 22975 12600 23020 12628
rect 23014 12588 23020 12600
rect 23072 12588 23078 12640
rect 30469 12631 30527 12637
rect 30469 12597 30481 12631
rect 30515 12628 30527 12631
rect 30650 12628 30656 12640
rect 30515 12600 30656 12628
rect 30515 12597 30527 12600
rect 30469 12591 30527 12597
rect 30650 12588 30656 12600
rect 30708 12588 30714 12640
rect 38197 12631 38255 12637
rect 38197 12597 38209 12631
rect 38243 12628 38255 12631
rect 38286 12628 38292 12640
rect 38243 12600 38292 12628
rect 38243 12597 38255 12600
rect 38197 12591 38255 12597
rect 38286 12588 38292 12600
rect 38344 12588 38350 12640
rect 38746 12628 38752 12640
rect 38707 12600 38752 12628
rect 38746 12588 38752 12600
rect 38804 12588 38810 12640
rect 48133 12631 48191 12637
rect 48133 12597 48145 12631
rect 48179 12628 48191 12631
rect 49050 12628 49056 12640
rect 48179 12600 49056 12628
rect 48179 12597 48191 12600
rect 48133 12591 48191 12597
rect 49050 12588 49056 12600
rect 49108 12588 49114 12640
rect 51718 12628 51724 12640
rect 51679 12600 51724 12628
rect 51718 12588 51724 12600
rect 51776 12588 51782 12640
rect 52454 12588 52460 12640
rect 52512 12628 52518 12640
rect 54297 12631 54355 12637
rect 54297 12628 54309 12631
rect 52512 12600 54309 12628
rect 52512 12588 52518 12600
rect 54297 12597 54309 12600
rect 54343 12628 54355 12631
rect 55416 12628 55444 12795
rect 56594 12792 56600 12804
rect 56652 12792 56658 12844
rect 56704 12841 56732 12872
rect 56778 12860 56784 12872
rect 56836 12860 56842 12912
rect 56689 12835 56747 12841
rect 56689 12801 56701 12835
rect 56735 12801 56747 12835
rect 56689 12795 56747 12801
rect 56870 12792 56876 12844
rect 56928 12832 56934 12844
rect 56965 12835 57023 12841
rect 56965 12832 56977 12835
rect 56928 12804 56977 12832
rect 56928 12792 56934 12804
rect 56965 12801 56977 12804
rect 57011 12801 57023 12835
rect 56965 12795 57023 12801
rect 56134 12724 56140 12776
rect 56192 12764 56198 12776
rect 56505 12767 56563 12773
rect 56505 12764 56517 12767
rect 56192 12736 56517 12764
rect 56192 12724 56198 12736
rect 56505 12733 56517 12736
rect 56551 12733 56563 12767
rect 56505 12727 56563 12733
rect 54343 12600 55444 12628
rect 54343 12597 54355 12600
rect 54297 12591 54355 12597
rect 1104 12538 58880 12560
rect 1104 12486 4214 12538
rect 4266 12486 4278 12538
rect 4330 12486 4342 12538
rect 4394 12486 4406 12538
rect 4458 12486 4470 12538
rect 4522 12486 34934 12538
rect 34986 12486 34998 12538
rect 35050 12486 35062 12538
rect 35114 12486 35126 12538
rect 35178 12486 35190 12538
rect 35242 12486 58880 12538
rect 1104 12464 58880 12486
rect 3142 12384 3148 12436
rect 3200 12424 3206 12436
rect 3789 12427 3847 12433
rect 3789 12424 3801 12427
rect 3200 12396 3801 12424
rect 3200 12384 3206 12396
rect 3789 12393 3801 12396
rect 3835 12393 3847 12427
rect 3789 12387 3847 12393
rect 4157 12427 4215 12433
rect 4157 12393 4169 12427
rect 4203 12424 4215 12427
rect 5902 12424 5908 12436
rect 4203 12396 5212 12424
rect 5863 12396 5908 12424
rect 4203 12393 4215 12396
rect 4157 12387 4215 12393
rect 1394 12356 1400 12368
rect 1355 12328 1400 12356
rect 1394 12316 1400 12328
rect 1452 12316 1458 12368
rect 4246 12220 4252 12232
rect 4207 12192 4252 12220
rect 4246 12180 4252 12192
rect 4304 12180 4310 12232
rect 5184 12229 5212 12396
rect 5902 12384 5908 12396
rect 5960 12384 5966 12436
rect 8662 12384 8668 12436
rect 8720 12424 8726 12436
rect 9125 12427 9183 12433
rect 9125 12424 9137 12427
rect 8720 12396 9137 12424
rect 8720 12384 8726 12396
rect 9125 12393 9137 12396
rect 9171 12393 9183 12427
rect 14461 12427 14519 12433
rect 14461 12424 14473 12427
rect 9125 12387 9183 12393
rect 13372 12396 14473 12424
rect 10410 12316 10416 12368
rect 10468 12356 10474 12368
rect 13372 12356 13400 12396
rect 14461 12393 14473 12396
rect 14507 12393 14519 12427
rect 14461 12387 14519 12393
rect 15933 12427 15991 12433
rect 15933 12393 15945 12427
rect 15979 12424 15991 12427
rect 17126 12424 17132 12436
rect 15979 12396 17132 12424
rect 15979 12393 15991 12396
rect 15933 12387 15991 12393
rect 10468 12328 13400 12356
rect 13449 12359 13507 12365
rect 10468 12316 10474 12328
rect 13449 12325 13461 12359
rect 13495 12356 13507 12359
rect 13538 12356 13544 12368
rect 13495 12328 13544 12356
rect 13495 12325 13507 12328
rect 13449 12319 13507 12325
rect 6546 12288 6552 12300
rect 5368 12260 6552 12288
rect 5368 12229 5396 12260
rect 6546 12248 6552 12260
rect 6604 12288 6610 12300
rect 8389 12291 8447 12297
rect 8389 12288 8401 12291
rect 6604 12260 8401 12288
rect 6604 12248 6610 12260
rect 8389 12257 8401 12260
rect 8435 12288 8447 12291
rect 8846 12288 8852 12300
rect 8435 12260 8852 12288
rect 8435 12257 8447 12260
rect 8389 12251 8447 12257
rect 8846 12248 8852 12260
rect 8904 12248 8910 12300
rect 12434 12248 12440 12300
rect 12492 12288 12498 12300
rect 13464 12288 13492 12319
rect 13538 12316 13544 12328
rect 13596 12316 13602 12368
rect 12492 12260 13492 12288
rect 12492 12248 12498 12260
rect 5169 12223 5227 12229
rect 5169 12189 5181 12223
rect 5215 12189 5227 12223
rect 5169 12183 5227 12189
rect 5353 12223 5411 12229
rect 5353 12189 5365 12223
rect 5399 12189 5411 12223
rect 5353 12183 5411 12189
rect 6084 12223 6142 12229
rect 6084 12189 6096 12223
rect 6130 12220 6142 12223
rect 6130 12192 6408 12220
rect 6130 12189 6142 12192
rect 6084 12183 6142 12189
rect 5184 12152 5212 12183
rect 5718 12152 5724 12164
rect 5184 12124 5724 12152
rect 5718 12112 5724 12124
rect 5776 12112 5782 12164
rect 6178 12152 6184 12164
rect 6139 12124 6184 12152
rect 6178 12112 6184 12124
rect 6236 12112 6242 12164
rect 6273 12155 6331 12161
rect 6273 12121 6285 12155
rect 6319 12121 6331 12155
rect 6380 12152 6408 12192
rect 6454 12180 6460 12232
rect 6512 12220 6518 12232
rect 7098 12220 7104 12232
rect 6512 12192 6557 12220
rect 7011 12192 7104 12220
rect 6512 12180 6518 12192
rect 7098 12180 7104 12192
rect 7156 12220 7162 12232
rect 8018 12220 8024 12232
rect 7156 12192 7788 12220
rect 7979 12192 8024 12220
rect 7156 12180 7162 12192
rect 6917 12155 6975 12161
rect 6917 12152 6929 12155
rect 6380 12124 6929 12152
rect 6273 12115 6331 12121
rect 6917 12121 6929 12124
rect 6963 12121 6975 12155
rect 7282 12152 7288 12164
rect 7243 12124 7288 12152
rect 6917 12115 6975 12121
rect 5261 12087 5319 12093
rect 5261 12053 5273 12087
rect 5307 12084 5319 12087
rect 6288 12084 6316 12115
rect 7282 12112 7288 12124
rect 7340 12112 7346 12164
rect 7760 12152 7788 12192
rect 8018 12180 8024 12192
rect 8076 12180 8082 12232
rect 8205 12223 8263 12229
rect 8205 12189 8217 12223
rect 8251 12220 8263 12223
rect 8938 12220 8944 12232
rect 8251 12192 8944 12220
rect 8251 12189 8263 12192
rect 8205 12183 8263 12189
rect 8938 12180 8944 12192
rect 8996 12220 9002 12232
rect 9309 12223 9367 12229
rect 9309 12220 9321 12223
rect 8996 12192 9321 12220
rect 8996 12180 9002 12192
rect 9309 12189 9321 12192
rect 9355 12189 9367 12223
rect 9309 12183 9367 12189
rect 9585 12223 9643 12229
rect 9585 12189 9597 12223
rect 9631 12220 9643 12223
rect 9858 12220 9864 12232
rect 9631 12192 9864 12220
rect 9631 12189 9643 12192
rect 9585 12183 9643 12189
rect 9858 12180 9864 12192
rect 9916 12180 9922 12232
rect 12636 12229 12664 12260
rect 12621 12223 12679 12229
rect 12621 12189 12633 12223
rect 12667 12189 12679 12223
rect 12621 12183 12679 12189
rect 12805 12223 12863 12229
rect 12805 12189 12817 12223
rect 12851 12189 12863 12223
rect 14476 12220 14504 12387
rect 17126 12384 17132 12396
rect 17184 12384 17190 12436
rect 21174 12384 21180 12436
rect 21232 12424 21238 12436
rect 22646 12424 22652 12436
rect 21232 12396 22652 12424
rect 21232 12384 21238 12396
rect 22646 12384 22652 12396
rect 22704 12384 22710 12436
rect 30190 12424 30196 12436
rect 28552 12396 30196 12424
rect 19334 12356 19340 12368
rect 14936 12328 19340 12356
rect 14936 12220 14964 12328
rect 19334 12316 19340 12328
rect 19392 12356 19398 12368
rect 21082 12356 21088 12368
rect 19392 12328 21088 12356
rect 19392 12316 19398 12328
rect 21082 12316 21088 12328
rect 21140 12316 21146 12368
rect 21192 12328 21680 12356
rect 21192 12288 21220 12328
rect 15672 12260 21220 12288
rect 21652 12288 21680 12328
rect 22189 12291 22247 12297
rect 22189 12288 22201 12291
rect 21652 12260 22201 12288
rect 15013 12223 15071 12229
rect 15013 12220 15025 12223
rect 14476 12192 15025 12220
rect 12805 12183 12863 12189
rect 15013 12189 15025 12192
rect 15059 12189 15071 12223
rect 15013 12183 15071 12189
rect 9674 12152 9680 12164
rect 7760 12124 9680 12152
rect 9674 12112 9680 12124
rect 9732 12112 9738 12164
rect 12820 12152 12848 12183
rect 15102 12180 15108 12232
rect 15160 12220 15166 12232
rect 15197 12223 15255 12229
rect 15197 12220 15209 12223
rect 15160 12192 15209 12220
rect 15160 12180 15166 12192
rect 15197 12189 15209 12192
rect 15243 12220 15255 12223
rect 15562 12220 15568 12232
rect 15243 12192 15568 12220
rect 15243 12189 15255 12192
rect 15197 12183 15255 12189
rect 15562 12180 15568 12192
rect 15620 12180 15626 12232
rect 15672 12152 15700 12260
rect 22189 12257 22201 12260
rect 22235 12257 22247 12291
rect 22189 12251 22247 12257
rect 16669 12223 16727 12229
rect 16669 12220 16681 12223
rect 16592 12192 16681 12220
rect 12820 12124 15700 12152
rect 15746 12112 15752 12164
rect 15804 12152 15810 12164
rect 15841 12155 15899 12161
rect 15841 12152 15853 12155
rect 15804 12124 15853 12152
rect 15804 12112 15810 12124
rect 15841 12121 15853 12124
rect 15887 12152 15899 12155
rect 16206 12152 16212 12164
rect 15887 12124 16212 12152
rect 15887 12121 15899 12124
rect 15841 12115 15899 12121
rect 16206 12112 16212 12124
rect 16264 12112 16270 12164
rect 5307 12056 6316 12084
rect 9493 12087 9551 12093
rect 5307 12053 5319 12056
rect 5261 12047 5319 12053
rect 9493 12053 9505 12087
rect 9539 12084 9551 12087
rect 10137 12087 10195 12093
rect 10137 12084 10149 12087
rect 9539 12056 10149 12084
rect 9539 12053 9551 12056
rect 9493 12047 9551 12053
rect 10137 12053 10149 12056
rect 10183 12084 10195 12087
rect 10226 12084 10232 12096
rect 10183 12056 10232 12084
rect 10183 12053 10195 12056
rect 10137 12047 10195 12053
rect 10226 12044 10232 12056
rect 10284 12044 10290 12096
rect 11793 12087 11851 12093
rect 11793 12053 11805 12087
rect 11839 12084 11851 12087
rect 11882 12084 11888 12096
rect 11839 12056 11888 12084
rect 11839 12053 11851 12056
rect 11793 12047 11851 12053
rect 11882 12044 11888 12056
rect 11940 12044 11946 12096
rect 15105 12087 15163 12093
rect 15105 12053 15117 12087
rect 15151 12084 15163 12087
rect 15654 12084 15660 12096
rect 15151 12056 15660 12084
rect 15151 12053 15163 12056
rect 15105 12047 15163 12053
rect 15654 12044 15660 12056
rect 15712 12044 15718 12096
rect 16482 12084 16488 12096
rect 16443 12056 16488 12084
rect 16482 12044 16488 12056
rect 16540 12044 16546 12096
rect 16592 12084 16620 12192
rect 16669 12189 16681 12192
rect 16715 12189 16727 12223
rect 17034 12220 17040 12232
rect 16995 12192 17040 12220
rect 16669 12183 16727 12189
rect 17034 12180 17040 12192
rect 17092 12180 17098 12232
rect 19426 12220 19432 12232
rect 19387 12192 19432 12220
rect 19426 12180 19432 12192
rect 19484 12180 19490 12232
rect 20073 12223 20131 12229
rect 20073 12189 20085 12223
rect 20119 12189 20131 12223
rect 20073 12183 20131 12189
rect 16758 12152 16764 12164
rect 16719 12124 16764 12152
rect 16758 12112 16764 12124
rect 16816 12112 16822 12164
rect 16853 12155 16911 12161
rect 16853 12121 16865 12155
rect 16899 12152 16911 12155
rect 17126 12152 17132 12164
rect 16899 12124 17132 12152
rect 16899 12121 16911 12124
rect 16853 12115 16911 12121
rect 17126 12112 17132 12124
rect 17184 12152 17190 12164
rect 17770 12152 17776 12164
rect 17184 12124 17776 12152
rect 17184 12112 17190 12124
rect 17770 12112 17776 12124
rect 17828 12112 17834 12164
rect 18782 12112 18788 12164
rect 18840 12152 18846 12164
rect 19613 12155 19671 12161
rect 19613 12152 19625 12155
rect 18840 12124 19625 12152
rect 18840 12112 18846 12124
rect 19613 12121 19625 12124
rect 19659 12121 19671 12155
rect 19613 12115 19671 12121
rect 17586 12084 17592 12096
rect 16592 12056 17592 12084
rect 17586 12044 17592 12056
rect 17644 12044 17650 12096
rect 18506 12084 18512 12096
rect 18467 12056 18512 12084
rect 18506 12044 18512 12056
rect 18564 12044 18570 12096
rect 19242 12084 19248 12096
rect 19203 12056 19248 12084
rect 19242 12044 19248 12056
rect 19300 12044 19306 12096
rect 20088 12084 20116 12183
rect 20162 12180 20168 12232
rect 20220 12220 20226 12232
rect 20346 12220 20352 12232
rect 20220 12192 20265 12220
rect 20307 12192 20352 12220
rect 20220 12180 20226 12192
rect 20346 12180 20352 12192
rect 20404 12180 20410 12232
rect 20441 12223 20499 12229
rect 20441 12189 20453 12223
rect 20487 12220 20499 12223
rect 21174 12220 21180 12232
rect 20487 12192 21180 12220
rect 20487 12189 20499 12192
rect 20441 12183 20499 12189
rect 21174 12180 21180 12192
rect 21232 12180 21238 12232
rect 21361 12223 21419 12229
rect 21361 12189 21373 12223
rect 21407 12189 21419 12223
rect 21361 12183 21419 12189
rect 21545 12223 21603 12229
rect 21545 12189 21557 12223
rect 21591 12220 21603 12223
rect 21729 12223 21787 12229
rect 21591 12192 21680 12220
rect 21591 12189 21603 12192
rect 21545 12183 21603 12189
rect 20622 12152 20628 12164
rect 20583 12124 20628 12152
rect 20622 12112 20628 12124
rect 20680 12112 20686 12164
rect 20990 12112 20996 12164
rect 21048 12152 21054 12164
rect 21376 12152 21404 12183
rect 21048 12124 21404 12152
rect 21048 12112 21054 12124
rect 21450 12112 21456 12164
rect 21508 12152 21514 12164
rect 21652 12152 21680 12192
rect 21729 12189 21741 12223
rect 21775 12220 21787 12223
rect 22094 12220 22100 12232
rect 21775 12192 22100 12220
rect 21775 12189 21787 12192
rect 21729 12183 21787 12189
rect 22094 12180 22100 12192
rect 22152 12180 22158 12232
rect 22370 12220 22376 12232
rect 22331 12192 22376 12220
rect 22370 12180 22376 12192
rect 22428 12180 22434 12232
rect 22462 12180 22468 12232
rect 22520 12220 22526 12232
rect 22557 12223 22615 12229
rect 22557 12220 22569 12223
rect 22520 12192 22569 12220
rect 22520 12180 22526 12192
rect 22557 12189 22569 12192
rect 22603 12189 22615 12223
rect 22557 12183 22615 12189
rect 22649 12223 22707 12229
rect 22649 12189 22661 12223
rect 22695 12220 22707 12223
rect 23109 12223 23167 12229
rect 23109 12220 23121 12223
rect 22695 12192 23121 12220
rect 22695 12189 22707 12192
rect 22649 12183 22707 12189
rect 23109 12189 23121 12192
rect 23155 12220 23167 12223
rect 24210 12220 24216 12232
rect 23155 12192 24216 12220
rect 23155 12189 23167 12192
rect 23109 12183 23167 12189
rect 24210 12180 24216 12192
rect 24268 12180 24274 12232
rect 24670 12180 24676 12232
rect 24728 12220 24734 12232
rect 25041 12223 25099 12229
rect 25041 12220 25053 12223
rect 24728 12192 25053 12220
rect 24728 12180 24734 12192
rect 25041 12189 25053 12192
rect 25087 12189 25099 12223
rect 25041 12183 25099 12189
rect 25682 12180 25688 12232
rect 25740 12220 25746 12232
rect 28552 12220 28580 12396
rect 30190 12384 30196 12396
rect 30248 12384 30254 12436
rect 30282 12384 30288 12436
rect 30340 12424 30346 12436
rect 32490 12424 32496 12436
rect 30340 12396 31754 12424
rect 32451 12396 32496 12424
rect 30340 12384 30346 12396
rect 28810 12316 28816 12368
rect 28868 12356 28874 12368
rect 28997 12359 29055 12365
rect 28868 12328 28948 12356
rect 28868 12316 28874 12328
rect 28626 12248 28632 12300
rect 28684 12288 28690 12300
rect 28920 12288 28948 12328
rect 28997 12325 29009 12359
rect 29043 12356 29055 12359
rect 30650 12356 30656 12368
rect 29043 12328 30656 12356
rect 29043 12325 29055 12328
rect 28997 12319 29055 12325
rect 30650 12316 30656 12328
rect 30708 12316 30714 12368
rect 30837 12359 30895 12365
rect 30837 12325 30849 12359
rect 30883 12325 30895 12359
rect 31726 12356 31754 12396
rect 32490 12384 32496 12396
rect 32548 12384 32554 12436
rect 34790 12384 34796 12436
rect 34848 12424 34854 12436
rect 34885 12427 34943 12433
rect 34885 12424 34897 12427
rect 34848 12396 34897 12424
rect 34848 12384 34854 12396
rect 34885 12393 34897 12396
rect 34931 12393 34943 12427
rect 37550 12424 37556 12436
rect 37511 12396 37556 12424
rect 34885 12387 34943 12393
rect 37550 12384 37556 12396
rect 37608 12384 37614 12436
rect 40405 12359 40463 12365
rect 40405 12356 40417 12359
rect 31726 12328 40417 12356
rect 30837 12319 30895 12325
rect 40405 12325 40417 12328
rect 40451 12356 40463 12359
rect 46017 12359 46075 12365
rect 40451 12328 41092 12356
rect 40451 12325 40463 12328
rect 40405 12319 40463 12325
rect 28684 12260 28856 12288
rect 28920 12260 29868 12288
rect 28684 12248 28690 12260
rect 28828 12229 28856 12260
rect 28721 12223 28779 12229
rect 28721 12220 28733 12223
rect 25740 12192 28733 12220
rect 25740 12180 25746 12192
rect 28721 12189 28733 12192
rect 28767 12189 28779 12223
rect 28721 12183 28779 12189
rect 28813 12223 28871 12229
rect 28813 12189 28825 12223
rect 28859 12189 28871 12223
rect 28813 12183 28871 12189
rect 28920 12192 29132 12220
rect 21910 12152 21916 12164
rect 21508 12124 21553 12152
rect 21652 12124 21916 12152
rect 21508 12112 21514 12124
rect 21910 12112 21916 12124
rect 21968 12112 21974 12164
rect 28920 12152 28948 12192
rect 22066 12124 28948 12152
rect 28997 12155 29055 12161
rect 21177 12087 21235 12093
rect 21177 12084 21189 12087
rect 20088 12056 21189 12084
rect 21177 12053 21189 12056
rect 21223 12053 21235 12087
rect 21177 12047 21235 12053
rect 21266 12044 21272 12096
rect 21324 12084 21330 12096
rect 22066 12084 22094 12124
rect 28997 12121 29009 12155
rect 29043 12121 29055 12155
rect 29104 12152 29132 12192
rect 29638 12180 29644 12232
rect 29696 12220 29702 12232
rect 29840 12229 29868 12260
rect 30006 12248 30012 12300
rect 30064 12288 30070 12300
rect 30852 12288 30880 12319
rect 34514 12288 34520 12300
rect 30064 12260 30604 12288
rect 30852 12260 34520 12288
rect 30064 12248 30070 12260
rect 29733 12223 29791 12229
rect 29733 12220 29745 12223
rect 29696 12192 29745 12220
rect 29696 12180 29702 12192
rect 29733 12189 29745 12192
rect 29779 12189 29791 12223
rect 29733 12183 29791 12189
rect 29825 12223 29883 12229
rect 29825 12189 29837 12223
rect 29871 12189 29883 12223
rect 30098 12220 30104 12232
rect 30059 12192 30104 12220
rect 29825 12183 29883 12189
rect 30098 12180 30104 12192
rect 30156 12180 30162 12232
rect 30576 12229 30604 12260
rect 34514 12248 34520 12260
rect 34572 12288 34578 12300
rect 38746 12288 38752 12300
rect 34572 12260 34928 12288
rect 34572 12248 34578 12260
rect 30561 12223 30619 12229
rect 30561 12189 30573 12223
rect 30607 12189 30619 12223
rect 30834 12220 30840 12232
rect 30795 12192 30840 12220
rect 30561 12183 30619 12189
rect 30834 12180 30840 12192
rect 30892 12180 30898 12232
rect 31754 12220 31760 12232
rect 31726 12180 31760 12220
rect 31812 12220 31818 12232
rect 32493 12223 32551 12229
rect 32493 12220 32505 12223
rect 31812 12192 32505 12220
rect 31812 12180 31818 12192
rect 32493 12189 32505 12192
rect 32539 12189 32551 12223
rect 32493 12183 32551 12189
rect 32585 12223 32643 12229
rect 32585 12189 32597 12223
rect 32631 12189 32643 12223
rect 32585 12183 32643 12189
rect 29914 12152 29920 12164
rect 29104 12124 29684 12152
rect 29875 12124 29920 12152
rect 28997 12115 29055 12121
rect 21324 12056 22094 12084
rect 25133 12087 25191 12093
rect 21324 12044 21330 12056
rect 25133 12053 25145 12087
rect 25179 12084 25191 12087
rect 25774 12084 25780 12096
rect 25179 12056 25780 12084
rect 25179 12053 25191 12056
rect 25133 12047 25191 12053
rect 25774 12044 25780 12056
rect 25832 12044 25838 12096
rect 29012 12084 29040 12115
rect 29549 12087 29607 12093
rect 29549 12084 29561 12087
rect 29012 12056 29561 12084
rect 29549 12053 29561 12056
rect 29595 12053 29607 12087
rect 29656 12084 29684 12124
rect 29914 12112 29920 12124
rect 29972 12112 29978 12164
rect 31389 12155 31447 12161
rect 31389 12152 31401 12155
rect 30024 12124 31401 12152
rect 30024 12084 30052 12124
rect 31389 12121 31401 12124
rect 31435 12152 31447 12155
rect 31726 12152 31754 12180
rect 32600 12152 32628 12183
rect 34698 12152 34704 12164
rect 31435 12124 31754 12152
rect 31956 12124 32628 12152
rect 34659 12124 34704 12152
rect 31435 12121 31447 12124
rect 31389 12115 31447 12121
rect 31956 12096 31984 12124
rect 34698 12112 34704 12124
rect 34756 12112 34762 12164
rect 34900 12161 34928 12260
rect 38212 12260 38752 12288
rect 38212 12229 38240 12260
rect 38746 12248 38752 12260
rect 38804 12248 38810 12300
rect 41064 12297 41092 12328
rect 46017 12325 46029 12359
rect 46063 12325 46075 12359
rect 46017 12319 46075 12325
rect 51445 12359 51503 12365
rect 51445 12325 51457 12359
rect 51491 12356 51503 12359
rect 51491 12328 52316 12356
rect 51491 12325 51503 12328
rect 51445 12319 51503 12325
rect 41049 12291 41107 12297
rect 41049 12257 41061 12291
rect 41095 12257 41107 12291
rect 46032 12288 46060 12319
rect 49237 12291 49295 12297
rect 46032 12260 48820 12288
rect 41049 12251 41107 12257
rect 38197 12223 38255 12229
rect 38197 12189 38209 12223
rect 38243 12189 38255 12223
rect 38197 12183 38255 12189
rect 38286 12180 38292 12232
rect 38344 12220 38350 12232
rect 38473 12223 38531 12229
rect 38344 12192 38389 12220
rect 38344 12180 38350 12192
rect 38473 12189 38485 12223
rect 38519 12189 38531 12223
rect 38473 12183 38531 12189
rect 34900 12155 34959 12161
rect 34900 12124 34913 12155
rect 34901 12121 34913 12124
rect 34947 12121 34959 12155
rect 34901 12115 34959 12121
rect 37182 12112 37188 12164
rect 37240 12152 37246 12164
rect 38378 12152 38384 12164
rect 37240 12124 38384 12152
rect 37240 12112 37246 12124
rect 38378 12112 38384 12124
rect 38436 12152 38442 12164
rect 38488 12152 38516 12183
rect 40678 12180 40684 12232
rect 40736 12220 40742 12232
rect 41138 12220 41144 12232
rect 40736 12192 41144 12220
rect 40736 12180 40742 12192
rect 41138 12180 41144 12192
rect 41196 12180 41202 12232
rect 45738 12220 45744 12232
rect 45699 12192 45744 12220
rect 45738 12180 45744 12192
rect 45796 12180 45802 12232
rect 48590 12220 48596 12232
rect 48551 12192 48596 12220
rect 48590 12180 48596 12192
rect 48648 12180 48654 12232
rect 48792 12229 48820 12260
rect 49237 12257 49249 12291
rect 49283 12288 49295 12291
rect 51353 12291 51411 12297
rect 51353 12288 51365 12291
rect 49283 12260 51365 12288
rect 49283 12257 49295 12260
rect 49237 12251 49295 12257
rect 51353 12257 51365 12260
rect 51399 12288 51411 12291
rect 51718 12288 51724 12300
rect 51399 12260 51724 12288
rect 51399 12257 51411 12260
rect 51353 12251 51411 12257
rect 51718 12248 51724 12260
rect 51776 12248 51782 12300
rect 48777 12223 48835 12229
rect 48777 12189 48789 12223
rect 48823 12189 48835 12223
rect 49050 12220 49056 12232
rect 49011 12192 49056 12220
rect 48777 12183 48835 12189
rect 38436 12124 38516 12152
rect 38657 12155 38715 12161
rect 38436 12112 38442 12124
rect 38657 12121 38669 12155
rect 38703 12152 38715 12155
rect 43806 12152 43812 12164
rect 38703 12124 43812 12152
rect 38703 12121 38715 12124
rect 38657 12115 38715 12121
rect 43806 12112 43812 12124
rect 43864 12112 43870 12164
rect 45370 12112 45376 12164
rect 45428 12152 45434 12164
rect 46017 12155 46075 12161
rect 46017 12152 46029 12155
rect 45428 12124 46029 12152
rect 45428 12112 45434 12124
rect 46017 12121 46029 12124
rect 46063 12121 46075 12155
rect 48792 12152 48820 12183
rect 49050 12180 49056 12192
rect 49108 12180 49114 12232
rect 51442 12180 51448 12232
rect 51500 12220 51506 12232
rect 51500 12192 51545 12220
rect 51500 12180 51506 12192
rect 51626 12180 51632 12232
rect 51684 12220 51690 12232
rect 52288 12229 52316 12328
rect 56520 12260 57284 12288
rect 56520 12232 56548 12260
rect 52089 12223 52147 12229
rect 52089 12220 52101 12223
rect 51684 12192 52101 12220
rect 51684 12180 51690 12192
rect 52089 12189 52101 12192
rect 52135 12189 52147 12223
rect 52089 12183 52147 12189
rect 52273 12223 52331 12229
rect 52273 12189 52285 12223
rect 52319 12220 52331 12223
rect 52454 12220 52460 12232
rect 52319 12192 52460 12220
rect 52319 12189 52331 12192
rect 52273 12183 52331 12189
rect 52454 12180 52460 12192
rect 52512 12180 52518 12232
rect 56413 12223 56471 12229
rect 56413 12189 56425 12223
rect 56459 12220 56471 12223
rect 56502 12220 56508 12232
rect 56459 12192 56508 12220
rect 56459 12189 56471 12192
rect 56413 12183 56471 12189
rect 56502 12180 56508 12192
rect 56560 12180 56566 12232
rect 57057 12223 57115 12229
rect 57057 12189 57069 12223
rect 57103 12220 57115 12223
rect 57146 12220 57152 12232
rect 57103 12192 57152 12220
rect 57103 12189 57115 12192
rect 57057 12183 57115 12189
rect 57146 12180 57152 12192
rect 57204 12180 57210 12232
rect 57256 12229 57284 12260
rect 57790 12248 57796 12300
rect 57848 12288 57854 12300
rect 57885 12291 57943 12297
rect 57885 12288 57897 12291
rect 57848 12260 57897 12288
rect 57848 12248 57854 12260
rect 57885 12257 57897 12260
rect 57931 12257 57943 12291
rect 57885 12251 57943 12257
rect 57241 12223 57299 12229
rect 57241 12189 57253 12223
rect 57287 12189 57299 12223
rect 58158 12220 58164 12232
rect 58119 12192 58164 12220
rect 57241 12183 57299 12189
rect 58158 12180 58164 12192
rect 58216 12180 58222 12232
rect 48958 12152 48964 12164
rect 48792 12124 48964 12152
rect 46017 12115 46075 12121
rect 48958 12112 48964 12124
rect 49016 12112 49022 12164
rect 51166 12152 51172 12164
rect 51127 12124 51172 12152
rect 51166 12112 51172 12124
rect 51224 12152 51230 12164
rect 51644 12152 51672 12180
rect 51902 12152 51908 12164
rect 51224 12124 51672 12152
rect 51863 12124 51908 12152
rect 51224 12112 51230 12124
rect 51902 12112 51908 12124
rect 51960 12112 51966 12164
rect 56226 12152 56232 12164
rect 56187 12124 56232 12152
rect 56226 12112 56232 12124
rect 56284 12112 56290 12164
rect 29656 12056 30052 12084
rect 30653 12087 30711 12093
rect 29549 12047 29607 12053
rect 30653 12053 30665 12087
rect 30699 12084 30711 12087
rect 30742 12084 30748 12096
rect 30699 12056 30748 12084
rect 30699 12053 30711 12056
rect 30653 12047 30711 12053
rect 30742 12044 30748 12056
rect 30800 12044 30806 12096
rect 31938 12084 31944 12096
rect 31899 12056 31944 12084
rect 31938 12044 31944 12056
rect 31996 12044 32002 12096
rect 32861 12087 32919 12093
rect 32861 12053 32873 12087
rect 32907 12084 32919 12087
rect 33778 12084 33784 12096
rect 32907 12056 33784 12084
rect 32907 12053 32919 12056
rect 32861 12047 32919 12053
rect 33778 12044 33784 12056
rect 33836 12044 33842 12096
rect 35069 12087 35127 12093
rect 35069 12053 35081 12087
rect 35115 12084 35127 12087
rect 35342 12084 35348 12096
rect 35115 12056 35348 12084
rect 35115 12053 35127 12056
rect 35069 12047 35127 12053
rect 35342 12044 35348 12056
rect 35400 12044 35406 12096
rect 41509 12087 41567 12093
rect 41509 12053 41521 12087
rect 41555 12084 41567 12087
rect 43162 12084 43168 12096
rect 41555 12056 43168 12084
rect 41555 12053 41567 12056
rect 41509 12047 41567 12053
rect 43162 12044 43168 12056
rect 43220 12044 43226 12096
rect 43714 12044 43720 12096
rect 43772 12084 43778 12096
rect 45830 12084 45836 12096
rect 43772 12056 45836 12084
rect 43772 12044 43778 12056
rect 45830 12044 45836 12056
rect 45888 12044 45894 12096
rect 56594 12084 56600 12096
rect 56555 12056 56600 12084
rect 56594 12044 56600 12056
rect 56652 12044 56658 12096
rect 57054 12084 57060 12096
rect 57015 12056 57060 12084
rect 57054 12044 57060 12056
rect 57112 12044 57118 12096
rect 1104 11994 58880 12016
rect 1104 11942 19574 11994
rect 19626 11942 19638 11994
rect 19690 11942 19702 11994
rect 19754 11942 19766 11994
rect 19818 11942 19830 11994
rect 19882 11942 50294 11994
rect 50346 11942 50358 11994
rect 50410 11942 50422 11994
rect 50474 11942 50486 11994
rect 50538 11942 50550 11994
rect 50602 11942 58880 11994
rect 1104 11920 58880 11942
rect 4246 11840 4252 11892
rect 4304 11880 4310 11892
rect 5629 11883 5687 11889
rect 5629 11880 5641 11883
rect 4304 11852 5641 11880
rect 4304 11840 4310 11852
rect 5629 11849 5641 11852
rect 5675 11849 5687 11883
rect 5629 11843 5687 11849
rect 5718 11840 5724 11892
rect 5776 11880 5782 11892
rect 6457 11883 6515 11889
rect 6457 11880 6469 11883
rect 5776 11852 6469 11880
rect 5776 11840 5782 11852
rect 6457 11849 6469 11852
rect 6503 11849 6515 11883
rect 6457 11843 6515 11849
rect 7282 11840 7288 11892
rect 7340 11880 7346 11892
rect 8389 11883 8447 11889
rect 8389 11880 8401 11883
rect 7340 11852 8401 11880
rect 7340 11840 7346 11852
rect 8389 11849 8401 11852
rect 8435 11849 8447 11883
rect 8938 11880 8944 11892
rect 8899 11852 8944 11880
rect 8389 11843 8447 11849
rect 8938 11840 8944 11852
rect 8996 11840 9002 11892
rect 17310 11840 17316 11892
rect 17368 11880 17374 11892
rect 18782 11880 18788 11892
rect 17368 11852 18788 11880
rect 17368 11840 17374 11852
rect 18782 11840 18788 11852
rect 18840 11840 18846 11892
rect 19334 11880 19340 11892
rect 19295 11852 19340 11880
rect 19334 11840 19340 11852
rect 19392 11840 19398 11892
rect 19981 11883 20039 11889
rect 19981 11849 19993 11883
rect 20027 11880 20039 11883
rect 20162 11880 20168 11892
rect 20027 11852 20168 11880
rect 20027 11849 20039 11852
rect 19981 11843 20039 11849
rect 20162 11840 20168 11852
rect 20220 11840 20226 11892
rect 21266 11880 21272 11892
rect 21100 11852 21272 11880
rect 3602 11812 3608 11824
rect 3344 11784 3608 11812
rect 3053 11747 3111 11753
rect 3053 11713 3065 11747
rect 3099 11713 3111 11747
rect 3053 11707 3111 11713
rect 3145 11747 3203 11753
rect 3145 11713 3157 11747
rect 3191 11744 3203 11747
rect 3234 11744 3240 11756
rect 3191 11716 3240 11744
rect 3191 11713 3203 11716
rect 3145 11707 3203 11713
rect 3068 11676 3096 11707
rect 3234 11704 3240 11716
rect 3292 11704 3298 11756
rect 3344 11753 3372 11784
rect 3602 11772 3608 11784
rect 3660 11772 3666 11824
rect 5736 11812 5764 11840
rect 8956 11812 8984 11840
rect 12624 11824 12676 11830
rect 4080 11784 5764 11812
rect 8312 11784 8984 11812
rect 9125 11815 9183 11821
rect 3329 11747 3387 11753
rect 3329 11713 3341 11747
rect 3375 11713 3387 11747
rect 3329 11707 3387 11713
rect 3421 11747 3479 11753
rect 3421 11713 3433 11747
rect 3467 11744 3479 11747
rect 3786 11744 3792 11756
rect 3467 11716 3792 11744
rect 3467 11713 3479 11716
rect 3421 11707 3479 11713
rect 3786 11704 3792 11716
rect 3844 11704 3850 11756
rect 3878 11704 3884 11756
rect 3936 11744 3942 11756
rect 4080 11753 4108 11784
rect 4065 11747 4123 11753
rect 3936 11716 3981 11744
rect 3936 11704 3942 11716
rect 4065 11713 4077 11747
rect 4111 11713 4123 11747
rect 4065 11707 4123 11713
rect 5629 11747 5687 11753
rect 5629 11713 5641 11747
rect 5675 11713 5687 11747
rect 5629 11707 5687 11713
rect 5813 11747 5871 11753
rect 5813 11713 5825 11747
rect 5859 11744 5871 11747
rect 6178 11744 6184 11756
rect 5859 11716 6184 11744
rect 5859 11713 5871 11716
rect 5813 11707 5871 11713
rect 3973 11679 4031 11685
rect 3973 11676 3985 11679
rect 3068 11648 3985 11676
rect 3973 11645 3985 11648
rect 4019 11645 4031 11679
rect 5644 11676 5672 11707
rect 6178 11704 6184 11716
rect 6236 11744 6242 11756
rect 6362 11744 6368 11756
rect 6236 11716 6368 11744
rect 6236 11704 6242 11716
rect 6362 11704 6368 11716
rect 6420 11704 6426 11756
rect 6549 11747 6607 11753
rect 6549 11713 6561 11747
rect 6595 11744 6607 11747
rect 7098 11744 7104 11756
rect 6595 11716 7104 11744
rect 6595 11713 6607 11716
rect 6549 11707 6607 11713
rect 6564 11676 6592 11707
rect 7098 11704 7104 11716
rect 7156 11704 7162 11756
rect 8312 11753 8340 11784
rect 9125 11781 9137 11815
rect 9171 11812 9183 11815
rect 9674 11812 9680 11824
rect 9171 11784 9680 11812
rect 9171 11781 9183 11784
rect 9125 11775 9183 11781
rect 9674 11772 9680 11784
rect 9732 11812 9738 11824
rect 10042 11812 10048 11824
rect 9732 11784 10048 11812
rect 9732 11772 9738 11784
rect 10042 11772 10048 11784
rect 10100 11772 10106 11824
rect 16298 11812 16304 11824
rect 12624 11766 12676 11772
rect 15488 11784 16304 11812
rect 8297 11747 8355 11753
rect 8297 11713 8309 11747
rect 8343 11713 8355 11747
rect 8297 11707 8355 11713
rect 8481 11747 8539 11753
rect 8481 11713 8493 11747
rect 8527 11713 8539 11747
rect 9306 11744 9312 11756
rect 9267 11716 9312 11744
rect 8481 11707 8539 11713
rect 5644 11648 6592 11676
rect 7837 11679 7895 11685
rect 3973 11639 4031 11645
rect 7837 11645 7849 11679
rect 7883 11676 7895 11679
rect 8018 11676 8024 11688
rect 7883 11648 8024 11676
rect 7883 11645 7895 11648
rect 7837 11639 7895 11645
rect 8018 11636 8024 11648
rect 8076 11676 8082 11688
rect 8496 11676 8524 11707
rect 9306 11704 9312 11716
rect 9364 11704 9370 11756
rect 11882 11744 11888 11756
rect 11843 11716 11888 11744
rect 11882 11704 11888 11716
rect 11940 11704 11946 11756
rect 12342 11744 12348 11756
rect 12303 11716 12348 11744
rect 12342 11704 12348 11716
rect 12400 11704 12406 11756
rect 15378 11744 15384 11756
rect 15291 11716 15384 11744
rect 15378 11704 15384 11716
rect 15436 11704 15442 11756
rect 15488 11753 15516 11784
rect 16298 11772 16304 11784
rect 16356 11812 16362 11824
rect 18800 11812 18828 11840
rect 21100 11812 21128 11852
rect 21266 11840 21272 11852
rect 21324 11840 21330 11892
rect 21913 11883 21971 11889
rect 21913 11849 21925 11883
rect 21959 11880 21971 11883
rect 29638 11880 29644 11892
rect 21959 11852 22094 11880
rect 21959 11849 21971 11852
rect 21913 11843 21971 11849
rect 16356 11784 16620 11812
rect 18800 11784 21128 11812
rect 21177 11815 21235 11821
rect 16356 11772 16362 11784
rect 15473 11747 15531 11753
rect 15473 11713 15485 11747
rect 15519 11713 15531 11747
rect 15654 11744 15660 11756
rect 15615 11716 15660 11744
rect 15473 11707 15531 11713
rect 15654 11704 15660 11716
rect 15712 11704 15718 11756
rect 15749 11747 15807 11753
rect 15749 11713 15761 11747
rect 15795 11744 15807 11747
rect 16482 11744 16488 11756
rect 15795 11716 16488 11744
rect 15795 11713 15807 11716
rect 15749 11707 15807 11713
rect 16482 11704 16488 11716
rect 16540 11704 16546 11756
rect 10226 11676 10232 11688
rect 8076 11648 10232 11676
rect 8076 11636 8082 11648
rect 10226 11636 10232 11648
rect 10284 11636 10290 11688
rect 15396 11676 15424 11704
rect 16114 11676 16120 11688
rect 15396 11648 16120 11676
rect 16114 11636 16120 11648
rect 16172 11636 16178 11688
rect 16592 11676 16620 11784
rect 21177 11781 21189 11815
rect 21223 11812 21235 11815
rect 21450 11812 21456 11824
rect 21223 11784 21456 11812
rect 21223 11781 21235 11784
rect 21177 11775 21235 11781
rect 21450 11772 21456 11784
rect 21508 11772 21514 11824
rect 22066 11812 22094 11852
rect 25608 11852 29644 11880
rect 22741 11815 22799 11821
rect 22741 11812 22753 11815
rect 22066 11784 22753 11812
rect 22741 11781 22753 11784
rect 22787 11812 22799 11815
rect 23566 11812 23572 11824
rect 22787 11784 23572 11812
rect 22787 11781 22799 11784
rect 22741 11775 22799 11781
rect 23566 11772 23572 11784
rect 23624 11772 23630 11824
rect 16666 11704 16672 11756
rect 16724 11744 16730 11756
rect 16807 11747 16865 11753
rect 16807 11744 16819 11747
rect 16724 11716 16819 11744
rect 16724 11704 16730 11716
rect 16807 11713 16819 11716
rect 16853 11713 16865 11747
rect 16942 11744 16948 11756
rect 16903 11716 16948 11744
rect 16807 11707 16865 11713
rect 16942 11704 16948 11716
rect 17000 11704 17006 11756
rect 17037 11747 17095 11753
rect 17037 11713 17049 11747
rect 17083 11744 17095 11747
rect 17126 11744 17132 11756
rect 17083 11716 17132 11744
rect 17083 11713 17095 11716
rect 17037 11707 17095 11713
rect 17126 11704 17132 11716
rect 17184 11704 17190 11756
rect 17221 11747 17279 11753
rect 17221 11713 17233 11747
rect 17267 11713 17279 11747
rect 17221 11707 17279 11713
rect 17236 11676 17264 11707
rect 19334 11704 19340 11756
rect 19392 11744 19398 11756
rect 19889 11747 19947 11753
rect 19889 11744 19901 11747
rect 19392 11716 19901 11744
rect 19392 11704 19398 11716
rect 19889 11713 19901 11716
rect 19935 11713 19947 11747
rect 19889 11707 19947 11713
rect 20073 11747 20131 11753
rect 20073 11713 20085 11747
rect 20119 11744 20131 11747
rect 20438 11744 20444 11756
rect 20119 11716 20444 11744
rect 20119 11713 20131 11716
rect 20073 11707 20131 11713
rect 20438 11704 20444 11716
rect 20496 11704 20502 11756
rect 22278 11704 22284 11756
rect 22336 11744 22342 11756
rect 22373 11747 22431 11753
rect 22373 11744 22385 11747
rect 22336 11716 22385 11744
rect 22336 11704 22342 11716
rect 22373 11713 22385 11716
rect 22419 11713 22431 11747
rect 22373 11707 22431 11713
rect 22466 11747 22524 11753
rect 22466 11713 22478 11747
rect 22512 11713 22524 11747
rect 22646 11744 22652 11756
rect 22607 11716 22652 11744
rect 22466 11707 22524 11713
rect 22094 11676 22100 11688
rect 16592 11648 22100 11676
rect 22094 11636 22100 11648
rect 22152 11676 22158 11688
rect 22481 11676 22509 11707
rect 22646 11704 22652 11716
rect 22704 11704 22710 11756
rect 22830 11704 22836 11756
rect 22888 11753 22894 11756
rect 22888 11744 22896 11753
rect 22888 11716 22981 11744
rect 22888 11707 22896 11716
rect 22888 11704 22894 11707
rect 23658 11704 23664 11756
rect 23716 11744 23722 11756
rect 23753 11747 23811 11753
rect 23753 11744 23765 11747
rect 23716 11716 23765 11744
rect 23716 11704 23722 11716
rect 23753 11713 23765 11716
rect 23799 11744 23811 11747
rect 24486 11744 24492 11756
rect 23799 11716 24492 11744
rect 23799 11713 23811 11716
rect 23753 11707 23811 11713
rect 24486 11704 24492 11716
rect 24544 11704 24550 11756
rect 24946 11704 24952 11756
rect 25004 11744 25010 11756
rect 25608 11753 25636 11852
rect 25774 11812 25780 11824
rect 25735 11784 25780 11812
rect 25774 11772 25780 11784
rect 25832 11772 25838 11824
rect 27798 11772 27804 11824
rect 27856 11812 27862 11824
rect 28258 11812 28264 11824
rect 27856 11784 28264 11812
rect 27856 11772 27862 11784
rect 28258 11772 28264 11784
rect 28316 11812 28322 11824
rect 28445 11815 28503 11821
rect 28445 11812 28457 11815
rect 28316 11784 28457 11812
rect 28316 11772 28322 11784
rect 28445 11781 28457 11784
rect 28491 11781 28503 11815
rect 28445 11775 28503 11781
rect 25593 11747 25651 11753
rect 25593 11744 25605 11747
rect 25004 11716 25605 11744
rect 25004 11704 25010 11716
rect 25593 11713 25605 11716
rect 25639 11713 25651 11747
rect 25593 11707 25651 11713
rect 25685 11747 25743 11753
rect 25685 11713 25697 11747
rect 25731 11713 25743 11747
rect 25685 11707 25743 11713
rect 22152 11648 22509 11676
rect 22853 11676 22881 11704
rect 23934 11676 23940 11688
rect 22853 11648 23940 11676
rect 22152 11636 22158 11648
rect 23934 11636 23940 11648
rect 23992 11636 23998 11688
rect 25222 11636 25228 11688
rect 25280 11676 25286 11688
rect 25700 11676 25728 11707
rect 25280 11648 25728 11676
rect 25792 11676 25820 11772
rect 25958 11744 25964 11756
rect 25919 11716 25964 11744
rect 25958 11704 25964 11716
rect 26016 11704 26022 11756
rect 27614 11704 27620 11756
rect 27672 11744 27678 11756
rect 28166 11744 28172 11756
rect 27672 11716 28172 11744
rect 27672 11704 27678 11716
rect 28166 11704 28172 11716
rect 28224 11704 28230 11756
rect 28552 11753 28580 11852
rect 29638 11840 29644 11852
rect 29696 11840 29702 11892
rect 29733 11883 29791 11889
rect 29733 11849 29745 11883
rect 29779 11880 29791 11883
rect 29779 11852 30052 11880
rect 29779 11849 29791 11852
rect 29733 11843 29791 11849
rect 30024 11812 30052 11852
rect 30098 11840 30104 11892
rect 30156 11880 30162 11892
rect 30285 11883 30343 11889
rect 30285 11880 30297 11883
rect 30156 11852 30297 11880
rect 30156 11840 30162 11852
rect 30285 11849 30297 11852
rect 30331 11849 30343 11883
rect 30285 11843 30343 11849
rect 32217 11883 32275 11889
rect 32217 11849 32229 11883
rect 32263 11880 32275 11883
rect 32490 11880 32496 11892
rect 32263 11852 32496 11880
rect 32263 11849 32275 11852
rect 32217 11843 32275 11849
rect 32490 11840 32496 11852
rect 32548 11840 32554 11892
rect 33686 11880 33692 11892
rect 33060 11852 33692 11880
rect 30469 11815 30527 11821
rect 30469 11812 30481 11815
rect 29380 11784 29776 11812
rect 30024 11784 30481 11812
rect 28353 11747 28411 11753
rect 28353 11713 28365 11747
rect 28399 11713 28411 11747
rect 28353 11707 28411 11713
rect 28537 11747 28595 11753
rect 28537 11713 28549 11747
rect 28583 11713 28595 11747
rect 29178 11744 29184 11756
rect 29139 11716 29184 11744
rect 28537 11707 28595 11713
rect 27982 11676 27988 11688
rect 25792 11648 27988 11676
rect 25280 11636 25286 11648
rect 6454 11568 6460 11620
rect 6512 11608 6518 11620
rect 7098 11608 7104 11620
rect 6512 11580 7104 11608
rect 6512 11568 6518 11580
rect 7098 11568 7104 11580
rect 7156 11568 7162 11620
rect 14826 11568 14832 11620
rect 14884 11608 14890 11620
rect 15102 11608 15108 11620
rect 14884 11580 15108 11608
rect 14884 11568 14890 11580
rect 15102 11568 15108 11580
rect 15160 11608 15166 11620
rect 18506 11608 18512 11620
rect 15160 11580 18512 11608
rect 15160 11568 15166 11580
rect 18506 11568 18512 11580
rect 18564 11608 18570 11620
rect 18564 11580 23244 11608
rect 18564 11568 18570 11580
rect 2869 11543 2927 11549
rect 2869 11509 2881 11543
rect 2915 11540 2927 11543
rect 3694 11540 3700 11552
rect 2915 11512 3700 11540
rect 2915 11509 2927 11512
rect 2869 11503 2927 11509
rect 3694 11500 3700 11512
rect 3752 11500 3758 11552
rect 9858 11540 9864 11552
rect 9819 11512 9864 11540
rect 9858 11500 9864 11512
rect 9916 11500 9922 11552
rect 13170 11500 13176 11552
rect 13228 11540 13234 11552
rect 15197 11543 15255 11549
rect 15197 11540 15209 11543
rect 13228 11512 15209 11540
rect 13228 11500 13234 11512
rect 15197 11509 15209 11512
rect 15243 11509 15255 11543
rect 15197 11503 15255 11509
rect 15838 11500 15844 11552
rect 15896 11540 15902 11552
rect 16669 11543 16727 11549
rect 16669 11540 16681 11543
rect 15896 11512 16681 11540
rect 15896 11500 15902 11512
rect 16669 11509 16681 11512
rect 16715 11509 16727 11543
rect 21082 11540 21088 11552
rect 21043 11512 21088 11540
rect 16669 11503 16727 11509
rect 21082 11500 21088 11512
rect 21140 11500 21146 11552
rect 23014 11540 23020 11552
rect 22975 11512 23020 11540
rect 23014 11500 23020 11512
rect 23072 11500 23078 11552
rect 23216 11540 23244 11580
rect 23290 11568 23296 11620
rect 23348 11608 23354 11620
rect 23569 11611 23627 11617
rect 23569 11608 23581 11611
rect 23348 11580 23581 11608
rect 23348 11568 23354 11580
rect 23569 11577 23581 11580
rect 23615 11577 23627 11611
rect 25590 11608 25596 11620
rect 23569 11571 23627 11577
rect 25240 11580 25596 11608
rect 25240 11540 25268 11580
rect 25590 11568 25596 11580
rect 25648 11568 25654 11620
rect 23216 11512 25268 11540
rect 25314 11500 25320 11552
rect 25372 11540 25378 11552
rect 25409 11543 25467 11549
rect 25409 11540 25421 11543
rect 25372 11512 25421 11540
rect 25372 11500 25378 11512
rect 25409 11509 25421 11512
rect 25455 11509 25467 11543
rect 25700 11540 25728 11648
rect 27982 11636 27988 11648
rect 28040 11676 28046 11688
rect 28368 11676 28396 11707
rect 29178 11704 29184 11716
rect 29236 11704 29242 11756
rect 29380 11753 29408 11784
rect 29365 11747 29423 11753
rect 29365 11713 29377 11747
rect 29411 11713 29423 11747
rect 29365 11707 29423 11713
rect 29457 11747 29515 11753
rect 29457 11713 29469 11747
rect 29503 11713 29515 11747
rect 29457 11707 29515 11713
rect 29549 11747 29607 11753
rect 29549 11713 29561 11747
rect 29595 11744 29607 11747
rect 29638 11744 29644 11756
rect 29595 11716 29644 11744
rect 29595 11713 29607 11716
rect 29549 11707 29607 11713
rect 29380 11676 29408 11707
rect 28040 11648 29408 11676
rect 29472 11676 29500 11707
rect 29638 11704 29644 11716
rect 29696 11704 29702 11756
rect 29748 11744 29776 11784
rect 30469 11781 30481 11784
rect 30515 11781 30527 11815
rect 30469 11775 30527 11781
rect 30650 11772 30656 11824
rect 30708 11812 30714 11824
rect 33060 11812 33088 11852
rect 33686 11840 33692 11852
rect 33744 11880 33750 11892
rect 33797 11883 33855 11889
rect 33797 11880 33809 11883
rect 33744 11852 33809 11880
rect 33744 11840 33750 11852
rect 33797 11849 33809 11852
rect 33843 11849 33855 11883
rect 33797 11843 33855 11849
rect 34609 11883 34667 11889
rect 34609 11849 34621 11883
rect 34655 11880 34667 11883
rect 34790 11880 34796 11892
rect 34655 11852 34796 11880
rect 34655 11849 34667 11852
rect 34609 11843 34667 11849
rect 34790 11840 34796 11852
rect 34848 11840 34854 11892
rect 38565 11883 38623 11889
rect 38565 11849 38577 11883
rect 38611 11880 38623 11883
rect 45370 11880 45376 11892
rect 38611 11852 41414 11880
rect 45331 11852 45376 11880
rect 38611 11849 38623 11852
rect 38565 11843 38623 11849
rect 33594 11812 33600 11824
rect 30708 11784 33088 11812
rect 33555 11784 33600 11812
rect 30708 11772 30714 11784
rect 33594 11772 33600 11784
rect 33652 11772 33658 11824
rect 36262 11772 36268 11824
rect 36320 11812 36326 11824
rect 37737 11815 37795 11821
rect 37737 11812 37749 11815
rect 36320 11784 37749 11812
rect 36320 11772 36326 11784
rect 37737 11781 37749 11784
rect 37783 11781 37795 11815
rect 37737 11775 37795 11781
rect 38286 11772 38292 11824
rect 38344 11812 38350 11824
rect 38473 11815 38531 11821
rect 38473 11812 38485 11815
rect 38344 11784 38485 11812
rect 38344 11772 38350 11784
rect 38473 11781 38485 11784
rect 38519 11781 38531 11815
rect 38473 11775 38531 11781
rect 38657 11815 38715 11821
rect 38657 11781 38669 11815
rect 38703 11812 38715 11815
rect 38746 11812 38752 11824
rect 38703 11784 38752 11812
rect 38703 11781 38715 11784
rect 38657 11775 38715 11781
rect 38746 11772 38752 11784
rect 38804 11772 38810 11824
rect 41386 11812 41414 11852
rect 45370 11840 45376 11852
rect 45428 11840 45434 11892
rect 49053 11883 49111 11889
rect 49053 11849 49065 11883
rect 49099 11880 49111 11883
rect 51166 11880 51172 11892
rect 49099 11852 51172 11880
rect 49099 11849 49111 11852
rect 49053 11843 49111 11849
rect 51166 11840 51172 11852
rect 51224 11840 51230 11892
rect 58158 11880 58164 11892
rect 58119 11852 58164 11880
rect 58158 11840 58164 11852
rect 58216 11840 58222 11892
rect 43070 11812 43076 11824
rect 41386 11784 43076 11812
rect 43070 11772 43076 11784
rect 43128 11812 43134 11824
rect 43714 11812 43720 11824
rect 43128 11784 43484 11812
rect 43675 11784 43720 11812
rect 43128 11772 43134 11784
rect 29914 11744 29920 11756
rect 29748 11716 29920 11744
rect 29914 11704 29920 11716
rect 29972 11704 29978 11756
rect 30190 11744 30196 11756
rect 30151 11716 30196 11744
rect 30190 11704 30196 11716
rect 30248 11704 30254 11756
rect 34514 11744 34520 11756
rect 34475 11716 34520 11744
rect 34514 11704 34520 11716
rect 34572 11704 34578 11756
rect 34698 11704 34704 11756
rect 34756 11744 34762 11756
rect 34793 11747 34851 11753
rect 34793 11744 34805 11747
rect 34756 11716 34805 11744
rect 34756 11704 34762 11716
rect 34793 11713 34805 11716
rect 34839 11744 34851 11747
rect 36078 11744 36084 11756
rect 34839 11716 36084 11744
rect 34839 11713 34851 11716
rect 34793 11707 34851 11713
rect 36078 11704 36084 11716
rect 36136 11704 36142 11756
rect 38378 11744 38384 11756
rect 38339 11716 38384 11744
rect 38378 11704 38384 11716
rect 38436 11704 38442 11756
rect 39114 11744 39120 11756
rect 39075 11716 39120 11744
rect 39114 11704 39120 11716
rect 39172 11704 39178 11756
rect 43162 11744 43168 11756
rect 43123 11716 43168 11744
rect 43162 11704 43168 11716
rect 43220 11704 43226 11756
rect 43456 11753 43484 11784
rect 43714 11772 43720 11784
rect 43772 11772 43778 11824
rect 53469 11815 53527 11821
rect 44928 11784 46244 11812
rect 43441 11747 43499 11753
rect 43441 11713 43453 11747
rect 43487 11713 43499 11747
rect 43806 11744 43812 11756
rect 43767 11716 43812 11744
rect 43441 11707 43499 11713
rect 43806 11704 43812 11716
rect 43864 11704 43870 11756
rect 44928 11688 44956 11784
rect 45005 11747 45063 11753
rect 45005 11713 45017 11747
rect 45051 11744 45063 11747
rect 45462 11744 45468 11756
rect 45051 11716 45468 11744
rect 45051 11713 45063 11716
rect 45005 11707 45063 11713
rect 45462 11704 45468 11716
rect 45520 11704 45526 11756
rect 46106 11744 46112 11756
rect 46067 11716 46112 11744
rect 46106 11704 46112 11716
rect 46164 11704 46170 11756
rect 46216 11753 46244 11784
rect 53469 11781 53481 11815
rect 53515 11812 53527 11815
rect 54662 11812 54668 11824
rect 53515 11784 54668 11812
rect 53515 11781 53527 11784
rect 53469 11775 53527 11781
rect 54662 11772 54668 11784
rect 54720 11772 54726 11824
rect 56226 11772 56232 11824
rect 56284 11812 56290 11824
rect 56284 11784 57100 11812
rect 56284 11772 56290 11784
rect 46201 11747 46259 11753
rect 46201 11713 46213 11747
rect 46247 11713 46259 11747
rect 46201 11707 46259 11713
rect 48685 11747 48743 11753
rect 48685 11713 48697 11747
rect 48731 11744 48743 11747
rect 49050 11744 49056 11756
rect 48731 11716 49056 11744
rect 48731 11713 48743 11716
rect 48685 11707 48743 11713
rect 49050 11704 49056 11716
rect 49108 11704 49114 11756
rect 53653 11747 53711 11753
rect 53653 11713 53665 11747
rect 53699 11744 53711 11747
rect 53834 11744 53840 11756
rect 53699 11716 53840 11744
rect 53699 11713 53711 11716
rect 53653 11707 53711 11713
rect 53834 11704 53840 11716
rect 53892 11704 53898 11756
rect 56042 11744 56048 11756
rect 56003 11716 56048 11744
rect 56042 11704 56048 11716
rect 56100 11704 56106 11756
rect 56686 11744 56692 11756
rect 56647 11716 56692 11744
rect 56686 11704 56692 11716
rect 56744 11704 56750 11756
rect 57072 11753 57100 11784
rect 57057 11747 57115 11753
rect 57057 11713 57069 11747
rect 57103 11713 57115 11747
rect 57057 11707 57115 11713
rect 57146 11704 57152 11756
rect 57204 11744 57210 11756
rect 57241 11747 57299 11753
rect 57241 11744 57253 11747
rect 57204 11716 57253 11744
rect 57204 11704 57210 11716
rect 57241 11713 57253 11716
rect 57287 11713 57299 11747
rect 57241 11707 57299 11713
rect 30558 11676 30564 11688
rect 29472 11648 30564 11676
rect 28040 11636 28046 11648
rect 30558 11636 30564 11648
rect 30616 11636 30622 11688
rect 44910 11676 44916 11688
rect 44871 11648 44916 11676
rect 44910 11636 44916 11648
rect 44968 11636 44974 11688
rect 45922 11676 45928 11688
rect 45883 11648 45928 11676
rect 45922 11636 45928 11648
rect 45980 11636 45986 11688
rect 46017 11679 46075 11685
rect 46017 11645 46029 11679
rect 46063 11645 46075 11679
rect 46017 11639 46075 11645
rect 37921 11611 37979 11617
rect 37921 11577 37933 11611
rect 37967 11608 37979 11611
rect 38470 11608 38476 11620
rect 37967 11580 38476 11608
rect 37967 11577 37979 11580
rect 37921 11571 37979 11577
rect 38470 11568 38476 11580
rect 38528 11568 38534 11620
rect 27614 11540 27620 11552
rect 25700 11512 27620 11540
rect 25409 11503 25467 11509
rect 27614 11500 27620 11512
rect 27672 11500 27678 11552
rect 28721 11543 28779 11549
rect 28721 11509 28733 11543
rect 28767 11540 28779 11543
rect 29362 11540 29368 11552
rect 28767 11512 29368 11540
rect 28767 11509 28779 11512
rect 28721 11503 28779 11509
rect 29362 11500 29368 11512
rect 29420 11500 29426 11552
rect 30469 11543 30527 11549
rect 30469 11509 30481 11543
rect 30515 11540 30527 11543
rect 31478 11540 31484 11552
rect 30515 11512 31484 11540
rect 30515 11509 30527 11512
rect 30469 11503 30527 11509
rect 31478 11500 31484 11512
rect 31536 11500 31542 11552
rect 33778 11540 33784 11552
rect 33739 11512 33784 11540
rect 33778 11500 33784 11512
rect 33836 11500 33842 11552
rect 33965 11543 34023 11549
rect 33965 11509 33977 11543
rect 34011 11540 34023 11543
rect 34698 11540 34704 11552
rect 34011 11512 34704 11540
rect 34011 11509 34023 11512
rect 33965 11503 34023 11509
rect 34698 11500 34704 11512
rect 34756 11500 34762 11552
rect 34793 11543 34851 11549
rect 34793 11509 34805 11543
rect 34839 11540 34851 11543
rect 35434 11540 35440 11552
rect 34839 11512 35440 11540
rect 34839 11509 34851 11512
rect 34793 11503 34851 11509
rect 35434 11500 35440 11512
rect 35492 11500 35498 11552
rect 39298 11540 39304 11552
rect 39259 11512 39304 11540
rect 39298 11500 39304 11512
rect 39356 11500 39362 11552
rect 39850 11500 39856 11552
rect 39908 11540 39914 11552
rect 46032 11540 46060 11639
rect 48590 11636 48596 11688
rect 48648 11676 48654 11688
rect 48777 11679 48835 11685
rect 48777 11676 48789 11679
rect 48648 11648 48789 11676
rect 48648 11636 48654 11648
rect 48777 11645 48789 11648
rect 48823 11645 48835 11679
rect 48777 11639 48835 11645
rect 48869 11679 48927 11685
rect 48869 11645 48881 11679
rect 48915 11676 48927 11679
rect 48958 11676 48964 11688
rect 48915 11648 48964 11676
rect 48915 11645 48927 11648
rect 48869 11639 48927 11645
rect 48958 11636 48964 11648
rect 49016 11636 49022 11688
rect 56594 11676 56600 11688
rect 56555 11648 56600 11676
rect 56594 11636 56600 11648
rect 56652 11636 56658 11688
rect 39908 11512 46060 11540
rect 46385 11543 46443 11549
rect 39908 11500 39914 11512
rect 46385 11509 46397 11543
rect 46431 11540 46443 11543
rect 47946 11540 47952 11552
rect 46431 11512 47952 11540
rect 46431 11509 46443 11512
rect 46385 11503 46443 11509
rect 47946 11500 47952 11512
rect 48004 11500 48010 11552
rect 53282 11540 53288 11552
rect 53243 11512 53288 11540
rect 53282 11500 53288 11512
rect 53340 11500 53346 11552
rect 1104 11450 58880 11472
rect 1104 11398 4214 11450
rect 4266 11398 4278 11450
rect 4330 11398 4342 11450
rect 4394 11398 4406 11450
rect 4458 11398 4470 11450
rect 4522 11398 34934 11450
rect 34986 11398 34998 11450
rect 35050 11398 35062 11450
rect 35114 11398 35126 11450
rect 35178 11398 35190 11450
rect 35242 11398 58880 11450
rect 1104 11376 58880 11398
rect 2866 11336 2872 11348
rect 2827 11308 2872 11336
rect 2866 11296 2872 11308
rect 2924 11296 2930 11348
rect 3602 11296 3608 11348
rect 3660 11336 3666 11348
rect 3789 11339 3847 11345
rect 3789 11336 3801 11339
rect 3660 11308 3801 11336
rect 3660 11296 3666 11308
rect 3789 11305 3801 11308
rect 3835 11305 3847 11339
rect 22278 11336 22284 11348
rect 22239 11308 22284 11336
rect 3789 11299 3847 11305
rect 22278 11296 22284 11308
rect 22336 11296 22342 11348
rect 22370 11296 22376 11348
rect 22428 11336 22434 11348
rect 25317 11339 25375 11345
rect 25317 11336 25329 11339
rect 22428 11308 25329 11336
rect 22428 11296 22434 11308
rect 25317 11305 25329 11308
rect 25363 11305 25375 11339
rect 25317 11299 25375 11305
rect 25590 11296 25596 11348
rect 25648 11336 25654 11348
rect 30374 11336 30380 11348
rect 25648 11308 30380 11336
rect 25648 11296 25654 11308
rect 30374 11296 30380 11308
rect 30432 11296 30438 11348
rect 41046 11336 41052 11348
rect 35176 11308 41052 11336
rect 16758 11268 16764 11280
rect 16592 11240 16764 11268
rect 3878 11200 3884 11212
rect 2976 11172 3884 11200
rect 2866 11092 2872 11144
rect 2924 11132 2930 11144
rect 2976 11141 3004 11172
rect 3878 11160 3884 11172
rect 3936 11160 3942 11212
rect 11882 11160 11888 11212
rect 11940 11200 11946 11212
rect 11977 11203 12035 11209
rect 11977 11200 11989 11203
rect 11940 11172 11989 11200
rect 11940 11160 11946 11172
rect 11977 11169 11989 11172
rect 12023 11169 12035 11203
rect 15657 11203 15715 11209
rect 15657 11200 15669 11203
rect 11977 11163 12035 11169
rect 14660 11172 15669 11200
rect 2961 11135 3019 11141
rect 2961 11132 2973 11135
rect 2924 11104 2973 11132
rect 2924 11092 2930 11104
rect 2961 11101 2973 11104
rect 3007 11101 3019 11135
rect 2961 11095 3019 11101
rect 3789 11135 3847 11141
rect 3789 11101 3801 11135
rect 3835 11101 3847 11135
rect 3789 11095 3847 11101
rect 3973 11135 4031 11141
rect 3973 11101 3985 11135
rect 4019 11132 4031 11135
rect 4062 11132 4068 11144
rect 4019 11104 4068 11132
rect 4019 11101 4031 11104
rect 3973 11095 4031 11101
rect 3145 11067 3203 11073
rect 3145 11033 3157 11067
rect 3191 11033 3203 11067
rect 3804 11064 3832 11095
rect 4062 11092 4068 11104
rect 4120 11092 4126 11144
rect 12161 11135 12219 11141
rect 12161 11101 12173 11135
rect 12207 11132 12219 11135
rect 12342 11132 12348 11144
rect 12207 11104 12348 11132
rect 12207 11101 12219 11104
rect 12161 11095 12219 11101
rect 12342 11092 12348 11104
rect 12400 11092 12406 11144
rect 14660 11141 14688 11172
rect 15657 11169 15669 11172
rect 15703 11169 15715 11203
rect 16390 11200 16396 11212
rect 15657 11163 15715 11169
rect 15948 11172 16396 11200
rect 14645 11135 14703 11141
rect 14645 11101 14657 11135
rect 14691 11101 14703 11135
rect 14645 11095 14703 11101
rect 14921 11135 14979 11141
rect 14921 11101 14933 11135
rect 14967 11132 14979 11135
rect 15102 11132 15108 11144
rect 14967 11104 15108 11132
rect 14967 11101 14979 11104
rect 14921 11095 14979 11101
rect 15102 11092 15108 11104
rect 15160 11092 15166 11144
rect 15838 11132 15844 11144
rect 15799 11104 15844 11132
rect 15838 11092 15844 11104
rect 15896 11092 15902 11144
rect 3804 11036 4108 11064
rect 3145 11027 3203 11033
rect 3160 10996 3188 11027
rect 4080 11008 4108 11036
rect 14274 11024 14280 11076
rect 14332 11064 14338 11076
rect 14461 11067 14519 11073
rect 14461 11064 14473 11067
rect 14332 11036 14473 11064
rect 14332 11024 14338 11036
rect 14461 11033 14473 11036
rect 14507 11033 14519 11067
rect 14461 11027 14519 11033
rect 14829 11067 14887 11073
rect 14829 11033 14841 11067
rect 14875 11064 14887 11067
rect 15194 11064 15200 11076
rect 14875 11036 15200 11064
rect 14875 11033 14887 11036
rect 14829 11027 14887 11033
rect 15194 11024 15200 11036
rect 15252 11064 15258 11076
rect 15948 11064 15976 11172
rect 16390 11160 16396 11172
rect 16448 11160 16454 11212
rect 16114 11132 16120 11144
rect 16075 11104 16120 11132
rect 16114 11092 16120 11104
rect 16172 11092 16178 11144
rect 16592 11141 16620 11240
rect 16758 11228 16764 11240
rect 16816 11268 16822 11280
rect 16816 11240 20024 11268
rect 16816 11228 16822 11240
rect 17586 11200 17592 11212
rect 17499 11172 17592 11200
rect 17586 11160 17592 11172
rect 17644 11200 17650 11212
rect 19334 11200 19340 11212
rect 17644 11172 19340 11200
rect 17644 11160 17650 11172
rect 19334 11160 19340 11172
rect 19392 11160 19398 11212
rect 19996 11144 20024 11240
rect 24210 11228 24216 11280
rect 24268 11268 24274 11280
rect 30653 11271 30711 11277
rect 30653 11268 30665 11271
rect 24268 11240 30665 11268
rect 24268 11228 24274 11240
rect 30653 11237 30665 11240
rect 30699 11268 30711 11271
rect 33965 11271 34023 11277
rect 30699 11240 31248 11268
rect 30699 11237 30711 11240
rect 30653 11231 30711 11237
rect 20990 11160 20996 11212
rect 21048 11200 21054 11212
rect 26510 11200 26516 11212
rect 21048 11172 22140 11200
rect 21048 11160 21054 11172
rect 16577 11135 16635 11141
rect 16577 11132 16589 11135
rect 16224 11104 16589 11132
rect 15252 11036 15976 11064
rect 16025 11067 16083 11073
rect 15252 11024 15258 11036
rect 16025 11033 16037 11067
rect 16071 11064 16083 11067
rect 16224 11064 16252 11104
rect 16577 11101 16589 11104
rect 16623 11101 16635 11135
rect 16577 11095 16635 11101
rect 16666 11092 16672 11144
rect 16724 11132 16730 11144
rect 16945 11135 17003 11141
rect 16945 11132 16957 11135
rect 16724 11104 16957 11132
rect 16724 11092 16730 11104
rect 16945 11101 16957 11104
rect 16991 11132 17003 11135
rect 17773 11135 17831 11141
rect 17773 11132 17785 11135
rect 16991 11104 17785 11132
rect 16991 11101 17003 11104
rect 16945 11095 17003 11101
rect 17773 11101 17785 11104
rect 17819 11132 17831 11135
rect 17862 11132 17868 11144
rect 17819 11104 17868 11132
rect 17819 11101 17831 11104
rect 17773 11095 17831 11101
rect 17862 11092 17868 11104
rect 17920 11092 17926 11144
rect 19978 11092 19984 11144
rect 20036 11132 20042 11144
rect 21082 11132 21088 11144
rect 20036 11104 21088 11132
rect 20036 11092 20042 11104
rect 21082 11092 21088 11104
rect 21140 11132 21146 11144
rect 22112 11141 22140 11172
rect 25516 11172 26516 11200
rect 21729 11135 21787 11141
rect 21729 11132 21741 11135
rect 21140 11104 21741 11132
rect 21140 11092 21146 11104
rect 21729 11101 21741 11104
rect 21775 11101 21787 11135
rect 21729 11095 21787 11101
rect 22097 11135 22155 11141
rect 22097 11101 22109 11135
rect 22143 11132 22155 11135
rect 22833 11135 22891 11141
rect 22833 11132 22845 11135
rect 22143 11104 22845 11132
rect 22143 11101 22155 11104
rect 22097 11095 22155 11101
rect 22833 11101 22845 11104
rect 22879 11101 22891 11135
rect 25314 11132 25320 11144
rect 25275 11104 25320 11132
rect 22833 11095 22891 11101
rect 25314 11092 25320 11104
rect 25372 11092 25378 11144
rect 25516 11141 25544 11172
rect 26510 11160 26516 11172
rect 26568 11200 26574 11212
rect 29178 11200 29184 11212
rect 26568 11172 29184 11200
rect 26568 11160 26574 11172
rect 29178 11160 29184 11172
rect 29236 11160 29242 11212
rect 29822 11160 29828 11212
rect 29880 11160 29886 11212
rect 31220 11209 31248 11240
rect 33965 11237 33977 11271
rect 34011 11268 34023 11271
rect 34011 11240 34836 11268
rect 34011 11237 34023 11240
rect 33965 11231 34023 11237
rect 31205 11203 31263 11209
rect 31205 11169 31217 11203
rect 31251 11200 31263 11203
rect 31938 11200 31944 11212
rect 31251 11172 31944 11200
rect 31251 11169 31263 11172
rect 31205 11163 31263 11169
rect 31938 11160 31944 11172
rect 31996 11160 32002 11212
rect 25501 11135 25559 11141
rect 25501 11101 25513 11135
rect 25547 11101 25559 11135
rect 25501 11095 25559 11101
rect 25593 11135 25651 11141
rect 25593 11101 25605 11135
rect 25639 11132 25651 11135
rect 25682 11132 25688 11144
rect 25639 11104 25688 11132
rect 25639 11101 25651 11104
rect 25593 11095 25651 11101
rect 25682 11092 25688 11104
rect 25740 11132 25746 11144
rect 27525 11135 27583 11141
rect 25740 11104 27476 11132
rect 25740 11092 25746 11104
rect 16071 11036 16252 11064
rect 16071 11033 16083 11036
rect 16025 11027 16083 11033
rect 16298 11024 16304 11076
rect 16356 11064 16362 11076
rect 16761 11067 16819 11073
rect 16761 11064 16773 11067
rect 16356 11036 16773 11064
rect 16356 11024 16362 11036
rect 16761 11033 16773 11036
rect 16807 11033 16819 11067
rect 16761 11027 16819 11033
rect 16853 11067 16911 11073
rect 16853 11033 16865 11067
rect 16899 11064 16911 11067
rect 20530 11064 20536 11076
rect 16899 11036 20536 11064
rect 16899 11033 16911 11036
rect 16853 11027 16911 11033
rect 20530 11024 20536 11036
rect 20588 11024 20594 11076
rect 21910 11064 21916 11076
rect 21871 11036 21916 11064
rect 21910 11024 21916 11036
rect 21968 11024 21974 11076
rect 22005 11067 22063 11073
rect 22005 11033 22017 11067
rect 22051 11064 22063 11067
rect 23658 11064 23664 11076
rect 22051 11036 23664 11064
rect 22051 11033 22063 11036
rect 22005 11027 22063 11033
rect 23658 11024 23664 11036
rect 23716 11024 23722 11076
rect 27448 11064 27476 11104
rect 27525 11101 27537 11135
rect 27571 11132 27583 11135
rect 27614 11132 27620 11144
rect 27571 11104 27620 11132
rect 27571 11101 27583 11104
rect 27525 11095 27583 11101
rect 27614 11092 27620 11104
rect 27672 11092 27678 11144
rect 27798 11132 27804 11144
rect 27759 11104 27804 11132
rect 27798 11092 27804 11104
rect 27856 11092 27862 11144
rect 27893 11135 27951 11141
rect 27893 11101 27905 11135
rect 27939 11132 27951 11135
rect 27982 11132 27988 11144
rect 27939 11104 27988 11132
rect 27939 11101 27951 11104
rect 27893 11095 27951 11101
rect 27982 11092 27988 11104
rect 28040 11092 28046 11144
rect 29840 11132 29868 11160
rect 34808 11144 34836 11240
rect 35176 11209 35204 11308
rect 41046 11296 41052 11308
rect 41104 11296 41110 11348
rect 42337 11339 42395 11345
rect 42337 11305 42349 11339
rect 42383 11336 42395 11339
rect 44910 11336 44916 11348
rect 42383 11308 44916 11336
rect 42383 11305 42395 11308
rect 42337 11299 42395 11305
rect 44910 11296 44916 11308
rect 44968 11296 44974 11348
rect 45830 11296 45836 11348
rect 45888 11336 45894 11348
rect 46109 11339 46167 11345
rect 46109 11336 46121 11339
rect 45888 11308 46121 11336
rect 45888 11296 45894 11308
rect 46109 11305 46121 11308
rect 46155 11305 46167 11339
rect 46109 11299 46167 11305
rect 46658 11296 46664 11348
rect 46716 11336 46722 11348
rect 47670 11336 47676 11348
rect 46716 11308 47676 11336
rect 46716 11296 46722 11308
rect 47670 11296 47676 11308
rect 47728 11296 47734 11348
rect 35802 11228 35808 11280
rect 35860 11268 35866 11280
rect 35989 11271 36047 11277
rect 35989 11268 36001 11271
rect 35860 11240 36001 11268
rect 35860 11228 35866 11240
rect 35989 11237 36001 11240
rect 36035 11237 36047 11271
rect 35989 11231 36047 11237
rect 36170 11228 36176 11280
rect 36228 11228 36234 11280
rect 39117 11271 39175 11277
rect 39117 11237 39129 11271
rect 39163 11268 39175 11271
rect 39163 11240 41414 11268
rect 39163 11237 39175 11240
rect 39117 11231 39175 11237
rect 35161 11203 35219 11209
rect 35161 11169 35173 11203
rect 35207 11169 35219 11203
rect 35342 11200 35348 11212
rect 35161 11163 35219 11169
rect 35268 11172 35348 11200
rect 30282 11132 30288 11144
rect 29840 11104 30288 11132
rect 30282 11092 30288 11104
rect 30340 11132 30346 11144
rect 31297 11135 31355 11141
rect 31297 11132 31309 11135
rect 30340 11104 31309 11132
rect 30340 11092 30346 11104
rect 31297 11101 31309 11104
rect 31343 11101 31355 11135
rect 31478 11132 31484 11144
rect 31439 11104 31484 11132
rect 31297 11095 31355 11101
rect 31478 11092 31484 11104
rect 31536 11092 31542 11144
rect 33686 11132 33692 11144
rect 33647 11104 33692 11132
rect 33686 11092 33692 11104
rect 33744 11092 33750 11144
rect 33778 11092 33784 11144
rect 33836 11132 33842 11144
rect 34790 11132 34796 11144
rect 33836 11104 33881 11132
rect 34751 11104 34796 11132
rect 33836 11092 33842 11104
rect 34790 11092 34796 11104
rect 34848 11092 34854 11144
rect 35268 11141 35296 11172
rect 35342 11160 35348 11172
rect 35400 11160 35406 11212
rect 36188 11200 36216 11228
rect 39022 11200 39028 11212
rect 36004 11172 36216 11200
rect 38764 11172 39028 11200
rect 34977 11135 35035 11141
rect 34977 11101 34989 11135
rect 35023 11101 35035 11135
rect 34977 11095 35035 11101
rect 35253 11135 35311 11141
rect 35253 11101 35265 11135
rect 35299 11101 35311 11135
rect 35434 11132 35440 11144
rect 35395 11104 35440 11132
rect 35253 11095 35311 11101
rect 27709 11067 27767 11073
rect 27709 11064 27721 11067
rect 27448 11036 27721 11064
rect 27709 11033 27721 11036
rect 27755 11033 27767 11067
rect 27709 11027 27767 11033
rect 31665 11067 31723 11073
rect 31665 11033 31677 11067
rect 31711 11064 31723 11067
rect 32674 11064 32680 11076
rect 31711 11036 32680 11064
rect 31711 11033 31723 11036
rect 31665 11027 31723 11033
rect 32674 11024 32680 11036
rect 32732 11024 32738 11076
rect 33594 11024 33600 11076
rect 33652 11064 33658 11076
rect 33965 11067 34023 11073
rect 33965 11064 33977 11067
rect 33652 11036 33977 11064
rect 33652 11024 33658 11036
rect 33965 11033 33977 11036
rect 34011 11064 34023 11067
rect 34011 11036 34652 11064
rect 34011 11033 34023 11036
rect 33965 11027 34023 11033
rect 3786 10996 3792 11008
rect 3160 10968 3792 10996
rect 3786 10956 3792 10968
rect 3844 10956 3850 11008
rect 4062 10956 4068 11008
rect 4120 10956 4126 11008
rect 9677 10999 9735 11005
rect 9677 10965 9689 10999
rect 9723 10996 9735 10999
rect 10134 10996 10140 11008
rect 9723 10968 10140 10996
rect 9723 10965 9735 10968
rect 9677 10959 9735 10965
rect 10134 10956 10140 10968
rect 10192 10956 10198 11008
rect 12342 10996 12348 11008
rect 12303 10968 12348 10996
rect 12342 10956 12348 10968
rect 12400 10956 12406 11008
rect 16942 10956 16948 11008
rect 17000 10996 17006 11008
rect 17129 10999 17187 11005
rect 17129 10996 17141 10999
rect 17000 10968 17141 10996
rect 17000 10956 17006 10968
rect 17129 10965 17141 10968
rect 17175 10965 17187 10999
rect 22922 10996 22928 11008
rect 22883 10968 22928 10996
rect 17129 10959 17187 10965
rect 22922 10956 22928 10968
rect 22980 10956 22986 11008
rect 28074 10996 28080 11008
rect 28035 10968 28080 10996
rect 28074 10956 28080 10968
rect 28132 10956 28138 11008
rect 34624 10996 34652 11036
rect 34698 11024 34704 11076
rect 34756 11064 34762 11076
rect 34992 11064 35020 11095
rect 35434 11092 35440 11104
rect 35492 11092 35498 11144
rect 36004 11141 36032 11172
rect 35989 11135 36047 11141
rect 35989 11101 36001 11135
rect 36035 11101 36047 11135
rect 35989 11095 36047 11101
rect 36004 11064 36032 11095
rect 36078 11092 36084 11144
rect 36136 11132 36142 11144
rect 36173 11135 36231 11141
rect 36173 11132 36185 11135
rect 36136 11104 36185 11132
rect 36136 11092 36142 11104
rect 36173 11101 36185 11104
rect 36219 11101 36231 11135
rect 38562 11132 38568 11144
rect 38523 11104 38568 11132
rect 36173 11095 36231 11101
rect 38562 11092 38568 11104
rect 38620 11092 38626 11144
rect 38764 11141 38792 11172
rect 39022 11160 39028 11172
rect 39080 11160 39086 11212
rect 40310 11200 40316 11212
rect 40271 11172 40316 11200
rect 40310 11160 40316 11172
rect 40368 11160 40374 11212
rect 38749 11135 38807 11141
rect 38749 11101 38761 11135
rect 38795 11101 38807 11135
rect 38930 11132 38936 11144
rect 38891 11104 38936 11132
rect 38749 11095 38807 11101
rect 38930 11092 38936 11104
rect 38988 11092 38994 11144
rect 41386 11132 41414 11240
rect 43162 11228 43168 11280
rect 43220 11228 43226 11280
rect 43180 11200 43208 11228
rect 45848 11200 45876 11296
rect 45922 11228 45928 11280
rect 45980 11268 45986 11280
rect 46293 11271 46351 11277
rect 46293 11268 46305 11271
rect 45980 11240 46305 11268
rect 45980 11228 45986 11240
rect 46293 11237 46305 11240
rect 46339 11268 46351 11271
rect 48590 11268 48596 11280
rect 46339 11240 48596 11268
rect 46339 11237 46351 11240
rect 46293 11231 46351 11237
rect 48590 11228 48596 11240
rect 48648 11228 48654 11280
rect 52730 11268 52736 11280
rect 52691 11240 52736 11268
rect 52730 11228 52736 11240
rect 52788 11228 52794 11280
rect 56962 11228 56968 11280
rect 57020 11268 57026 11280
rect 57020 11240 57744 11268
rect 57020 11228 57026 11240
rect 43180 11172 43484 11200
rect 45848 11172 46612 11200
rect 42153 11135 42211 11141
rect 42153 11132 42165 11135
rect 41386 11104 42165 11132
rect 42153 11101 42165 11104
rect 42199 11101 42211 11135
rect 42334 11132 42340 11144
rect 42295 11104 42340 11132
rect 42153 11095 42211 11101
rect 42334 11092 42340 11104
rect 42392 11092 42398 11144
rect 43070 11092 43076 11144
rect 43128 11132 43134 11144
rect 43456 11141 43484 11172
rect 43165 11135 43223 11141
rect 43165 11132 43177 11135
rect 43128 11104 43177 11132
rect 43128 11092 43134 11104
rect 43165 11101 43177 11104
rect 43211 11101 43223 11135
rect 43165 11095 43223 11101
rect 43441 11135 43499 11141
rect 43441 11101 43453 11135
rect 43487 11101 43499 11135
rect 43441 11095 43499 11101
rect 43625 11135 43683 11141
rect 43625 11101 43637 11135
rect 43671 11132 43683 11135
rect 45738 11132 45744 11144
rect 43671 11104 45744 11132
rect 43671 11101 43683 11104
rect 43625 11095 43683 11101
rect 45738 11092 45744 11104
rect 45796 11132 45802 11144
rect 46584 11132 46612 11172
rect 47670 11160 47676 11212
rect 47728 11200 47734 11212
rect 53282 11200 53288 11212
rect 47728 11172 48544 11200
rect 53243 11172 53288 11200
rect 47728 11160 47734 11172
rect 48516 11141 48544 11172
rect 53282 11160 53288 11172
rect 53340 11160 53346 11212
rect 54018 11200 54024 11212
rect 53979 11172 54024 11200
rect 54018 11160 54024 11172
rect 54076 11160 54082 11212
rect 57606 11200 57612 11212
rect 56888 11172 57612 11200
rect 48225 11135 48283 11141
rect 48225 11132 48237 11135
rect 45796 11104 46060 11132
rect 46584 11104 48237 11132
rect 45796 11092 45802 11104
rect 34756 11036 35020 11064
rect 35084 11036 36032 11064
rect 34756 11024 34762 11036
rect 35084 10996 35112 11036
rect 38470 11024 38476 11076
rect 38528 11064 38534 11076
rect 38841 11067 38899 11073
rect 38841 11064 38853 11067
rect 38528 11036 38853 11064
rect 38528 11024 38534 11036
rect 38841 11033 38853 11036
rect 38887 11064 38899 11067
rect 39850 11064 39856 11076
rect 38887 11036 39856 11064
rect 38887 11033 38899 11036
rect 38841 11027 38899 11033
rect 39850 11024 39856 11036
rect 39908 11024 39914 11076
rect 43257 11067 43315 11073
rect 43257 11033 43269 11067
rect 43303 11064 43315 11067
rect 43806 11064 43812 11076
rect 43303 11036 43812 11064
rect 43303 11033 43315 11036
rect 43257 11027 43315 11033
rect 43806 11024 43812 11036
rect 43864 11064 43870 11076
rect 43864 11036 45324 11064
rect 43864 11024 43870 11036
rect 34624 10968 35112 10996
rect 35526 10956 35532 11008
rect 35584 10996 35590 11008
rect 41414 10996 41420 11008
rect 35584 10968 41420 10996
rect 35584 10956 35590 10968
rect 41414 10956 41420 10968
rect 41472 10956 41478 11008
rect 45296 10996 45324 11036
rect 45370 11024 45376 11076
rect 45428 11064 45434 11076
rect 45925 11067 45983 11073
rect 45925 11064 45937 11067
rect 45428 11036 45937 11064
rect 45428 11024 45434 11036
rect 45925 11033 45937 11036
rect 45971 11033 45983 11067
rect 46032 11064 46060 11104
rect 48225 11101 48237 11104
rect 48271 11101 48283 11135
rect 48225 11095 48283 11101
rect 48501 11135 48559 11141
rect 48501 11101 48513 11135
rect 48547 11101 48559 11135
rect 48501 11095 48559 11101
rect 46125 11067 46183 11073
rect 46125 11064 46137 11067
rect 46032 11036 46137 11064
rect 45925 11027 45983 11033
rect 46125 11033 46137 11036
rect 46171 11033 46183 11067
rect 48240 11064 48268 11095
rect 48590 11092 48596 11144
rect 48648 11132 48654 11144
rect 49145 11135 49203 11141
rect 49145 11132 49157 11135
rect 48648 11104 49157 11132
rect 48648 11092 48654 11104
rect 49145 11101 49157 11104
rect 49191 11101 49203 11135
rect 49145 11095 49203 11101
rect 49329 11135 49387 11141
rect 49329 11101 49341 11135
rect 49375 11101 49387 11135
rect 49329 11095 49387 11101
rect 48682 11064 48688 11076
rect 46125 11027 46183 11033
rect 46216 11036 48176 11064
rect 48240 11036 48544 11064
rect 48643 11036 48688 11064
rect 46216 10996 46244 11036
rect 45296 10968 46244 10996
rect 48148 10996 48176 11036
rect 48317 10999 48375 11005
rect 48317 10996 48329 10999
rect 48148 10968 48329 10996
rect 48317 10965 48329 10968
rect 48363 10996 48375 10999
rect 48406 10996 48412 11008
rect 48363 10968 48412 10996
rect 48363 10965 48375 10968
rect 48317 10959 48375 10965
rect 48406 10956 48412 10968
rect 48464 10956 48470 11008
rect 48516 10996 48544 11036
rect 48682 11024 48688 11036
rect 48740 11024 48746 11076
rect 49344 11064 49372 11095
rect 51534 11092 51540 11144
rect 51592 11132 51598 11144
rect 51721 11135 51779 11141
rect 51721 11132 51733 11135
rect 51592 11104 51733 11132
rect 51592 11092 51598 11104
rect 51721 11101 51733 11104
rect 51767 11101 51779 11135
rect 53006 11132 53012 11144
rect 52967 11104 53012 11132
rect 51721 11095 51779 11101
rect 53006 11092 53012 11104
rect 53064 11092 53070 11144
rect 53745 11135 53803 11141
rect 53745 11101 53757 11135
rect 53791 11132 53803 11135
rect 53834 11132 53840 11144
rect 53791 11104 53840 11132
rect 53791 11101 53803 11104
rect 53745 11095 53803 11101
rect 53834 11092 53840 11104
rect 53892 11092 53898 11144
rect 54662 11092 54668 11144
rect 54720 11132 54726 11144
rect 56229 11135 56287 11141
rect 56229 11132 56241 11135
rect 54720 11104 56241 11132
rect 54720 11092 54726 11104
rect 56229 11101 56241 11104
rect 56275 11101 56287 11135
rect 56229 11095 56287 11101
rect 56413 11135 56471 11141
rect 56413 11101 56425 11135
rect 56459 11132 56471 11135
rect 56502 11132 56508 11144
rect 56459 11104 56508 11132
rect 56459 11101 56471 11104
rect 56413 11095 56471 11101
rect 56502 11092 56508 11104
rect 56560 11092 56566 11144
rect 56888 11141 56916 11172
rect 57606 11160 57612 11172
rect 57664 11160 57670 11212
rect 56689 11135 56747 11141
rect 56689 11101 56701 11135
rect 56735 11101 56747 11135
rect 56689 11095 56747 11101
rect 56873 11135 56931 11141
rect 56873 11101 56885 11135
rect 56919 11101 56931 11135
rect 56873 11095 56931 11101
rect 57333 11135 57391 11141
rect 57333 11101 57345 11135
rect 57379 11132 57391 11135
rect 57422 11132 57428 11144
rect 57379 11104 57428 11132
rect 57379 11101 57391 11104
rect 57333 11095 57391 11101
rect 48792 11036 49372 11064
rect 56704 11064 56732 11095
rect 57422 11092 57428 11104
rect 57480 11092 57486 11144
rect 57517 11135 57575 11141
rect 57517 11101 57529 11135
rect 57563 11132 57575 11135
rect 57716 11132 57744 11240
rect 57977 11135 58035 11141
rect 57977 11132 57989 11135
rect 57563 11104 57989 11132
rect 57563 11101 57575 11104
rect 57517 11095 57575 11101
rect 57977 11101 57989 11104
rect 58023 11101 58035 11135
rect 57977 11095 58035 11101
rect 58069 11067 58127 11073
rect 58069 11064 58081 11067
rect 56704 11036 58081 11064
rect 48792 10996 48820 11036
rect 58069 11033 58081 11036
rect 58115 11033 58127 11067
rect 58069 11027 58127 11033
rect 48516 10968 48820 10996
rect 48958 10956 48964 11008
rect 49016 10996 49022 11008
rect 49145 10999 49203 11005
rect 49145 10996 49157 10999
rect 49016 10968 49157 10996
rect 49016 10956 49022 10968
rect 49145 10965 49157 10968
rect 49191 10965 49203 10999
rect 51810 10996 51816 11008
rect 51771 10968 51816 10996
rect 49145 10959 49203 10965
rect 51810 10956 51816 10968
rect 51868 10956 51874 11008
rect 56962 10956 56968 11008
rect 57020 10996 57026 11008
rect 57425 10999 57483 11005
rect 57425 10996 57437 10999
rect 57020 10968 57437 10996
rect 57020 10956 57026 10968
rect 57425 10965 57437 10968
rect 57471 10965 57483 10999
rect 57425 10959 57483 10965
rect 1104 10906 58880 10928
rect 1104 10854 19574 10906
rect 19626 10854 19638 10906
rect 19690 10854 19702 10906
rect 19754 10854 19766 10906
rect 19818 10854 19830 10906
rect 19882 10854 50294 10906
rect 50346 10854 50358 10906
rect 50410 10854 50422 10906
rect 50474 10854 50486 10906
rect 50538 10854 50550 10906
rect 50602 10854 58880 10906
rect 1104 10832 58880 10854
rect 2501 10795 2559 10801
rect 2501 10761 2513 10795
rect 2547 10792 2559 10795
rect 2774 10792 2780 10804
rect 2547 10764 2780 10792
rect 2547 10761 2559 10764
rect 2501 10755 2559 10761
rect 2774 10752 2780 10764
rect 2832 10752 2838 10804
rect 3878 10752 3884 10804
rect 3936 10792 3942 10804
rect 4065 10795 4123 10801
rect 4065 10792 4077 10795
rect 3936 10764 4077 10792
rect 3936 10752 3942 10764
rect 4065 10761 4077 10764
rect 4111 10761 4123 10795
rect 6362 10792 6368 10804
rect 6323 10764 6368 10792
rect 4065 10755 4123 10761
rect 6362 10752 6368 10764
rect 6420 10752 6426 10804
rect 9125 10795 9183 10801
rect 9125 10761 9137 10795
rect 9171 10792 9183 10795
rect 9306 10792 9312 10804
rect 9171 10764 9312 10792
rect 9171 10761 9183 10764
rect 9125 10755 9183 10761
rect 9306 10752 9312 10764
rect 9364 10752 9370 10804
rect 10042 10792 10048 10804
rect 10003 10764 10048 10792
rect 10042 10752 10048 10764
rect 10100 10752 10106 10804
rect 14369 10795 14427 10801
rect 14369 10761 14381 10795
rect 14415 10792 14427 10795
rect 15194 10792 15200 10804
rect 14415 10764 15200 10792
rect 14415 10761 14427 10764
rect 14369 10755 14427 10761
rect 15194 10752 15200 10764
rect 15252 10752 15258 10804
rect 16114 10752 16120 10804
rect 16172 10792 16178 10804
rect 17034 10792 17040 10804
rect 16172 10764 17040 10792
rect 16172 10752 16178 10764
rect 17034 10752 17040 10764
rect 17092 10752 17098 10804
rect 24762 10792 24768 10804
rect 23032 10764 24768 10792
rect 11793 10727 11851 10733
rect 9324 10696 10180 10724
rect 1394 10656 1400 10668
rect 1355 10628 1400 10656
rect 1394 10616 1400 10628
rect 1452 10616 1458 10668
rect 3329 10659 3387 10665
rect 3329 10625 3341 10659
rect 3375 10656 3387 10659
rect 3694 10656 3700 10668
rect 3375 10628 3700 10656
rect 3375 10625 3387 10628
rect 3329 10619 3387 10625
rect 3694 10616 3700 10628
rect 3752 10616 3758 10668
rect 4062 10616 4068 10668
rect 4120 10656 4126 10668
rect 4249 10659 4307 10665
rect 4249 10656 4261 10659
rect 4120 10628 4261 10656
rect 4120 10616 4126 10628
rect 4249 10625 4261 10628
rect 4295 10625 4307 10659
rect 4249 10619 4307 10625
rect 6549 10659 6607 10665
rect 6549 10625 6561 10659
rect 6595 10656 6607 10659
rect 6822 10656 6828 10668
rect 6595 10628 6828 10656
rect 6595 10625 6607 10628
rect 6549 10619 6607 10625
rect 6822 10616 6828 10628
rect 6880 10616 6886 10668
rect 9324 10665 9352 10696
rect 10152 10668 10180 10696
rect 11793 10693 11805 10727
rect 11839 10724 11851 10727
rect 15102 10724 15108 10736
rect 11839 10696 13216 10724
rect 15063 10696 15108 10724
rect 11839 10693 11851 10696
rect 11793 10687 11851 10693
rect 13188 10668 13216 10696
rect 15102 10684 15108 10696
rect 15160 10724 15166 10736
rect 15565 10727 15623 10733
rect 15565 10724 15577 10727
rect 15160 10696 15577 10724
rect 15160 10684 15166 10696
rect 15565 10693 15577 10696
rect 15611 10693 15623 10727
rect 15565 10687 15623 10693
rect 19429 10727 19487 10733
rect 19429 10693 19441 10727
rect 19475 10724 19487 10727
rect 20070 10724 20076 10736
rect 19475 10696 20076 10724
rect 19475 10693 19487 10696
rect 19429 10687 19487 10693
rect 20070 10684 20076 10696
rect 20128 10684 20134 10736
rect 23032 10733 23060 10764
rect 24762 10752 24768 10764
rect 24820 10792 24826 10804
rect 27430 10792 27436 10804
rect 24820 10764 26188 10792
rect 27343 10764 27436 10792
rect 24820 10752 24826 10764
rect 23017 10727 23075 10733
rect 23017 10693 23029 10727
rect 23063 10693 23075 10727
rect 23017 10687 23075 10693
rect 23109 10727 23167 10733
rect 23109 10693 23121 10727
rect 23155 10724 23167 10727
rect 24302 10724 24308 10736
rect 23155 10696 24308 10724
rect 23155 10693 23167 10696
rect 23109 10687 23167 10693
rect 24302 10684 24308 10696
rect 24360 10684 24366 10736
rect 24394 10684 24400 10736
rect 24452 10724 24458 10736
rect 26160 10733 26188 10764
rect 27430 10752 27436 10764
rect 27488 10792 27494 10804
rect 27488 10764 28994 10792
rect 27488 10752 27494 10764
rect 25317 10727 25375 10733
rect 25317 10724 25329 10727
rect 24452 10696 25329 10724
rect 24452 10684 24458 10696
rect 25317 10693 25329 10696
rect 25363 10693 25375 10727
rect 25317 10687 25375 10693
rect 26145 10727 26203 10733
rect 26145 10693 26157 10727
rect 26191 10693 26203 10727
rect 26145 10687 26203 10693
rect 9309 10659 9367 10665
rect 9309 10625 9321 10659
rect 9355 10625 9367 10659
rect 9953 10659 10011 10665
rect 9953 10656 9965 10659
rect 9309 10619 9367 10625
rect 9508 10628 9965 10656
rect 9508 10600 9536 10628
rect 9953 10625 9965 10628
rect 9999 10625 10011 10659
rect 9953 10619 10011 10625
rect 10134 10616 10140 10668
rect 10192 10656 10198 10668
rect 12158 10656 12164 10668
rect 10192 10628 10285 10656
rect 12119 10628 12164 10656
rect 10192 10616 10198 10628
rect 12158 10616 12164 10628
rect 12216 10616 12222 10668
rect 12342 10656 12348 10668
rect 12303 10628 12348 10656
rect 12342 10616 12348 10628
rect 12400 10656 12406 10668
rect 12989 10659 13047 10665
rect 12989 10656 13001 10659
rect 12400 10628 13001 10656
rect 12400 10616 12406 10628
rect 12989 10625 13001 10628
rect 13035 10625 13047 10659
rect 13170 10656 13176 10668
rect 13131 10628 13176 10656
rect 12989 10619 13047 10625
rect 13170 10616 13176 10628
rect 13228 10616 13234 10668
rect 19291 10659 19349 10665
rect 19291 10656 19303 10659
rect 18616 10628 19303 10656
rect 3234 10588 3240 10600
rect 3195 10560 3240 10588
rect 3234 10548 3240 10560
rect 3292 10548 3298 10600
rect 4433 10591 4491 10597
rect 4433 10557 4445 10591
rect 4479 10588 4491 10591
rect 5994 10588 6000 10600
rect 4479 10560 6000 10588
rect 4479 10557 4491 10560
rect 4433 10551 4491 10557
rect 5994 10548 6000 10560
rect 6052 10588 6058 10600
rect 6733 10591 6791 10597
rect 6733 10588 6745 10591
rect 6052 10560 6745 10588
rect 6052 10548 6058 10560
rect 6733 10557 6745 10560
rect 6779 10557 6791 10591
rect 9490 10588 9496 10600
rect 9451 10560 9496 10588
rect 6733 10551 6791 10557
rect 9490 10548 9496 10560
rect 9548 10548 9554 10600
rect 10152 10588 10180 10616
rect 10686 10588 10692 10600
rect 10152 10560 10692 10588
rect 10686 10548 10692 10560
rect 10744 10548 10750 10600
rect 12176 10588 12204 10616
rect 12176 10560 13032 10588
rect 1581 10523 1639 10529
rect 1581 10489 1593 10523
rect 1627 10520 1639 10523
rect 6638 10520 6644 10532
rect 1627 10492 6644 10520
rect 1627 10489 1639 10492
rect 1581 10483 1639 10489
rect 6638 10480 6644 10492
rect 6696 10480 6702 10532
rect 11514 10412 11520 10464
rect 11572 10452 11578 10464
rect 11885 10455 11943 10461
rect 11885 10452 11897 10455
rect 11572 10424 11897 10452
rect 11572 10412 11578 10424
rect 11885 10421 11897 10424
rect 11931 10421 11943 10455
rect 11885 10415 11943 10421
rect 12434 10412 12440 10464
rect 12492 10452 12498 10464
rect 13004 10461 13032 10560
rect 12805 10455 12863 10461
rect 12805 10452 12817 10455
rect 12492 10424 12817 10452
rect 12492 10412 12498 10424
rect 12805 10421 12817 10424
rect 12851 10421 12863 10455
rect 12805 10415 12863 10421
rect 12989 10455 13047 10461
rect 12989 10421 13001 10455
rect 13035 10421 13047 10455
rect 12989 10415 13047 10421
rect 15746 10412 15752 10464
rect 15804 10452 15810 10464
rect 18616 10461 18644 10628
rect 19291 10625 19303 10628
rect 19337 10625 19349 10659
rect 19291 10619 19349 10625
rect 19521 10659 19579 10665
rect 19521 10625 19533 10659
rect 19567 10625 19579 10659
rect 19702 10656 19708 10668
rect 19663 10628 19708 10656
rect 19521 10619 19579 10625
rect 18601 10455 18659 10461
rect 18601 10452 18613 10455
rect 15804 10424 18613 10452
rect 15804 10412 15810 10424
rect 18601 10421 18613 10424
rect 18647 10421 18659 10455
rect 18601 10415 18659 10421
rect 18690 10412 18696 10464
rect 18748 10452 18754 10464
rect 19153 10455 19211 10461
rect 19153 10452 19165 10455
rect 18748 10424 19165 10452
rect 18748 10412 18754 10424
rect 19153 10421 19165 10424
rect 19199 10421 19211 10455
rect 19306 10452 19334 10619
rect 19536 10588 19564 10619
rect 19702 10616 19708 10628
rect 19760 10616 19766 10668
rect 19797 10659 19855 10665
rect 19797 10625 19809 10659
rect 19843 10656 19855 10659
rect 22922 10656 22928 10668
rect 19843 10628 22094 10656
rect 22835 10628 22928 10656
rect 19843 10625 19855 10628
rect 19797 10619 19855 10625
rect 20346 10588 20352 10600
rect 19536 10560 20352 10588
rect 20346 10548 20352 10560
rect 20404 10548 20410 10600
rect 22066 10520 22094 10628
rect 22922 10616 22928 10628
rect 22980 10616 22986 10668
rect 23290 10656 23296 10668
rect 23251 10628 23296 10656
rect 23290 10616 23296 10628
rect 23348 10616 23354 10668
rect 25133 10659 25191 10665
rect 25133 10625 25145 10659
rect 25179 10625 25191 10659
rect 25133 10619 25191 10625
rect 22940 10588 22968 10616
rect 23658 10588 23664 10600
rect 22940 10560 23664 10588
rect 23658 10548 23664 10560
rect 23716 10548 23722 10600
rect 25148 10588 25176 10619
rect 25222 10616 25228 10668
rect 25280 10656 25286 10668
rect 25501 10659 25559 10665
rect 25280 10628 25325 10656
rect 25280 10616 25286 10628
rect 25501 10625 25513 10659
rect 25547 10656 25559 10659
rect 25958 10656 25964 10668
rect 25547 10628 25964 10656
rect 25547 10625 25559 10628
rect 25501 10619 25559 10625
rect 25958 10616 25964 10628
rect 26016 10616 26022 10668
rect 27448 10665 27476 10752
rect 28966 10724 28994 10764
rect 29454 10752 29460 10804
rect 29512 10792 29518 10804
rect 42429 10795 42487 10801
rect 42429 10792 42441 10795
rect 29512 10764 29684 10792
rect 29512 10752 29518 10764
rect 29656 10733 29684 10764
rect 30024 10764 42441 10792
rect 29641 10727 29699 10733
rect 28966 10696 29500 10724
rect 27448 10659 27533 10665
rect 27448 10628 27487 10659
rect 27475 10625 27487 10628
rect 27521 10625 27533 10659
rect 27475 10619 27533 10625
rect 27893 10659 27951 10665
rect 27893 10625 27905 10659
rect 27939 10656 27951 10659
rect 28074 10656 28080 10668
rect 27939 10628 28080 10656
rect 27939 10625 27951 10628
rect 27893 10619 27951 10625
rect 28074 10616 28080 10628
rect 28132 10616 28138 10668
rect 29362 10656 29368 10668
rect 29323 10628 29368 10656
rect 29362 10616 29368 10628
rect 29420 10616 29426 10668
rect 29472 10665 29500 10696
rect 29641 10693 29653 10727
rect 29687 10693 29699 10727
rect 29641 10687 29699 10693
rect 29458 10659 29516 10665
rect 29458 10625 29470 10659
rect 29504 10625 29516 10659
rect 29730 10656 29736 10668
rect 29691 10628 29736 10656
rect 29458 10619 29516 10625
rect 29730 10616 29736 10628
rect 29788 10616 29794 10668
rect 29914 10665 29920 10668
rect 29871 10659 29920 10665
rect 29871 10625 29883 10659
rect 29917 10625 29920 10659
rect 29871 10619 29920 10625
rect 29914 10616 29920 10619
rect 29972 10616 29978 10668
rect 25406 10588 25412 10600
rect 25148 10560 25412 10588
rect 25406 10548 25412 10560
rect 25464 10548 25470 10600
rect 27341 10591 27399 10597
rect 27341 10557 27353 10591
rect 27387 10588 27399 10591
rect 27706 10588 27712 10600
rect 27387 10560 27712 10588
rect 27387 10557 27399 10560
rect 27341 10551 27399 10557
rect 27706 10548 27712 10560
rect 27764 10548 27770 10600
rect 28718 10548 28724 10600
rect 28776 10588 28782 10600
rect 30024 10588 30052 10764
rect 42429 10761 42441 10764
rect 42475 10792 42487 10795
rect 43162 10792 43168 10804
rect 42475 10764 43168 10792
rect 42475 10761 42487 10764
rect 42429 10755 42487 10761
rect 43162 10752 43168 10764
rect 43220 10752 43226 10804
rect 47670 10752 47676 10804
rect 47728 10792 47734 10804
rect 47949 10795 48007 10801
rect 47949 10792 47961 10795
rect 47728 10764 47961 10792
rect 47728 10752 47734 10764
rect 47949 10761 47961 10764
rect 47995 10761 48007 10795
rect 47949 10755 48007 10761
rect 52733 10795 52791 10801
rect 52733 10761 52745 10795
rect 52779 10792 52791 10795
rect 53006 10792 53012 10804
rect 52779 10764 53012 10792
rect 52779 10761 52791 10764
rect 52733 10755 52791 10761
rect 31478 10684 31484 10736
rect 31536 10724 31542 10736
rect 31536 10696 34100 10724
rect 31536 10684 31542 10696
rect 32677 10659 32735 10665
rect 32677 10656 32689 10659
rect 28776 10560 30052 10588
rect 31726 10628 32689 10656
rect 28776 10548 28782 10560
rect 22741 10523 22799 10529
rect 22741 10520 22753 10523
rect 22066 10492 22753 10520
rect 22741 10489 22753 10492
rect 22787 10489 22799 10523
rect 22741 10483 22799 10489
rect 23934 10480 23940 10532
rect 23992 10520 23998 10532
rect 27798 10520 27804 10532
rect 23992 10492 26188 10520
rect 27759 10492 27804 10520
rect 23992 10480 23998 10492
rect 24118 10452 24124 10464
rect 19306 10424 24124 10452
rect 19153 10415 19211 10421
rect 24118 10412 24124 10424
rect 24176 10412 24182 10464
rect 24302 10452 24308 10464
rect 24263 10424 24308 10452
rect 24302 10412 24308 10424
rect 24360 10412 24366 10464
rect 24946 10452 24952 10464
rect 24907 10424 24952 10452
rect 24946 10412 24952 10424
rect 25004 10412 25010 10464
rect 26050 10452 26056 10464
rect 26011 10424 26056 10452
rect 26050 10412 26056 10424
rect 26108 10412 26114 10464
rect 26160 10452 26188 10492
rect 27798 10480 27804 10492
rect 27856 10480 27862 10532
rect 30009 10523 30067 10529
rect 30009 10489 30021 10523
rect 30055 10520 30067 10523
rect 31726 10520 31754 10628
rect 32677 10625 32689 10628
rect 32723 10625 32735 10659
rect 33594 10656 33600 10668
rect 33555 10628 33600 10656
rect 32677 10619 32735 10625
rect 33594 10616 33600 10628
rect 33652 10616 33658 10668
rect 30055 10492 31754 10520
rect 34072 10520 34100 10696
rect 34698 10684 34704 10736
rect 34756 10724 34762 10736
rect 34885 10727 34943 10733
rect 34885 10724 34897 10727
rect 34756 10696 34897 10724
rect 34756 10684 34762 10696
rect 34885 10693 34897 10696
rect 34931 10693 34943 10727
rect 39669 10727 39727 10733
rect 39669 10724 39681 10727
rect 34885 10687 34943 10693
rect 36648 10696 37596 10724
rect 35161 10659 35219 10665
rect 35161 10625 35173 10659
rect 35207 10656 35219 10659
rect 35434 10656 35440 10668
rect 35207 10628 35440 10656
rect 35207 10625 35219 10628
rect 35161 10619 35219 10625
rect 35434 10616 35440 10628
rect 35492 10616 35498 10668
rect 36648 10665 36676 10696
rect 36633 10659 36691 10665
rect 36633 10625 36645 10659
rect 36679 10625 36691 10659
rect 37366 10656 37372 10668
rect 37327 10628 37372 10656
rect 36633 10619 36691 10625
rect 37366 10616 37372 10628
rect 37424 10616 37430 10668
rect 37568 10665 37596 10696
rect 38948 10696 39681 10724
rect 38948 10668 38976 10696
rect 39669 10693 39681 10696
rect 39715 10693 39727 10727
rect 39850 10724 39856 10736
rect 39811 10696 39856 10724
rect 39669 10687 39727 10693
rect 39850 10684 39856 10696
rect 39908 10684 39914 10736
rect 41138 10724 41144 10736
rect 39960 10696 41144 10724
rect 37553 10659 37611 10665
rect 37553 10625 37565 10659
rect 37599 10656 37611 10659
rect 38930 10656 38936 10668
rect 37599 10628 38792 10656
rect 38891 10628 38936 10656
rect 37599 10625 37611 10628
rect 37553 10619 37611 10625
rect 34790 10548 34796 10600
rect 34848 10588 34854 10600
rect 34977 10591 35035 10597
rect 34977 10588 34989 10591
rect 34848 10560 34989 10588
rect 34848 10548 34854 10560
rect 34977 10557 34989 10560
rect 35023 10557 35035 10591
rect 36357 10591 36415 10597
rect 36357 10588 36369 10591
rect 34977 10551 35035 10557
rect 35084 10560 36369 10588
rect 35084 10520 35112 10560
rect 36357 10557 36369 10560
rect 36403 10557 36415 10591
rect 38286 10588 38292 10600
rect 38247 10560 38292 10588
rect 36357 10551 36415 10557
rect 38286 10548 38292 10560
rect 38344 10548 38350 10600
rect 38764 10588 38792 10628
rect 38930 10616 38936 10628
rect 38988 10616 38994 10668
rect 39209 10659 39267 10665
rect 39209 10625 39221 10659
rect 39255 10656 39267 10659
rect 39868 10656 39896 10684
rect 39255 10628 39896 10656
rect 39255 10625 39267 10628
rect 39209 10619 39267 10625
rect 39960 10588 39988 10696
rect 40310 10616 40316 10668
rect 40368 10656 40374 10668
rect 40696 10665 40724 10696
rect 41138 10684 41144 10696
rect 41196 10684 41202 10736
rect 40681 10659 40739 10665
rect 40368 10628 40632 10656
rect 40368 10616 40374 10628
rect 40604 10597 40632 10628
rect 40681 10625 40693 10659
rect 40727 10625 40739 10659
rect 47964 10656 47992 10755
rect 53006 10752 53012 10764
rect 53064 10752 53070 10804
rect 53834 10752 53840 10804
rect 53892 10792 53898 10804
rect 54021 10795 54079 10801
rect 54021 10792 54033 10795
rect 53892 10764 54033 10792
rect 53892 10752 53898 10764
rect 54021 10761 54033 10764
rect 54067 10761 54079 10795
rect 54021 10755 54079 10761
rect 56226 10752 56232 10804
rect 56284 10792 56290 10804
rect 56321 10795 56379 10801
rect 56321 10792 56333 10795
rect 56284 10764 56333 10792
rect 56284 10752 56290 10764
rect 56321 10761 56333 10764
rect 56367 10761 56379 10795
rect 56321 10755 56379 10761
rect 51810 10684 51816 10736
rect 51868 10724 51874 10736
rect 53101 10727 53159 10733
rect 53101 10724 53113 10727
rect 51868 10696 53113 10724
rect 51868 10684 51874 10696
rect 53101 10693 53113 10696
rect 53147 10693 53159 10727
rect 55122 10724 55128 10736
rect 53101 10687 53159 10693
rect 53852 10696 55128 10724
rect 48593 10659 48651 10665
rect 48593 10656 48605 10659
rect 47964 10628 48605 10656
rect 40681 10619 40739 10625
rect 48593 10625 48605 10628
rect 48639 10625 48651 10659
rect 48958 10656 48964 10668
rect 48919 10628 48964 10656
rect 48593 10619 48651 10625
rect 48958 10616 48964 10628
rect 49016 10616 49022 10668
rect 51718 10656 51724 10668
rect 51679 10628 51724 10656
rect 51718 10616 51724 10628
rect 51776 10616 51782 10668
rect 52086 10656 52092 10668
rect 52047 10628 52092 10656
rect 52086 10616 52092 10628
rect 52144 10656 52150 10668
rect 52917 10659 52975 10665
rect 52917 10656 52929 10659
rect 52144 10628 52929 10656
rect 52144 10616 52150 10628
rect 52917 10625 52929 10628
rect 52963 10625 52975 10659
rect 52917 10619 52975 10625
rect 53193 10659 53251 10665
rect 53193 10625 53205 10659
rect 53239 10625 53251 10659
rect 53650 10656 53656 10668
rect 53611 10628 53656 10656
rect 53193 10619 53251 10625
rect 38764 10560 39988 10588
rect 40589 10591 40647 10597
rect 40589 10557 40601 10591
rect 40635 10557 40647 10591
rect 49510 10588 49516 10600
rect 49471 10560 49516 10588
rect 40589 10551 40647 10557
rect 49510 10548 49516 10560
rect 49568 10548 49574 10600
rect 51534 10548 51540 10600
rect 51592 10588 51598 10600
rect 51629 10591 51687 10597
rect 51629 10588 51641 10591
rect 51592 10560 51641 10588
rect 51592 10548 51598 10560
rect 51629 10557 51641 10560
rect 51675 10557 51687 10591
rect 53208 10588 53236 10619
rect 53650 10616 53656 10628
rect 53708 10616 53714 10668
rect 53852 10665 53880 10696
rect 55122 10684 55128 10696
rect 55180 10724 55186 10736
rect 55953 10727 56011 10733
rect 55953 10724 55965 10727
rect 55180 10696 55965 10724
rect 55180 10684 55186 10696
rect 55953 10693 55965 10696
rect 55999 10693 56011 10727
rect 55953 10687 56011 10693
rect 56137 10727 56195 10733
rect 56137 10693 56149 10727
rect 56183 10724 56195 10727
rect 56870 10724 56876 10736
rect 56183 10696 56876 10724
rect 56183 10693 56195 10696
rect 56137 10687 56195 10693
rect 56870 10684 56876 10696
rect 56928 10684 56934 10736
rect 53837 10659 53895 10665
rect 53837 10625 53849 10659
rect 53883 10625 53895 10659
rect 53837 10619 53895 10625
rect 54110 10616 54116 10668
rect 54168 10656 54174 10668
rect 54481 10659 54539 10665
rect 54481 10656 54493 10659
rect 54168 10628 54493 10656
rect 54168 10616 54174 10628
rect 54481 10625 54493 10628
rect 54527 10625 54539 10659
rect 54662 10656 54668 10668
rect 54623 10628 54668 10656
rect 54481 10619 54539 10625
rect 54662 10616 54668 10628
rect 54720 10616 54726 10668
rect 56778 10616 56784 10668
rect 56836 10656 56842 10668
rect 56965 10659 57023 10665
rect 56965 10656 56977 10659
rect 56836 10628 56977 10656
rect 56836 10616 56842 10628
rect 56965 10625 56977 10628
rect 57011 10625 57023 10659
rect 56965 10619 57023 10625
rect 57149 10659 57207 10665
rect 57149 10625 57161 10659
rect 57195 10656 57207 10659
rect 57422 10656 57428 10668
rect 57195 10628 57428 10656
rect 57195 10625 57207 10628
rect 57149 10619 57207 10625
rect 57422 10616 57428 10628
rect 57480 10616 57486 10668
rect 57606 10616 57612 10668
rect 57664 10656 57670 10668
rect 57885 10659 57943 10665
rect 57885 10656 57897 10659
rect 57664 10628 57897 10656
rect 57664 10616 57670 10628
rect 57885 10625 57897 10628
rect 57931 10625 57943 10659
rect 57885 10619 57943 10625
rect 54018 10588 54024 10600
rect 53208 10560 54024 10588
rect 51629 10551 51687 10557
rect 54018 10548 54024 10560
rect 54076 10548 54082 10600
rect 35250 10520 35256 10532
rect 34072 10492 35112 10520
rect 35176 10492 35256 10520
rect 30055 10489 30067 10492
rect 30009 10483 30067 10489
rect 29822 10452 29828 10464
rect 26160 10424 29828 10452
rect 29822 10412 29828 10424
rect 29880 10412 29886 10464
rect 30282 10412 30288 10464
rect 30340 10452 30346 10464
rect 30837 10455 30895 10461
rect 30837 10452 30849 10455
rect 30340 10424 30849 10452
rect 30340 10412 30346 10424
rect 30837 10421 30849 10424
rect 30883 10421 30895 10455
rect 30837 10415 30895 10421
rect 31018 10412 31024 10464
rect 31076 10452 31082 10464
rect 35176 10461 35204 10492
rect 35250 10480 35256 10492
rect 35308 10480 35314 10532
rect 38930 10520 38936 10532
rect 38891 10492 38936 10520
rect 38930 10480 38936 10492
rect 38988 10480 38994 10532
rect 32125 10455 32183 10461
rect 32125 10452 32137 10455
rect 31076 10424 32137 10452
rect 31076 10412 31082 10424
rect 32125 10421 32137 10424
rect 32171 10421 32183 10455
rect 32125 10415 32183 10421
rect 35161 10455 35219 10461
rect 35161 10421 35173 10455
rect 35207 10421 35219 10455
rect 35161 10415 35219 10421
rect 35345 10455 35403 10461
rect 35345 10421 35357 10455
rect 35391 10452 35403 10455
rect 35526 10452 35532 10464
rect 35391 10424 35532 10452
rect 35391 10421 35403 10424
rect 35345 10415 35403 10421
rect 35526 10412 35532 10424
rect 35584 10412 35590 10464
rect 39850 10412 39856 10464
rect 39908 10452 39914 10464
rect 39945 10455 40003 10461
rect 39945 10452 39957 10455
rect 39908 10424 39957 10452
rect 39908 10412 39914 10424
rect 39945 10421 39957 10424
rect 39991 10421 40003 10455
rect 40954 10452 40960 10464
rect 40915 10424 40960 10452
rect 39945 10415 40003 10421
rect 40954 10412 40960 10424
rect 41012 10412 41018 10464
rect 54570 10452 54576 10464
rect 54531 10424 54576 10452
rect 54570 10412 54576 10424
rect 54628 10412 54634 10464
rect 56502 10412 56508 10464
rect 56560 10452 56566 10464
rect 56781 10455 56839 10461
rect 56781 10452 56793 10455
rect 56560 10424 56793 10452
rect 56560 10412 56566 10424
rect 56781 10421 56793 10424
rect 56827 10421 56839 10455
rect 58066 10452 58072 10464
rect 58027 10424 58072 10452
rect 56781 10415 56839 10421
rect 58066 10412 58072 10424
rect 58124 10412 58130 10464
rect 1104 10362 58880 10384
rect 1104 10310 4214 10362
rect 4266 10310 4278 10362
rect 4330 10310 4342 10362
rect 4394 10310 4406 10362
rect 4458 10310 4470 10362
rect 4522 10310 34934 10362
rect 34986 10310 34998 10362
rect 35050 10310 35062 10362
rect 35114 10310 35126 10362
rect 35178 10310 35190 10362
rect 35242 10310 58880 10362
rect 1104 10288 58880 10310
rect 1394 10248 1400 10260
rect 1355 10220 1400 10248
rect 1394 10208 1400 10220
rect 1452 10208 1458 10260
rect 5813 10251 5871 10257
rect 5813 10217 5825 10251
rect 5859 10248 5871 10251
rect 5994 10248 6000 10260
rect 5859 10220 6000 10248
rect 5859 10217 5871 10220
rect 5813 10211 5871 10217
rect 5828 10180 5856 10211
rect 5994 10208 6000 10220
rect 6052 10208 6058 10260
rect 6641 10251 6699 10257
rect 6641 10217 6653 10251
rect 6687 10217 6699 10251
rect 6822 10248 6828 10260
rect 6783 10220 6828 10248
rect 6641 10211 6699 10217
rect 3988 10152 5856 10180
rect 5905 10183 5963 10189
rect 2866 10004 2872 10056
rect 2924 10044 2930 10056
rect 2961 10047 3019 10053
rect 2961 10044 2973 10047
rect 2924 10016 2973 10044
rect 2924 10004 2930 10016
rect 2961 10013 2973 10016
rect 3007 10013 3019 10047
rect 3142 10044 3148 10056
rect 3103 10016 3148 10044
rect 2961 10007 3019 10013
rect 3142 10004 3148 10016
rect 3200 10004 3206 10056
rect 3988 10053 4016 10152
rect 5905 10149 5917 10183
rect 5951 10180 5963 10183
rect 6656 10180 6684 10211
rect 6822 10208 6828 10220
rect 6880 10208 6886 10260
rect 9401 10251 9459 10257
rect 9401 10217 9413 10251
rect 9447 10248 9459 10251
rect 9490 10248 9496 10260
rect 9447 10220 9496 10248
rect 9447 10217 9459 10220
rect 9401 10211 9459 10217
rect 9490 10208 9496 10220
rect 9548 10208 9554 10260
rect 12158 10208 12164 10260
rect 12216 10248 12222 10260
rect 12253 10251 12311 10257
rect 12253 10248 12265 10251
rect 12216 10220 12265 10248
rect 12216 10208 12222 10220
rect 12253 10217 12265 10220
rect 12299 10217 12311 10251
rect 12253 10211 12311 10217
rect 21818 10208 21824 10260
rect 21876 10248 21882 10260
rect 22462 10248 22468 10260
rect 21876 10220 22468 10248
rect 21876 10208 21882 10220
rect 22462 10208 22468 10220
rect 22520 10248 22526 10260
rect 25314 10248 25320 10260
rect 22520 10220 25320 10248
rect 22520 10208 22526 10220
rect 25314 10208 25320 10220
rect 25372 10208 25378 10260
rect 31570 10208 31576 10260
rect 31628 10248 31634 10260
rect 36354 10248 36360 10260
rect 31628 10220 32168 10248
rect 36315 10220 36360 10248
rect 31628 10208 31634 10220
rect 6914 10180 6920 10192
rect 5951 10152 6920 10180
rect 5951 10149 5963 10152
rect 5905 10143 5963 10149
rect 6914 10140 6920 10152
rect 6972 10140 6978 10192
rect 19150 10140 19156 10192
rect 19208 10180 19214 10192
rect 19245 10183 19303 10189
rect 19245 10180 19257 10183
rect 19208 10152 19257 10180
rect 19208 10140 19214 10152
rect 19245 10149 19257 10152
rect 19291 10149 19303 10183
rect 19245 10143 19303 10149
rect 20346 10140 20352 10192
rect 20404 10180 20410 10192
rect 20901 10183 20959 10189
rect 20901 10180 20913 10183
rect 20404 10152 20913 10180
rect 20404 10140 20410 10152
rect 20901 10149 20913 10152
rect 20947 10180 20959 10183
rect 27430 10180 27436 10192
rect 20947 10152 27436 10180
rect 20947 10149 20959 10152
rect 20901 10143 20959 10149
rect 27430 10140 27436 10152
rect 27488 10140 27494 10192
rect 29730 10140 29736 10192
rect 29788 10180 29794 10192
rect 29917 10183 29975 10189
rect 29917 10180 29929 10183
rect 29788 10152 29929 10180
rect 29788 10140 29794 10152
rect 29917 10149 29929 10152
rect 29963 10149 29975 10183
rect 29917 10143 29975 10149
rect 5721 10115 5779 10121
rect 5721 10081 5733 10115
rect 5767 10112 5779 10115
rect 6362 10112 6368 10124
rect 5767 10084 6368 10112
rect 5767 10081 5779 10084
rect 5721 10075 5779 10081
rect 6362 10072 6368 10084
rect 6420 10112 6426 10124
rect 6420 10084 6500 10112
rect 6420 10072 6426 10084
rect 6472 10053 6500 10084
rect 8846 10072 8852 10124
rect 8904 10112 8910 10124
rect 9033 10115 9091 10121
rect 9033 10112 9045 10115
rect 8904 10084 9045 10112
rect 8904 10072 8910 10084
rect 9033 10081 9045 10084
rect 9079 10081 9091 10115
rect 12618 10112 12624 10124
rect 12579 10084 12624 10112
rect 9033 10075 9091 10081
rect 12618 10072 12624 10084
rect 12676 10072 12682 10124
rect 15013 10115 15071 10121
rect 15013 10081 15025 10115
rect 15059 10112 15071 10115
rect 18690 10112 18696 10124
rect 15059 10084 18696 10112
rect 15059 10081 15071 10084
rect 15013 10075 15071 10081
rect 18690 10072 18696 10084
rect 18748 10072 18754 10124
rect 21729 10115 21787 10121
rect 21729 10081 21741 10115
rect 21775 10112 21787 10115
rect 26237 10115 26295 10121
rect 21775 10084 22876 10112
rect 21775 10081 21787 10084
rect 21729 10075 21787 10081
rect 3789 10047 3847 10053
rect 3789 10013 3801 10047
rect 3835 10013 3847 10047
rect 3789 10007 3847 10013
rect 3973 10047 4031 10053
rect 3973 10013 3985 10047
rect 4019 10013 4031 10047
rect 3973 10007 4031 10013
rect 5997 10047 6055 10053
rect 5997 10013 6009 10047
rect 6043 10013 6055 10047
rect 5997 10007 6055 10013
rect 6457 10047 6515 10053
rect 6457 10013 6469 10047
rect 6503 10013 6515 10047
rect 6457 10007 6515 10013
rect 6641 10047 6699 10053
rect 6641 10013 6653 10047
rect 6687 10044 6699 10047
rect 8202 10044 8208 10056
rect 6687 10016 8208 10044
rect 6687 10013 6699 10016
rect 6641 10007 6699 10013
rect 3804 9976 3832 10007
rect 4062 9976 4068 9988
rect 3804 9948 4068 9976
rect 4062 9936 4068 9948
rect 4120 9936 4126 9988
rect 6012 9976 6040 10007
rect 6656 9976 6684 10007
rect 8202 10004 8208 10016
rect 8260 10004 8266 10056
rect 9125 10047 9183 10053
rect 9125 10013 9137 10047
rect 9171 10044 9183 10047
rect 12437 10047 12495 10053
rect 9171 10016 9628 10044
rect 9171 10013 9183 10016
rect 9125 10007 9183 10013
rect 6012 9948 6684 9976
rect 9600 9920 9628 10016
rect 12437 10013 12449 10047
rect 12483 10044 12495 10047
rect 14918 10044 14924 10056
rect 12483 10016 13124 10044
rect 14879 10016 14924 10044
rect 12483 10013 12495 10016
rect 12437 10007 12495 10013
rect 13096 9920 13124 10016
rect 14918 10004 14924 10016
rect 14976 10004 14982 10056
rect 15102 10004 15108 10056
rect 15160 10044 15166 10056
rect 15657 10047 15715 10053
rect 15657 10044 15669 10047
rect 15160 10016 15669 10044
rect 15160 10004 15166 10016
rect 15657 10013 15669 10016
rect 15703 10013 15715 10047
rect 15657 10007 15715 10013
rect 15933 10047 15991 10053
rect 15933 10013 15945 10047
rect 15979 10044 15991 10047
rect 16577 10047 16635 10053
rect 16577 10044 16589 10047
rect 15979 10016 16589 10044
rect 15979 10013 15991 10016
rect 15933 10007 15991 10013
rect 16577 10013 16589 10016
rect 16623 10013 16635 10047
rect 16577 10007 16635 10013
rect 16761 10047 16819 10053
rect 16761 10013 16773 10047
rect 16807 10044 16819 10047
rect 16942 10044 16948 10056
rect 16807 10016 16948 10044
rect 16807 10013 16819 10016
rect 16761 10007 16819 10013
rect 16942 10004 16948 10016
rect 17000 10004 17006 10056
rect 17034 10004 17040 10056
rect 17092 10044 17098 10056
rect 19242 10044 19248 10056
rect 17092 10016 17137 10044
rect 19203 10016 19248 10044
rect 17092 10004 17098 10016
rect 19242 10004 19248 10016
rect 19300 10004 19306 10056
rect 19429 10047 19487 10053
rect 19429 10013 19441 10047
rect 19475 10044 19487 10047
rect 20254 10044 20260 10056
rect 19475 10016 20260 10044
rect 19475 10013 19487 10016
rect 19429 10007 19487 10013
rect 20254 10004 20260 10016
rect 20312 10044 20318 10056
rect 20438 10044 20444 10056
rect 20312 10016 20444 10044
rect 20312 10004 20318 10016
rect 20438 10004 20444 10016
rect 20496 10044 20502 10056
rect 21637 10047 21695 10053
rect 21637 10044 21649 10047
rect 20496 10016 21649 10044
rect 20496 10004 20502 10016
rect 21637 10013 21649 10016
rect 21683 10013 21695 10047
rect 21818 10044 21824 10056
rect 21779 10016 21824 10044
rect 21637 10007 21695 10013
rect 21818 10004 21824 10016
rect 21876 10004 21882 10056
rect 22848 10053 22876 10084
rect 26237 10081 26249 10115
rect 26283 10112 26295 10115
rect 27522 10112 27528 10124
rect 26283 10084 27528 10112
rect 26283 10081 26295 10084
rect 26237 10075 26295 10081
rect 27522 10072 27528 10084
rect 27580 10072 27586 10124
rect 27614 10072 27620 10124
rect 27672 10112 27678 10124
rect 28169 10115 28227 10121
rect 28169 10112 28181 10115
rect 27672 10084 28181 10112
rect 27672 10072 27678 10084
rect 28169 10081 28181 10084
rect 28215 10081 28227 10115
rect 28169 10075 28227 10081
rect 29362 10072 29368 10124
rect 29420 10112 29426 10124
rect 29420 10084 31754 10112
rect 29420 10072 29426 10084
rect 22557 10047 22615 10053
rect 22557 10013 22569 10047
rect 22603 10013 22615 10047
rect 22557 10007 22615 10013
rect 22649 10047 22707 10053
rect 22649 10013 22661 10047
rect 22695 10044 22707 10047
rect 22833 10047 22891 10053
rect 22695 10016 22784 10044
rect 22695 10013 22707 10016
rect 22649 10007 22707 10013
rect 21085 9979 21143 9985
rect 21085 9945 21097 9979
rect 21131 9976 21143 9979
rect 22572 9976 22600 10007
rect 22756 9976 22784 10016
rect 22833 10013 22845 10047
rect 22879 10013 22891 10047
rect 22833 10007 22891 10013
rect 22925 10047 22983 10053
rect 22925 10013 22937 10047
rect 22971 10044 22983 10047
rect 24946 10044 24952 10056
rect 22971 10016 24952 10044
rect 22971 10013 22983 10016
rect 22925 10007 22983 10013
rect 24946 10004 24952 10016
rect 25004 10004 25010 10056
rect 26510 10044 26516 10056
rect 26471 10016 26516 10044
rect 26510 10004 26516 10016
rect 26568 10004 26574 10056
rect 28442 10044 28448 10056
rect 28403 10016 28448 10044
rect 28442 10004 28448 10016
rect 28500 10004 28506 10056
rect 30101 10047 30159 10053
rect 30101 10013 30113 10047
rect 30147 10044 30159 10047
rect 30742 10044 30748 10056
rect 30147 10016 30748 10044
rect 30147 10013 30159 10016
rect 30101 10007 30159 10013
rect 23382 9976 23388 9988
rect 21131 9948 22692 9976
rect 22756 9948 23388 9976
rect 21131 9945 21143 9948
rect 21085 9939 21143 9945
rect 22664 9920 22692 9948
rect 23382 9936 23388 9948
rect 23440 9936 23446 9988
rect 23658 9936 23664 9988
rect 23716 9976 23722 9988
rect 25498 9976 25504 9988
rect 23716 9948 25504 9976
rect 23716 9936 23722 9948
rect 25498 9936 25504 9948
rect 25556 9936 25562 9988
rect 25590 9936 25596 9988
rect 25648 9976 25654 9988
rect 25958 9976 25964 9988
rect 25648 9948 25964 9976
rect 25648 9936 25654 9948
rect 25958 9936 25964 9948
rect 26016 9976 26022 9988
rect 30116 9976 30144 10007
rect 30742 10004 30748 10016
rect 30800 10004 30806 10056
rect 26016 9948 30144 9976
rect 26016 9936 26022 9948
rect 3053 9911 3111 9917
rect 3053 9877 3065 9911
rect 3099 9908 3111 9911
rect 3418 9908 3424 9920
rect 3099 9880 3424 9908
rect 3099 9877 3111 9880
rect 3053 9871 3111 9877
rect 3418 9868 3424 9880
rect 3476 9868 3482 9920
rect 3786 9868 3792 9920
rect 3844 9908 3850 9920
rect 3881 9911 3939 9917
rect 3881 9908 3893 9911
rect 3844 9880 3893 9908
rect 3844 9868 3850 9880
rect 3881 9877 3893 9880
rect 3927 9877 3939 9911
rect 3881 9871 3939 9877
rect 9582 9868 9588 9920
rect 9640 9908 9646 9920
rect 9953 9911 10011 9917
rect 9953 9908 9965 9911
rect 9640 9880 9965 9908
rect 9640 9868 9646 9880
rect 9953 9877 9965 9880
rect 9999 9877 10011 9911
rect 9953 9871 10011 9877
rect 13078 9868 13084 9920
rect 13136 9908 13142 9920
rect 14093 9911 14151 9917
rect 14093 9908 14105 9911
rect 13136 9880 14105 9908
rect 13136 9868 13142 9880
rect 14093 9877 14105 9880
rect 14139 9877 14151 9911
rect 15746 9908 15752 9920
rect 15707 9880 15752 9908
rect 14093 9871 14151 9877
rect 15746 9868 15752 9880
rect 15804 9868 15810 9920
rect 16117 9911 16175 9917
rect 16117 9877 16129 9911
rect 16163 9908 16175 9911
rect 16574 9908 16580 9920
rect 16163 9880 16580 9908
rect 16163 9877 16175 9880
rect 16117 9871 16175 9877
rect 16574 9868 16580 9880
rect 16632 9868 16638 9920
rect 16850 9868 16856 9920
rect 16908 9908 16914 9920
rect 16945 9911 17003 9917
rect 16945 9908 16957 9911
rect 16908 9880 16957 9908
rect 16908 9868 16914 9880
rect 16945 9877 16957 9880
rect 16991 9877 17003 9911
rect 22370 9908 22376 9920
rect 22331 9880 22376 9908
rect 16945 9871 17003 9877
rect 22370 9868 22376 9880
rect 22428 9868 22434 9920
rect 22646 9868 22652 9920
rect 22704 9868 22710 9920
rect 24581 9911 24639 9917
rect 24581 9877 24593 9911
rect 24627 9908 24639 9911
rect 24762 9908 24768 9920
rect 24627 9880 24768 9908
rect 24627 9877 24639 9880
rect 24581 9871 24639 9877
rect 24762 9868 24768 9880
rect 24820 9868 24826 9920
rect 27706 9868 27712 9920
rect 27764 9908 27770 9920
rect 30834 9908 30840 9920
rect 27764 9880 30840 9908
rect 27764 9868 27770 9880
rect 30834 9868 30840 9880
rect 30892 9868 30898 9920
rect 31726 9908 31754 10084
rect 32140 9985 32168 10220
rect 36354 10208 36360 10220
rect 36412 10208 36418 10260
rect 38749 10251 38807 10257
rect 38749 10217 38761 10251
rect 38795 10248 38807 10251
rect 39298 10248 39304 10260
rect 38795 10220 39304 10248
rect 38795 10217 38807 10220
rect 38749 10211 38807 10217
rect 38764 10180 38792 10211
rect 39298 10208 39304 10220
rect 39356 10248 39362 10260
rect 39853 10251 39911 10257
rect 39853 10248 39865 10251
rect 39356 10220 39865 10248
rect 39356 10208 39362 10220
rect 39853 10217 39865 10220
rect 39899 10217 39911 10251
rect 39853 10211 39911 10217
rect 41046 10208 41052 10260
rect 41104 10248 41110 10260
rect 41104 10220 42196 10248
rect 41104 10208 41110 10220
rect 33520 10152 38792 10180
rect 38933 10183 38991 10189
rect 32674 10044 32680 10056
rect 32635 10016 32680 10044
rect 32674 10004 32680 10016
rect 32732 10004 32738 10056
rect 33045 10047 33103 10053
rect 33045 10013 33057 10047
rect 33091 10044 33103 10047
rect 33410 10044 33416 10056
rect 33091 10016 33416 10044
rect 33091 10013 33103 10016
rect 33045 10007 33103 10013
rect 32125 9979 32183 9985
rect 32125 9945 32137 9979
rect 32171 9976 32183 9979
rect 33060 9976 33088 10007
rect 33410 10004 33416 10016
rect 33468 10004 33474 10056
rect 32171 9948 33088 9976
rect 32171 9945 32183 9948
rect 32125 9939 32183 9945
rect 33520 9908 33548 10152
rect 38933 10149 38945 10183
rect 38979 10180 38991 10183
rect 41874 10180 41880 10192
rect 38979 10152 41880 10180
rect 38979 10149 38991 10152
rect 38933 10143 38991 10149
rect 41874 10140 41880 10152
rect 41932 10140 41938 10192
rect 40972 10084 41920 10112
rect 40972 10056 41000 10084
rect 36173 10047 36231 10053
rect 36173 10044 36185 10047
rect 35636 10016 36185 10044
rect 33686 9908 33692 9920
rect 31726 9880 33548 9908
rect 33647 9880 33692 9908
rect 33686 9868 33692 9880
rect 33744 9868 33750 9920
rect 35342 9868 35348 9920
rect 35400 9908 35406 9920
rect 35636 9917 35664 10016
rect 36173 10013 36185 10016
rect 36219 10013 36231 10047
rect 36538 10044 36544 10056
rect 36499 10016 36544 10044
rect 36173 10007 36231 10013
rect 36538 10004 36544 10016
rect 36596 10004 36602 10056
rect 40954 10044 40960 10056
rect 40915 10016 40960 10044
rect 40954 10004 40960 10016
rect 41012 10004 41018 10056
rect 41046 10004 41052 10056
rect 41104 10044 41110 10056
rect 41141 10047 41199 10053
rect 41141 10044 41153 10047
rect 41104 10016 41153 10044
rect 41104 10004 41110 10016
rect 41141 10013 41153 10016
rect 41187 10013 41199 10047
rect 41141 10007 41199 10013
rect 41233 10047 41291 10053
rect 41233 10013 41245 10047
rect 41279 10044 41291 10047
rect 41414 10044 41420 10056
rect 41279 10016 41420 10044
rect 41279 10013 41291 10016
rect 41233 10007 41291 10013
rect 41414 10004 41420 10016
rect 41472 10044 41478 10056
rect 41782 10044 41788 10056
rect 41472 10016 41788 10044
rect 41472 10004 41478 10016
rect 41782 10004 41788 10016
rect 41840 10004 41846 10056
rect 41892 10053 41920 10084
rect 42168 10053 42196 10220
rect 51718 10208 51724 10260
rect 51776 10248 51782 10260
rect 53469 10251 53527 10257
rect 53469 10248 53481 10251
rect 51776 10220 53481 10248
rect 51776 10208 51782 10220
rect 53469 10217 53481 10220
rect 53515 10248 53527 10251
rect 53650 10248 53656 10260
rect 53515 10220 53656 10248
rect 53515 10217 53527 10220
rect 53469 10211 53527 10217
rect 53650 10208 53656 10220
rect 53708 10208 53714 10260
rect 55677 10251 55735 10257
rect 55677 10217 55689 10251
rect 55723 10248 55735 10251
rect 56686 10248 56692 10260
rect 55723 10220 56692 10248
rect 55723 10217 55735 10220
rect 55677 10211 55735 10217
rect 56686 10208 56692 10220
rect 56744 10208 56750 10260
rect 43162 10112 43168 10124
rect 43123 10084 43168 10112
rect 43162 10072 43168 10084
rect 43220 10072 43226 10124
rect 45554 10112 45560 10124
rect 45515 10084 45560 10112
rect 45554 10072 45560 10084
rect 45612 10072 45618 10124
rect 46017 10115 46075 10121
rect 46017 10081 46029 10115
rect 46063 10112 46075 10115
rect 48501 10115 48559 10121
rect 48501 10112 48513 10115
rect 46063 10084 48513 10112
rect 46063 10081 46075 10084
rect 46017 10075 46075 10081
rect 48501 10081 48513 10084
rect 48547 10112 48559 10115
rect 49237 10115 49295 10121
rect 48547 10084 49188 10112
rect 48547 10081 48559 10084
rect 48501 10075 48559 10081
rect 41877 10047 41935 10053
rect 41877 10013 41889 10047
rect 41923 10013 41935 10047
rect 41877 10007 41935 10013
rect 42153 10047 42211 10053
rect 42153 10013 42165 10047
rect 42199 10013 42211 10047
rect 42153 10007 42211 10013
rect 42613 10047 42671 10053
rect 42613 10013 42625 10047
rect 42659 10013 42671 10047
rect 42613 10007 42671 10013
rect 42797 10047 42855 10053
rect 42797 10013 42809 10047
rect 42843 10044 42855 10047
rect 45649 10047 45707 10053
rect 45649 10044 45661 10047
rect 42843 10016 43024 10044
rect 42843 10013 42855 10016
rect 42797 10007 42855 10013
rect 38470 9936 38476 9988
rect 38528 9976 38534 9988
rect 38565 9979 38623 9985
rect 38565 9976 38577 9979
rect 38528 9948 38577 9976
rect 38528 9936 38534 9948
rect 38565 9945 38577 9948
rect 38611 9945 38623 9979
rect 38565 9939 38623 9945
rect 38654 9936 38660 9988
rect 38712 9976 38718 9988
rect 38765 9979 38823 9985
rect 38765 9976 38777 9979
rect 38712 9948 38777 9976
rect 38712 9936 38718 9948
rect 38765 9945 38777 9948
rect 38811 9945 38823 9979
rect 42628 9976 42656 10007
rect 42886 9976 42892 9988
rect 38765 9939 38823 9945
rect 41524 9948 42892 9976
rect 41524 9920 41552 9948
rect 42886 9936 42892 9948
rect 42944 9936 42950 9988
rect 35621 9911 35679 9917
rect 35621 9908 35633 9911
rect 35400 9880 35633 9908
rect 35400 9868 35406 9880
rect 35621 9877 35633 9880
rect 35667 9877 35679 9911
rect 36722 9908 36728 9920
rect 36683 9880 36728 9908
rect 35621 9871 35679 9877
rect 36722 9868 36728 9880
rect 36780 9868 36786 9920
rect 41233 9911 41291 9917
rect 41233 9877 41245 9911
rect 41279 9908 41291 9911
rect 41506 9908 41512 9920
rect 41279 9880 41512 9908
rect 41279 9877 41291 9880
rect 41233 9871 41291 9877
rect 41506 9868 41512 9880
rect 41564 9868 41570 9920
rect 41690 9908 41696 9920
rect 41651 9880 41696 9908
rect 41690 9868 41696 9880
rect 41748 9868 41754 9920
rect 41782 9868 41788 9920
rect 41840 9908 41846 9920
rect 42061 9911 42119 9917
rect 42061 9908 42073 9911
rect 41840 9880 42073 9908
rect 41840 9868 41846 9880
rect 42061 9877 42073 9880
rect 42107 9908 42119 9911
rect 42702 9908 42708 9920
rect 42107 9880 42708 9908
rect 42107 9877 42119 9880
rect 42061 9871 42119 9877
rect 42702 9868 42708 9880
rect 42760 9908 42766 9920
rect 42996 9908 43024 10016
rect 44192 10016 45661 10044
rect 44192 9920 44220 10016
rect 45649 10013 45661 10016
rect 45695 10013 45707 10047
rect 47762 10044 47768 10056
rect 47723 10016 47768 10044
rect 45649 10007 45707 10013
rect 47762 10004 47768 10016
rect 47820 10004 47826 10056
rect 48133 10047 48191 10053
rect 48133 10013 48145 10047
rect 48179 10044 48191 10047
rect 48406 10044 48412 10056
rect 48179 10016 48412 10044
rect 48179 10013 48191 10016
rect 48133 10007 48191 10013
rect 48406 10004 48412 10016
rect 48464 10004 48470 10056
rect 49160 10053 49188 10084
rect 49237 10081 49249 10115
rect 49283 10081 49295 10115
rect 49237 10075 49295 10081
rect 49513 10115 49571 10121
rect 49513 10081 49525 10115
rect 49559 10112 49571 10115
rect 55582 10112 55588 10124
rect 49559 10084 51074 10112
rect 55543 10084 55588 10112
rect 49559 10081 49571 10084
rect 49513 10075 49571 10081
rect 49145 10047 49203 10053
rect 49145 10013 49157 10047
rect 49191 10013 49203 10047
rect 49145 10007 49203 10013
rect 48424 9976 48452 10004
rect 49252 9976 49280 10075
rect 51046 10044 51074 10084
rect 55582 10072 55588 10084
rect 55640 10072 55646 10124
rect 55769 10115 55827 10121
rect 55769 10081 55781 10115
rect 55815 10112 55827 10115
rect 56502 10112 56508 10124
rect 55815 10084 56508 10112
rect 55815 10081 55827 10084
rect 55769 10075 55827 10081
rect 56502 10072 56508 10084
rect 56560 10112 56566 10124
rect 56560 10084 56824 10112
rect 56560 10072 56566 10084
rect 51537 10047 51595 10053
rect 51046 10016 51488 10044
rect 51166 9976 51172 9988
rect 48424 9948 49280 9976
rect 51127 9948 51172 9976
rect 51166 9936 51172 9948
rect 51224 9936 51230 9988
rect 51460 9976 51488 10016
rect 51537 10013 51549 10047
rect 51583 10044 51595 10047
rect 51810 10044 51816 10056
rect 51583 10016 51816 10044
rect 51583 10013 51595 10016
rect 51537 10007 51595 10013
rect 51810 10004 51816 10016
rect 51868 10004 51874 10056
rect 55861 10047 55919 10053
rect 55861 10013 55873 10047
rect 55907 10044 55919 10047
rect 55950 10044 55956 10056
rect 55907 10016 55956 10044
rect 55907 10013 55919 10016
rect 55861 10007 55919 10013
rect 55950 10004 55956 10016
rect 56008 10004 56014 10056
rect 56796 10053 56824 10084
rect 56781 10047 56839 10053
rect 56781 10013 56793 10047
rect 56827 10013 56839 10047
rect 56962 10044 56968 10056
rect 56923 10016 56968 10044
rect 56781 10007 56839 10013
rect 56962 10004 56968 10016
rect 57020 10004 57026 10056
rect 51721 9979 51779 9985
rect 51721 9976 51733 9979
rect 51460 9948 51733 9976
rect 51721 9945 51733 9948
rect 51767 9976 51779 9979
rect 52086 9976 52092 9988
rect 51767 9948 52092 9976
rect 51767 9945 51779 9948
rect 51721 9939 51779 9945
rect 52086 9936 52092 9948
rect 52144 9936 52150 9988
rect 42760 9880 43024 9908
rect 43073 9911 43131 9917
rect 42760 9868 42766 9880
rect 43073 9877 43085 9911
rect 43119 9908 43131 9911
rect 44174 9908 44180 9920
rect 43119 9880 44180 9908
rect 43119 9877 43131 9880
rect 43073 9871 43131 9877
rect 44174 9868 44180 9880
rect 44232 9868 44238 9920
rect 57146 9908 57152 9920
rect 57107 9880 57152 9908
rect 57146 9868 57152 9880
rect 57204 9868 57210 9920
rect 57606 9868 57612 9920
rect 57664 9908 57670 9920
rect 57701 9911 57759 9917
rect 57701 9908 57713 9911
rect 57664 9880 57713 9908
rect 57664 9868 57670 9880
rect 57701 9877 57713 9880
rect 57747 9877 57759 9911
rect 57701 9871 57759 9877
rect 1104 9818 58880 9840
rect 1104 9766 19574 9818
rect 19626 9766 19638 9818
rect 19690 9766 19702 9818
rect 19754 9766 19766 9818
rect 19818 9766 19830 9818
rect 19882 9766 50294 9818
rect 50346 9766 50358 9818
rect 50410 9766 50422 9818
rect 50474 9766 50486 9818
rect 50538 9766 50550 9818
rect 50602 9766 58880 9818
rect 1104 9744 58880 9766
rect 6362 9704 6368 9716
rect 6323 9676 6368 9704
rect 6362 9664 6368 9676
rect 6420 9664 6426 9716
rect 13998 9664 14004 9716
rect 14056 9704 14062 9716
rect 15289 9707 15347 9713
rect 15289 9704 15301 9707
rect 14056 9676 15301 9704
rect 14056 9664 14062 9676
rect 15289 9673 15301 9676
rect 15335 9704 15347 9707
rect 15746 9704 15752 9716
rect 15335 9676 15752 9704
rect 15335 9673 15347 9676
rect 15289 9667 15347 9673
rect 15746 9664 15752 9676
rect 15804 9664 15810 9716
rect 23290 9704 23296 9716
rect 18800 9676 20668 9704
rect 13728 9648 13780 9654
rect 6914 9596 6920 9648
rect 6972 9636 6978 9648
rect 8665 9639 8723 9645
rect 8665 9636 8677 9639
rect 6972 9608 8677 9636
rect 6972 9596 6978 9608
rect 8665 9605 8677 9608
rect 8711 9605 8723 9639
rect 9582 9636 9588 9648
rect 8665 9599 8723 9605
rect 9048 9608 9588 9636
rect 3050 9528 3056 9580
rect 3108 9568 3114 9580
rect 3145 9571 3203 9577
rect 3145 9568 3157 9571
rect 3108 9540 3157 9568
rect 3108 9528 3114 9540
rect 3145 9537 3157 9540
rect 3191 9537 3203 9571
rect 3418 9568 3424 9580
rect 3379 9540 3424 9568
rect 3145 9531 3203 9537
rect 3418 9528 3424 9540
rect 3476 9528 3482 9580
rect 3697 9571 3755 9577
rect 3697 9537 3709 9571
rect 3743 9537 3755 9571
rect 3697 9531 3755 9537
rect 3712 9500 3740 9531
rect 3786 9528 3792 9580
rect 3844 9568 3850 9580
rect 4065 9571 4123 9577
rect 3844 9540 3889 9568
rect 3844 9528 3850 9540
rect 4065 9537 4077 9571
rect 4111 9568 4123 9571
rect 4614 9568 4620 9580
rect 4111 9540 4620 9568
rect 4111 9537 4123 9540
rect 4065 9531 4123 9537
rect 4614 9528 4620 9540
rect 4672 9528 4678 9580
rect 6733 9571 6791 9577
rect 6733 9537 6745 9571
rect 6779 9537 6791 9571
rect 8846 9568 8852 9580
rect 8807 9540 8852 9568
rect 6733 9531 6791 9537
rect 3068 9472 3740 9500
rect 3068 9444 3096 9472
rect 6546 9460 6552 9512
rect 6604 9500 6610 9512
rect 6641 9503 6699 9509
rect 6641 9500 6653 9503
rect 6604 9472 6653 9500
rect 6604 9460 6610 9472
rect 6641 9469 6653 9472
rect 6687 9469 6699 9503
rect 6748 9500 6776 9531
rect 8846 9528 8852 9540
rect 8904 9528 8910 9580
rect 9048 9577 9076 9608
rect 9582 9596 9588 9608
rect 9640 9596 9646 9648
rect 17034 9596 17040 9648
rect 17092 9636 17098 9648
rect 17957 9639 18015 9645
rect 17957 9636 17969 9639
rect 17092 9608 17969 9636
rect 17092 9596 17098 9608
rect 17957 9605 17969 9608
rect 18003 9605 18015 9639
rect 17957 9599 18015 9605
rect 13728 9590 13780 9596
rect 9033 9571 9091 9577
rect 9033 9537 9045 9571
rect 9079 9537 9091 9571
rect 11514 9568 11520 9580
rect 11475 9540 11520 9568
rect 9033 9531 9091 9537
rect 11514 9528 11520 9540
rect 11572 9528 11578 9580
rect 11701 9571 11759 9577
rect 11701 9537 11713 9571
rect 11747 9568 11759 9571
rect 12434 9568 12440 9580
rect 11747 9540 12440 9568
rect 11747 9537 11759 9540
rect 11701 9531 11759 9537
rect 12434 9528 12440 9540
rect 12492 9528 12498 9580
rect 12618 9568 12624 9580
rect 12579 9540 12624 9568
rect 12618 9528 12624 9540
rect 12676 9528 12682 9580
rect 13078 9568 13084 9580
rect 13039 9540 13084 9568
rect 13078 9528 13084 9540
rect 13136 9528 13142 9580
rect 16942 9528 16948 9580
rect 17000 9568 17006 9580
rect 18800 9568 18828 9676
rect 20530 9636 20536 9648
rect 18892 9608 20392 9636
rect 18892 9577 18920 9608
rect 20364 9580 20392 9608
rect 20456 9608 20536 9636
rect 17000 9540 18828 9568
rect 17000 9528 17006 9540
rect 7006 9500 7012 9512
rect 6748 9472 7012 9500
rect 6641 9463 6699 9469
rect 7006 9460 7012 9472
rect 7064 9500 7070 9512
rect 11532 9500 11560 9528
rect 7064 9472 11560 9500
rect 18800 9500 18828 9540
rect 18877 9571 18935 9577
rect 18877 9537 18889 9571
rect 18923 9537 18935 9571
rect 18877 9531 18935 9537
rect 18969 9571 19027 9577
rect 18969 9537 18981 9571
rect 19015 9537 19027 9571
rect 19150 9568 19156 9580
rect 19111 9540 19156 9568
rect 18969 9531 19027 9537
rect 18984 9500 19012 9531
rect 19150 9528 19156 9540
rect 19208 9528 19214 9580
rect 19245 9571 19303 9577
rect 19245 9537 19257 9571
rect 19291 9537 19303 9571
rect 20346 9568 20352 9580
rect 20307 9540 20352 9568
rect 19245 9531 19303 9537
rect 18800 9472 19012 9500
rect 19260 9500 19288 9531
rect 20346 9528 20352 9540
rect 20404 9528 20410 9580
rect 20456 9577 20484 9608
rect 20530 9596 20536 9608
rect 20588 9596 20594 9648
rect 20640 9636 20668 9676
rect 21928 9676 23296 9704
rect 21928 9636 21956 9676
rect 23290 9664 23296 9676
rect 23348 9664 23354 9716
rect 25317 9707 25375 9713
rect 25317 9673 25329 9707
rect 25363 9673 25375 9707
rect 25317 9667 25375 9673
rect 28583 9707 28641 9713
rect 28583 9673 28595 9707
rect 28629 9704 28641 9707
rect 29086 9704 29092 9716
rect 28629 9676 29092 9704
rect 28629 9673 28641 9676
rect 28583 9667 28641 9673
rect 22922 9636 22928 9648
rect 20640 9608 21956 9636
rect 22883 9608 22928 9636
rect 22922 9596 22928 9608
rect 22980 9596 22986 9648
rect 23382 9636 23388 9648
rect 23032 9608 23388 9636
rect 20441 9571 20499 9577
rect 20441 9537 20453 9571
rect 20487 9537 20499 9571
rect 20622 9568 20628 9580
rect 20583 9540 20628 9568
rect 20441 9531 20499 9537
rect 20622 9528 20628 9540
rect 20680 9528 20686 9580
rect 20714 9528 20720 9580
rect 20772 9568 20778 9580
rect 20772 9540 20817 9568
rect 20772 9528 20778 9540
rect 22646 9528 22652 9580
rect 22704 9577 22710 9580
rect 22704 9571 22753 9577
rect 22704 9537 22707 9571
rect 22741 9537 22753 9571
rect 22704 9531 22753 9537
rect 22809 9571 22867 9577
rect 22809 9537 22821 9571
rect 22855 9568 22867 9571
rect 23032 9568 23060 9608
rect 23382 9596 23388 9608
rect 23440 9636 23446 9648
rect 23845 9639 23903 9645
rect 23845 9636 23857 9639
rect 23440 9608 23857 9636
rect 23440 9596 23446 9608
rect 23845 9605 23857 9608
rect 23891 9605 23903 9639
rect 23845 9599 23903 9605
rect 23937 9639 23995 9645
rect 23937 9605 23949 9639
rect 23983 9605 23995 9639
rect 23937 9599 23995 9605
rect 22855 9540 23060 9568
rect 23109 9571 23167 9577
rect 22855 9537 22867 9540
rect 22809 9531 22867 9537
rect 23109 9537 23121 9571
rect 23155 9568 23167 9571
rect 23290 9568 23296 9580
rect 23155 9540 23296 9568
rect 23155 9537 23167 9540
rect 23109 9531 23167 9537
rect 22704 9528 22710 9531
rect 23290 9528 23296 9540
rect 23348 9528 23354 9580
rect 23658 9528 23664 9580
rect 23716 9577 23722 9580
rect 23716 9571 23765 9577
rect 23716 9537 23719 9571
rect 23753 9537 23765 9571
rect 23716 9531 23765 9537
rect 23716 9528 23722 9531
rect 19260 9472 22692 9500
rect 7064 9460 7070 9472
rect 3050 9392 3056 9444
rect 3108 9392 3114 9444
rect 18141 9435 18199 9441
rect 18141 9401 18153 9435
rect 18187 9432 18199 9435
rect 22278 9432 22284 9444
rect 18187 9404 22284 9432
rect 18187 9401 18199 9404
rect 18141 9395 18199 9401
rect 22278 9392 22284 9404
rect 22336 9392 22342 9444
rect 22664 9432 22692 9472
rect 23569 9435 23627 9441
rect 23569 9432 23581 9435
rect 22664 9404 23581 9432
rect 23569 9401 23581 9404
rect 23615 9401 23627 9435
rect 23952 9432 23980 9599
rect 24026 9596 24032 9648
rect 24084 9636 24090 9648
rect 25332 9636 25360 9667
rect 29086 9664 29092 9676
rect 29144 9664 29150 9716
rect 29730 9664 29736 9716
rect 29788 9704 29794 9716
rect 35342 9704 35348 9716
rect 29788 9676 30052 9704
rect 35303 9676 35348 9704
rect 29788 9664 29794 9676
rect 24084 9608 25360 9636
rect 24084 9596 24090 9608
rect 25590 9596 25596 9648
rect 25648 9636 25654 9648
rect 25648 9608 25693 9636
rect 25792 9608 26648 9636
rect 25648 9596 25654 9608
rect 24121 9571 24179 9577
rect 24121 9537 24133 9571
rect 24167 9568 24179 9571
rect 24670 9568 24676 9580
rect 24167 9540 24256 9568
rect 24631 9540 24676 9568
rect 24167 9537 24179 9540
rect 24121 9531 24179 9537
rect 24228 9512 24256 9540
rect 24670 9528 24676 9540
rect 24728 9528 24734 9580
rect 24762 9528 24768 9580
rect 24820 9568 24826 9580
rect 24857 9571 24915 9577
rect 24857 9568 24869 9571
rect 24820 9540 24869 9568
rect 24820 9528 24826 9540
rect 24857 9537 24869 9540
rect 24903 9537 24915 9571
rect 25498 9568 25504 9580
rect 25459 9540 25504 9568
rect 24857 9531 24915 9537
rect 25498 9528 25504 9540
rect 25556 9528 25562 9580
rect 25682 9528 25688 9580
rect 25740 9568 25746 9580
rect 25792 9568 25820 9608
rect 25869 9571 25927 9577
rect 25740 9540 25833 9568
rect 25740 9528 25746 9540
rect 25869 9537 25881 9571
rect 25915 9568 25927 9571
rect 26510 9568 26516 9580
rect 25915 9540 26516 9568
rect 25915 9537 25927 9540
rect 25869 9531 25927 9537
rect 26510 9528 26516 9540
rect 26568 9528 26574 9580
rect 26620 9568 26648 9608
rect 27338 9596 27344 9648
rect 27396 9636 27402 9648
rect 27433 9639 27491 9645
rect 27433 9636 27445 9639
rect 27396 9608 27445 9636
rect 27396 9596 27402 9608
rect 27433 9605 27445 9608
rect 27479 9636 27491 9639
rect 28718 9636 28724 9648
rect 27479 9608 28724 9636
rect 27479 9605 27491 9608
rect 27433 9599 27491 9605
rect 28718 9596 28724 9608
rect 28776 9636 28782 9648
rect 29362 9636 29368 9648
rect 28776 9608 29368 9636
rect 28776 9596 28782 9608
rect 28626 9568 28632 9580
rect 26620 9540 28632 9568
rect 28626 9528 28632 9540
rect 28684 9528 28690 9580
rect 28828 9577 28856 9608
rect 29362 9596 29368 9608
rect 29420 9596 29426 9648
rect 29454 9596 29460 9648
rect 29512 9636 29518 9648
rect 29914 9636 29920 9648
rect 29512 9608 29920 9636
rect 29512 9596 29518 9608
rect 29914 9596 29920 9608
rect 29972 9596 29978 9648
rect 30024 9645 30052 9676
rect 35342 9664 35348 9676
rect 35400 9664 35406 9716
rect 36081 9707 36139 9713
rect 36081 9673 36093 9707
rect 36127 9673 36139 9707
rect 36081 9667 36139 9673
rect 43073 9707 43131 9713
rect 43073 9673 43085 9707
rect 43119 9673 43131 9707
rect 43073 9667 43131 9673
rect 30009 9639 30067 9645
rect 30009 9605 30021 9639
rect 30055 9605 30067 9639
rect 30009 9599 30067 9605
rect 28813 9571 28871 9577
rect 28813 9537 28825 9571
rect 28859 9537 28871 9571
rect 28813 9531 28871 9537
rect 28994 9528 29000 9580
rect 29052 9568 29058 9580
rect 29822 9577 29828 9580
rect 29641 9571 29699 9577
rect 29641 9568 29653 9571
rect 29052 9540 29653 9568
rect 29052 9528 29058 9540
rect 29641 9537 29653 9540
rect 29687 9537 29699 9571
rect 29641 9531 29699 9537
rect 29789 9571 29828 9577
rect 29789 9537 29801 9571
rect 29789 9531 29828 9537
rect 29822 9528 29828 9531
rect 29880 9528 29886 9580
rect 30106 9571 30164 9577
rect 30106 9537 30118 9571
rect 30152 9537 30164 9571
rect 35360 9568 35388 9664
rect 35894 9596 35900 9648
rect 35952 9636 35958 9648
rect 36096 9636 36124 9667
rect 35952 9608 36124 9636
rect 35952 9596 35958 9608
rect 41506 9596 41512 9648
rect 41564 9636 41570 9648
rect 42702 9636 42708 9648
rect 41564 9608 41920 9636
rect 42663 9608 42708 9636
rect 41564 9596 41570 9608
rect 35989 9571 36047 9577
rect 35989 9568 36001 9571
rect 35360 9540 36001 9568
rect 30106 9531 30164 9537
rect 35989 9537 36001 9540
rect 36035 9537 36047 9571
rect 36354 9568 36360 9580
rect 36315 9540 36360 9568
rect 35989 9531 36047 9537
rect 24210 9460 24216 9512
rect 24268 9500 24274 9512
rect 26050 9500 26056 9512
rect 24268 9472 26056 9500
rect 24268 9460 24274 9472
rect 26050 9460 26056 9472
rect 26108 9460 26114 9512
rect 27430 9460 27436 9512
rect 27488 9500 27494 9512
rect 29454 9500 29460 9512
rect 27488 9472 29460 9500
rect 27488 9460 27494 9472
rect 29454 9460 29460 9472
rect 29512 9500 29518 9512
rect 30121 9500 30149 9531
rect 36354 9528 36360 9540
rect 36412 9528 36418 9580
rect 41690 9568 41696 9580
rect 41651 9540 41696 9568
rect 41690 9528 41696 9540
rect 41748 9528 41754 9580
rect 41892 9577 41920 9608
rect 42702 9596 42708 9608
rect 42760 9596 42766 9648
rect 42910 9639 42968 9645
rect 42910 9605 42922 9639
rect 42956 9636 42968 9639
rect 43088 9636 43116 9667
rect 55122 9664 55128 9716
rect 55180 9704 55186 9716
rect 55217 9707 55275 9713
rect 55217 9704 55229 9707
rect 55180 9676 55229 9704
rect 55180 9664 55186 9676
rect 55217 9673 55229 9676
rect 55263 9673 55275 9707
rect 55217 9667 55275 9673
rect 43993 9639 44051 9645
rect 43993 9636 44005 9639
rect 42956 9608 43024 9636
rect 43088 9608 44005 9636
rect 42956 9605 42968 9608
rect 42910 9599 42968 9605
rect 41877 9571 41935 9577
rect 41877 9537 41889 9571
rect 41923 9537 41935 9571
rect 42996 9568 43024 9608
rect 43993 9605 44005 9608
rect 44039 9605 44051 9639
rect 44174 9636 44180 9648
rect 44135 9608 44180 9636
rect 43993 9599 44051 9605
rect 44174 9596 44180 9608
rect 44232 9636 44238 9648
rect 44232 9608 44864 9636
rect 44232 9596 44238 9608
rect 43162 9568 43168 9580
rect 42996 9540 43168 9568
rect 41877 9531 41935 9537
rect 43162 9528 43168 9540
rect 43220 9528 43226 9580
rect 44836 9577 44864 9608
rect 44821 9571 44879 9577
rect 44821 9537 44833 9571
rect 44867 9537 44879 9571
rect 44821 9531 44879 9537
rect 45465 9571 45523 9577
rect 45465 9537 45477 9571
rect 45511 9568 45523 9571
rect 45554 9568 45560 9580
rect 45511 9540 45560 9568
rect 45511 9537 45523 9540
rect 45465 9531 45523 9537
rect 45554 9528 45560 9540
rect 45612 9528 45618 9580
rect 45830 9568 45836 9580
rect 45791 9540 45836 9568
rect 45830 9528 45836 9540
rect 45888 9528 45894 9580
rect 46014 9568 46020 9580
rect 45975 9540 46020 9568
rect 46014 9528 46020 9540
rect 46072 9528 46078 9580
rect 54018 9568 54024 9580
rect 53979 9540 54024 9568
rect 54018 9528 54024 9540
rect 54076 9528 54082 9580
rect 55125 9571 55183 9577
rect 55125 9537 55137 9571
rect 55171 9537 55183 9571
rect 55306 9568 55312 9580
rect 55267 9540 55312 9568
rect 55125 9531 55183 9537
rect 36538 9500 36544 9512
rect 29512 9472 30149 9500
rect 36499 9472 36544 9500
rect 29512 9460 29518 9472
rect 36538 9460 36544 9472
rect 36596 9460 36602 9512
rect 55140 9500 55168 9531
rect 55306 9528 55312 9540
rect 55364 9568 55370 9580
rect 55950 9568 55956 9580
rect 55364 9540 55956 9568
rect 55364 9528 55370 9540
rect 55582 9500 55588 9512
rect 55140 9472 55588 9500
rect 55582 9460 55588 9472
rect 55640 9460 55646 9512
rect 55876 9509 55904 9540
rect 55950 9528 55956 9540
rect 56008 9528 56014 9580
rect 55861 9503 55919 9509
rect 55861 9469 55873 9503
rect 55907 9469 55919 9503
rect 55861 9463 55919 9469
rect 56226 9460 56232 9512
rect 56284 9500 56290 9512
rect 56321 9503 56379 9509
rect 56321 9500 56333 9503
rect 56284 9472 56333 9500
rect 56284 9460 56290 9472
rect 56321 9469 56333 9472
rect 56367 9469 56379 9503
rect 56321 9463 56379 9469
rect 24302 9432 24308 9444
rect 23952 9404 24308 9432
rect 23569 9395 23627 9401
rect 24302 9392 24308 9404
rect 24360 9432 24366 9444
rect 25682 9432 25688 9444
rect 24360 9404 25688 9432
rect 24360 9392 24366 9404
rect 25682 9392 25688 9404
rect 25740 9392 25746 9444
rect 44913 9435 44971 9441
rect 44913 9432 44925 9435
rect 29840 9404 44925 9432
rect 4433 9367 4491 9373
rect 4433 9333 4445 9367
rect 4479 9364 4491 9367
rect 4706 9364 4712 9376
rect 4479 9336 4712 9364
rect 4479 9333 4491 9336
rect 4433 9327 4491 9333
rect 4706 9324 4712 9336
rect 4764 9324 4770 9376
rect 10870 9324 10876 9376
rect 10928 9364 10934 9376
rect 11609 9367 11667 9373
rect 11609 9364 11621 9367
rect 10928 9336 11621 9364
rect 10928 9324 10934 9336
rect 11609 9333 11621 9336
rect 11655 9333 11667 9367
rect 15838 9364 15844 9376
rect 15799 9336 15844 9364
rect 11609 9327 11667 9333
rect 15838 9324 15844 9336
rect 15896 9324 15902 9376
rect 15930 9324 15936 9376
rect 15988 9364 15994 9376
rect 18693 9367 18751 9373
rect 18693 9364 18705 9367
rect 15988 9336 18705 9364
rect 15988 9324 15994 9336
rect 18693 9333 18705 9336
rect 18739 9333 18751 9367
rect 20162 9364 20168 9376
rect 20123 9336 20168 9364
rect 18693 9327 18751 9333
rect 20162 9324 20168 9336
rect 20220 9324 20226 9376
rect 22462 9324 22468 9376
rect 22520 9364 22526 9376
rect 22557 9367 22615 9373
rect 22557 9364 22569 9367
rect 22520 9336 22569 9364
rect 22520 9324 22526 9336
rect 22557 9333 22569 9336
rect 22603 9333 22615 9367
rect 24854 9364 24860 9376
rect 24815 9336 24860 9364
rect 22557 9327 22615 9333
rect 24854 9324 24860 9336
rect 24912 9324 24918 9376
rect 26878 9324 26884 9376
rect 26936 9364 26942 9376
rect 29840 9364 29868 9404
rect 44913 9401 44925 9404
rect 44959 9401 44971 9435
rect 55125 9435 55183 9441
rect 55125 9432 55137 9435
rect 44913 9395 44971 9401
rect 54312 9404 55137 9432
rect 26936 9336 29868 9364
rect 30285 9367 30343 9373
rect 26936 9324 26942 9336
rect 30285 9333 30297 9367
rect 30331 9364 30343 9367
rect 30558 9364 30564 9376
rect 30331 9336 30564 9364
rect 30331 9333 30343 9336
rect 30285 9327 30343 9333
rect 30558 9324 30564 9336
rect 30616 9324 30622 9376
rect 41785 9367 41843 9373
rect 41785 9333 41797 9367
rect 41831 9364 41843 9367
rect 42518 9364 42524 9376
rect 41831 9336 42524 9364
rect 41831 9333 41843 9336
rect 41785 9327 41843 9333
rect 42518 9324 42524 9336
rect 42576 9324 42582 9376
rect 42886 9364 42892 9376
rect 42847 9336 42892 9364
rect 42886 9324 42892 9336
rect 42944 9324 42950 9376
rect 44361 9367 44419 9373
rect 44361 9333 44373 9367
rect 44407 9364 44419 9367
rect 45922 9364 45928 9376
rect 44407 9336 45928 9364
rect 44407 9333 44419 9336
rect 44361 9327 44419 9333
rect 45922 9324 45928 9336
rect 45980 9324 45986 9376
rect 54312 9373 54340 9404
rect 55125 9401 55137 9404
rect 55171 9401 55183 9435
rect 55125 9395 55183 9401
rect 56045 9435 56103 9441
rect 56045 9401 56057 9435
rect 56091 9432 56103 9435
rect 56134 9432 56140 9444
rect 56091 9404 56140 9432
rect 56091 9401 56103 9404
rect 56045 9395 56103 9401
rect 56134 9392 56140 9404
rect 56192 9392 56198 9444
rect 54297 9367 54355 9373
rect 54297 9333 54309 9367
rect 54343 9333 54355 9367
rect 54478 9364 54484 9376
rect 54439 9336 54484 9364
rect 54297 9327 54355 9333
rect 54478 9324 54484 9336
rect 54536 9324 54542 9376
rect 1104 9274 58880 9296
rect 1104 9222 4214 9274
rect 4266 9222 4278 9274
rect 4330 9222 4342 9274
rect 4394 9222 4406 9274
rect 4458 9222 4470 9274
rect 4522 9222 34934 9274
rect 34986 9222 34998 9274
rect 35050 9222 35062 9274
rect 35114 9222 35126 9274
rect 35178 9222 35190 9274
rect 35242 9222 58880 9274
rect 1104 9200 58880 9222
rect 3234 9160 3240 9172
rect 3195 9132 3240 9160
rect 3234 9120 3240 9132
rect 3292 9120 3298 9172
rect 4062 9120 4068 9172
rect 4120 9160 4126 9172
rect 4157 9163 4215 9169
rect 4157 9160 4169 9163
rect 4120 9132 4169 9160
rect 4120 9120 4126 9132
rect 4157 9129 4169 9132
rect 4203 9129 4215 9163
rect 6546 9160 6552 9172
rect 6507 9132 6552 9160
rect 4157 9123 4215 9129
rect 6546 9120 6552 9132
rect 6604 9120 6610 9172
rect 8202 9160 8208 9172
rect 8163 9132 8208 9160
rect 8202 9120 8208 9132
rect 8260 9120 8266 9172
rect 8846 9120 8852 9172
rect 8904 9160 8910 9172
rect 8941 9163 8999 9169
rect 8941 9160 8953 9163
rect 8904 9132 8953 9160
rect 8904 9120 8910 9132
rect 8941 9129 8953 9132
rect 8987 9129 8999 9163
rect 8941 9123 8999 9129
rect 20349 9163 20407 9169
rect 20349 9129 20361 9163
rect 20395 9160 20407 9163
rect 20622 9160 20628 9172
rect 20395 9132 20628 9160
rect 20395 9129 20407 9132
rect 20349 9123 20407 9129
rect 20622 9120 20628 9132
rect 20680 9120 20686 9172
rect 25498 9120 25504 9172
rect 25556 9160 25562 9172
rect 28994 9160 29000 9172
rect 25556 9132 27752 9160
rect 28955 9132 29000 9160
rect 25556 9120 25562 9132
rect 10505 9095 10563 9101
rect 10505 9061 10517 9095
rect 10551 9061 10563 9095
rect 10505 9055 10563 9061
rect 8570 9024 8576 9036
rect 8220 8996 8576 9024
rect 2869 8959 2927 8965
rect 2869 8925 2881 8959
rect 2915 8956 2927 8959
rect 3142 8956 3148 8968
rect 2915 8928 3148 8956
rect 2915 8925 2927 8928
rect 2869 8919 2927 8925
rect 3142 8916 3148 8928
rect 3200 8956 3206 8968
rect 3602 8956 3608 8968
rect 3200 8928 3608 8956
rect 3200 8916 3206 8928
rect 3602 8916 3608 8928
rect 3660 8916 3666 8968
rect 6365 8959 6423 8965
rect 6365 8925 6377 8959
rect 6411 8956 6423 8959
rect 6454 8956 6460 8968
rect 6411 8928 6460 8956
rect 6411 8925 6423 8928
rect 6365 8919 6423 8925
rect 6454 8916 6460 8928
rect 6512 8916 6518 8968
rect 6549 8959 6607 8965
rect 6549 8925 6561 8959
rect 6595 8956 6607 8959
rect 6914 8956 6920 8968
rect 6595 8928 6920 8956
rect 6595 8925 6607 8928
rect 6549 8919 6607 8925
rect 6914 8916 6920 8928
rect 6972 8916 6978 8968
rect 8220 8965 8248 8996
rect 8570 8984 8576 8996
rect 8628 9024 8634 9036
rect 9401 9027 9459 9033
rect 9401 9024 9413 9027
rect 8628 8996 9413 9024
rect 8628 8984 8634 8996
rect 9401 8993 9413 8996
rect 9447 9024 9459 9027
rect 10042 9024 10048 9036
rect 9447 8996 10048 9024
rect 9447 8993 9459 8996
rect 9401 8987 9459 8993
rect 10042 8984 10048 8996
rect 10100 8984 10106 9036
rect 8205 8959 8263 8965
rect 8205 8925 8217 8959
rect 8251 8925 8263 8959
rect 8205 8919 8263 8925
rect 8389 8959 8447 8965
rect 8389 8925 8401 8959
rect 8435 8956 8447 8959
rect 9309 8959 9367 8965
rect 9309 8956 9321 8959
rect 8435 8928 9321 8956
rect 8435 8925 8447 8928
rect 8389 8919 8447 8925
rect 9309 8925 9321 8928
rect 9355 8956 9367 8959
rect 10520 8956 10548 9055
rect 10594 9052 10600 9104
rect 10652 9092 10658 9104
rect 24397 9095 24455 9101
rect 24397 9092 24409 9095
rect 10652 9064 20392 9092
rect 10652 9052 10658 9064
rect 10962 9024 10968 9036
rect 10923 8996 10968 9024
rect 10962 8984 10968 8996
rect 11020 8984 11026 9036
rect 15105 9027 15163 9033
rect 15105 8993 15117 9027
rect 15151 9024 15163 9027
rect 15930 9024 15936 9036
rect 15151 8996 15936 9024
rect 15151 8993 15163 8996
rect 15105 8987 15163 8993
rect 15930 8984 15936 8996
rect 15988 8984 15994 9036
rect 17494 9024 17500 9036
rect 17455 8996 17500 9024
rect 17494 8984 17500 8996
rect 17552 8984 17558 9036
rect 10870 8956 10876 8968
rect 9355 8928 10548 8956
rect 10831 8928 10876 8956
rect 9355 8925 9367 8928
rect 9309 8919 9367 8925
rect 10870 8916 10876 8928
rect 10928 8916 10934 8968
rect 14918 8916 14924 8968
rect 14976 8956 14982 8968
rect 15013 8959 15071 8965
rect 15013 8956 15025 8959
rect 14976 8928 15025 8956
rect 14976 8916 14982 8928
rect 15013 8925 15025 8928
rect 15059 8925 15071 8959
rect 15013 8919 15071 8925
rect 16761 8959 16819 8965
rect 16761 8925 16773 8959
rect 16807 8956 16819 8959
rect 17218 8956 17224 8968
rect 16807 8928 17224 8956
rect 16807 8925 16819 8928
rect 16761 8919 16819 8925
rect 3050 8888 3056 8900
rect 3011 8860 3056 8888
rect 3050 8848 3056 8860
rect 3108 8848 3114 8900
rect 3786 8888 3792 8900
rect 3747 8860 3792 8888
rect 3786 8848 3792 8860
rect 3844 8848 3850 8900
rect 3878 8848 3884 8900
rect 3936 8888 3942 8900
rect 3973 8891 4031 8897
rect 3973 8888 3985 8891
rect 3936 8860 3985 8888
rect 3936 8848 3942 8860
rect 3973 8857 3985 8860
rect 4019 8857 4031 8891
rect 10042 8888 10048 8900
rect 10003 8860 10048 8888
rect 3973 8851 4031 8857
rect 10042 8848 10048 8860
rect 10100 8848 10106 8900
rect 15028 8888 15056 8919
rect 17218 8916 17224 8928
rect 17276 8956 17282 8968
rect 17405 8959 17463 8965
rect 17405 8956 17417 8959
rect 17276 8928 17417 8956
rect 17276 8916 17282 8928
rect 17405 8925 17417 8928
rect 17451 8925 17463 8959
rect 17405 8919 17463 8925
rect 19242 8916 19248 8968
rect 19300 8956 19306 8968
rect 19337 8959 19395 8965
rect 19337 8956 19349 8959
rect 19300 8928 19349 8956
rect 19300 8916 19306 8928
rect 19337 8925 19349 8928
rect 19383 8925 19395 8959
rect 19518 8956 19524 8968
rect 19479 8928 19524 8956
rect 19337 8919 19395 8925
rect 19518 8916 19524 8928
rect 19576 8916 19582 8968
rect 20165 8959 20223 8965
rect 20165 8925 20177 8959
rect 20211 8956 20223 8959
rect 20254 8956 20260 8968
rect 20211 8928 20260 8956
rect 20211 8925 20223 8928
rect 20165 8919 20223 8925
rect 20254 8916 20260 8928
rect 20312 8916 20318 8968
rect 20364 8965 20392 9064
rect 20824 9064 24409 9092
rect 20824 8965 20852 9064
rect 24397 9061 24409 9064
rect 24443 9092 24455 9095
rect 24670 9092 24676 9104
rect 24443 9064 24676 9092
rect 24443 9061 24455 9064
rect 24397 9055 24455 9061
rect 24670 9052 24676 9064
rect 24728 9092 24734 9104
rect 25590 9092 25596 9104
rect 24728 9064 25596 9092
rect 24728 9052 24734 9064
rect 25590 9052 25596 9064
rect 25648 9052 25654 9104
rect 20898 8984 20904 9036
rect 20956 9024 20962 9036
rect 24210 9024 24216 9036
rect 20956 8996 24216 9024
rect 20956 8984 20962 8996
rect 20349 8959 20407 8965
rect 20349 8925 20361 8959
rect 20395 8956 20407 8959
rect 20809 8959 20867 8965
rect 20809 8956 20821 8959
rect 20395 8928 20821 8956
rect 20395 8925 20407 8928
rect 20349 8919 20407 8925
rect 20809 8925 20821 8928
rect 20855 8925 20867 8959
rect 22462 8956 22468 8968
rect 22423 8928 22468 8956
rect 20809 8919 20867 8925
rect 22462 8916 22468 8928
rect 22520 8916 22526 8968
rect 22756 8965 22784 8996
rect 24210 8984 24216 8996
rect 24268 8984 24274 9036
rect 24854 8984 24860 9036
rect 24912 9024 24918 9036
rect 24912 8996 27384 9024
rect 24912 8984 24918 8996
rect 22557 8959 22615 8965
rect 22557 8925 22569 8959
rect 22603 8925 22615 8959
rect 22557 8919 22615 8925
rect 22741 8959 22799 8965
rect 22741 8925 22753 8959
rect 22787 8925 22799 8959
rect 22741 8919 22799 8925
rect 22833 8959 22891 8965
rect 22833 8925 22845 8959
rect 22879 8925 22891 8959
rect 22833 8919 22891 8925
rect 15838 8888 15844 8900
rect 15028 8860 15844 8888
rect 15838 8848 15844 8860
rect 15896 8888 15902 8900
rect 19429 8891 19487 8897
rect 15896 8860 17908 8888
rect 15896 8848 15902 8860
rect 14185 8823 14243 8829
rect 14185 8789 14197 8823
rect 14231 8820 14243 8823
rect 14458 8820 14464 8832
rect 14231 8792 14464 8820
rect 14231 8789 14243 8792
rect 14185 8783 14243 8789
rect 14458 8780 14464 8792
rect 14516 8780 14522 8832
rect 17678 8780 17684 8832
rect 17736 8820 17742 8832
rect 17773 8823 17831 8829
rect 17773 8820 17785 8823
rect 17736 8792 17785 8820
rect 17736 8780 17742 8792
rect 17773 8789 17785 8792
rect 17819 8789 17831 8823
rect 17880 8820 17908 8860
rect 19429 8857 19441 8891
rect 19475 8888 19487 8891
rect 22572 8888 22600 8919
rect 19475 8860 22600 8888
rect 22848 8888 22876 8919
rect 23014 8916 23020 8968
rect 23072 8956 23078 8968
rect 24949 8959 25007 8965
rect 24949 8956 24961 8959
rect 23072 8928 24961 8956
rect 23072 8916 23078 8928
rect 24949 8925 24961 8928
rect 24995 8925 25007 8959
rect 24949 8919 25007 8925
rect 25038 8916 25044 8968
rect 25096 8956 25102 8968
rect 25225 8959 25283 8965
rect 25225 8956 25237 8959
rect 25096 8928 25237 8956
rect 25096 8916 25102 8928
rect 25225 8925 25237 8928
rect 25271 8925 25283 8959
rect 25225 8919 25283 8925
rect 25240 8888 25268 8919
rect 26050 8916 26056 8968
rect 26108 8956 26114 8968
rect 26237 8959 26295 8965
rect 26237 8956 26249 8959
rect 26108 8928 26249 8956
rect 26108 8916 26114 8928
rect 26237 8925 26249 8928
rect 26283 8925 26295 8959
rect 26237 8919 26295 8925
rect 26326 8916 26332 8968
rect 26384 8956 26390 8968
rect 26605 8959 26663 8965
rect 26605 8956 26617 8959
rect 26384 8928 26617 8956
rect 26384 8916 26390 8928
rect 26605 8925 26617 8928
rect 26651 8925 26663 8959
rect 27246 8956 27252 8968
rect 27207 8928 27252 8956
rect 26605 8919 26663 8925
rect 27246 8916 27252 8928
rect 27304 8916 27310 8968
rect 27356 8965 27384 8996
rect 27341 8959 27399 8965
rect 27341 8925 27353 8959
rect 27387 8925 27399 8959
rect 27522 8956 27528 8968
rect 27483 8928 27528 8956
rect 27341 8919 27399 8925
rect 27522 8916 27528 8928
rect 27580 8916 27586 8968
rect 27617 8959 27675 8965
rect 27617 8925 27629 8959
rect 27663 8925 27675 8959
rect 27617 8919 27675 8925
rect 26421 8891 26479 8897
rect 26421 8888 26433 8891
rect 22848 8860 25176 8888
rect 25240 8860 26433 8888
rect 19475 8857 19487 8860
rect 19429 8851 19487 8857
rect 20254 8820 20260 8832
rect 17880 8792 20260 8820
rect 17773 8783 17831 8789
rect 20254 8780 20260 8792
rect 20312 8780 20318 8832
rect 22278 8780 22284 8832
rect 22336 8820 22342 8832
rect 22848 8820 22876 8860
rect 22336 8792 22876 8820
rect 22336 8780 22342 8792
rect 23014 8780 23020 8832
rect 23072 8820 23078 8832
rect 25148 8820 25176 8860
rect 26421 8857 26433 8860
rect 26467 8857 26479 8891
rect 26421 8851 26479 8857
rect 26510 8848 26516 8900
rect 26568 8888 26574 8900
rect 27632 8888 27660 8919
rect 26568 8860 26613 8888
rect 26712 8860 27660 8888
rect 26568 8848 26574 8860
rect 26712 8820 26740 8860
rect 27356 8832 27384 8860
rect 23072 8792 23117 8820
rect 25148 8792 26740 8820
rect 26789 8823 26847 8829
rect 23072 8780 23078 8792
rect 26789 8789 26801 8823
rect 26835 8820 26847 8823
rect 27246 8820 27252 8832
rect 26835 8792 27252 8820
rect 26835 8789 26847 8792
rect 26789 8783 26847 8789
rect 27246 8780 27252 8792
rect 27304 8780 27310 8832
rect 27338 8780 27344 8832
rect 27396 8780 27402 8832
rect 27724 8820 27752 9132
rect 28994 9120 29000 9132
rect 29052 9120 29058 9172
rect 29086 9120 29092 9172
rect 29144 9160 29150 9172
rect 30561 9163 30619 9169
rect 29144 9132 29776 9160
rect 29144 9120 29150 9132
rect 27801 9095 27859 9101
rect 27801 9061 27813 9095
rect 27847 9092 27859 9095
rect 29638 9092 29644 9104
rect 27847 9064 29644 9092
rect 27847 9061 27859 9064
rect 27801 9055 27859 9061
rect 29638 9052 29644 9064
rect 29696 9052 29702 9104
rect 29748 9024 29776 9132
rect 30561 9129 30573 9163
rect 30607 9160 30619 9163
rect 33226 9160 33232 9172
rect 30607 9132 33232 9160
rect 30607 9129 30619 9132
rect 30561 9123 30619 9129
rect 33226 9120 33232 9132
rect 33284 9120 33290 9172
rect 36354 9120 36360 9172
rect 36412 9160 36418 9172
rect 37461 9163 37519 9169
rect 37461 9160 37473 9163
rect 36412 9132 37473 9160
rect 36412 9120 36418 9132
rect 37461 9129 37473 9132
rect 37507 9129 37519 9163
rect 37461 9123 37519 9129
rect 42889 9163 42947 9169
rect 42889 9129 42901 9163
rect 42935 9160 42947 9163
rect 43162 9160 43168 9172
rect 42935 9132 43168 9160
rect 42935 9129 42947 9132
rect 42889 9123 42947 9129
rect 43162 9120 43168 9132
rect 43220 9120 43226 9172
rect 54018 9120 54024 9172
rect 54076 9160 54082 9172
rect 54389 9163 54447 9169
rect 54389 9160 54401 9163
rect 54076 9132 54401 9160
rect 54076 9120 54082 9132
rect 54389 9129 54401 9132
rect 54435 9129 54447 9163
rect 54389 9123 54447 9129
rect 32769 9095 32827 9101
rect 32769 9061 32781 9095
rect 32815 9061 32827 9095
rect 32769 9055 32827 9061
rect 28460 8996 29592 9024
rect 29748 8996 29832 9024
rect 28460 8965 28488 8996
rect 28445 8959 28503 8965
rect 28445 8925 28457 8959
rect 28491 8925 28503 8959
rect 28626 8956 28632 8968
rect 28587 8928 28632 8956
rect 28445 8919 28503 8925
rect 28460 8888 28488 8919
rect 28626 8916 28632 8928
rect 28684 8916 28690 8968
rect 29564 8965 29592 8996
rect 29804 8965 29832 8996
rect 30926 8984 30932 9036
rect 30984 9024 30990 9036
rect 32309 9027 32367 9033
rect 32309 9024 32321 9027
rect 30984 8996 32321 9024
rect 30984 8984 30990 8996
rect 32309 8993 32321 8996
rect 32355 8993 32367 9027
rect 32784 9024 32812 9055
rect 33134 9052 33140 9104
rect 33192 9092 33198 9104
rect 33321 9095 33379 9101
rect 33321 9092 33333 9095
rect 33192 9064 33333 9092
rect 33192 9052 33198 9064
rect 33321 9061 33333 9064
rect 33367 9061 33379 9095
rect 36722 9092 36728 9104
rect 36683 9064 36728 9092
rect 33321 9055 33379 9061
rect 36722 9052 36728 9064
rect 36780 9052 36786 9104
rect 36909 9095 36967 9101
rect 36909 9061 36921 9095
rect 36955 9092 36967 9095
rect 40126 9092 40132 9104
rect 36955 9064 40132 9092
rect 36955 9061 36967 9064
rect 36909 9055 36967 9061
rect 40126 9052 40132 9064
rect 40184 9092 40190 9104
rect 45554 9092 45560 9104
rect 40184 9064 40540 9092
rect 40184 9052 40190 9064
rect 34606 9024 34612 9036
rect 32784 8996 34612 9024
rect 32309 8987 32367 8993
rect 34606 8984 34612 8996
rect 34664 9024 34670 9036
rect 34664 8996 34928 9024
rect 34664 8984 34670 8996
rect 28813 8959 28871 8965
rect 28534 8888 28540 8900
rect 28460 8860 28540 8888
rect 28534 8848 28540 8860
rect 28592 8848 28598 8900
rect 28718 8897 28724 8946
rect 28717 8894 28724 8897
rect 28776 8894 28782 8946
rect 28813 8925 28825 8959
rect 28859 8925 28871 8959
rect 28813 8919 28871 8925
rect 29549 8959 29607 8965
rect 29549 8925 29561 8959
rect 29595 8925 29607 8959
rect 29804 8959 29875 8965
rect 29804 8928 29829 8959
rect 29549 8919 29607 8925
rect 29817 8925 29829 8928
rect 29863 8925 29875 8959
rect 29817 8919 29875 8925
rect 29917 8959 29975 8965
rect 29917 8925 29929 8959
rect 29963 8925 29975 8959
rect 30834 8956 30840 8968
rect 30795 8928 30840 8956
rect 29917 8919 29975 8925
rect 28717 8891 28775 8894
rect 28717 8857 28729 8891
rect 28763 8857 28775 8891
rect 28717 8851 28775 8857
rect 28828 8820 28856 8919
rect 28902 8848 28908 8900
rect 28960 8888 28966 8900
rect 28960 8848 28994 8888
rect 29454 8848 29460 8900
rect 29512 8888 29518 8900
rect 29733 8891 29791 8897
rect 29733 8888 29745 8891
rect 29512 8860 29745 8888
rect 29512 8848 29518 8860
rect 29733 8857 29745 8860
rect 29779 8857 29791 8891
rect 29733 8851 29791 8857
rect 27724 8792 28856 8820
rect 28966 8820 28994 8848
rect 29932 8820 29960 8919
rect 30834 8916 30840 8928
rect 30892 8956 30898 8968
rect 32122 8956 32128 8968
rect 30892 8928 32128 8956
rect 30892 8916 30898 8928
rect 32122 8916 32128 8928
rect 32180 8916 32186 8968
rect 32401 8959 32459 8965
rect 32401 8925 32413 8959
rect 32447 8956 32459 8959
rect 33134 8956 33140 8968
rect 32447 8928 33140 8956
rect 32447 8925 32459 8928
rect 32401 8919 32459 8925
rect 33134 8916 33140 8928
rect 33192 8916 33198 8968
rect 33686 8916 33692 8968
rect 33744 8956 33750 8968
rect 34422 8956 34428 8968
rect 33744 8928 34428 8956
rect 33744 8916 33750 8928
rect 34422 8916 34428 8928
rect 34480 8956 34486 8968
rect 34793 8959 34851 8965
rect 34793 8956 34805 8959
rect 34480 8928 34805 8956
rect 34480 8916 34486 8928
rect 34793 8925 34805 8928
rect 34839 8925 34851 8959
rect 34900 8942 34928 8996
rect 35894 8984 35900 9036
rect 35952 9024 35958 9036
rect 36262 9024 36268 9036
rect 35952 8996 36268 9024
rect 35952 8984 35958 8996
rect 36262 8984 36268 8996
rect 36320 9024 36326 9036
rect 36449 9027 36507 9033
rect 36449 9024 36461 9027
rect 36320 8996 36461 9024
rect 36320 8984 36326 8996
rect 36449 8993 36461 8996
rect 36495 8993 36507 9027
rect 36449 8987 36507 8993
rect 37829 9027 37887 9033
rect 37829 8993 37841 9027
rect 37875 9024 37887 9027
rect 37918 9024 37924 9036
rect 37875 8996 37924 9024
rect 37875 8993 37887 8996
rect 37829 8987 37887 8993
rect 37918 8984 37924 8996
rect 37976 9024 37982 9036
rect 38286 9024 38292 9036
rect 37976 8996 38292 9024
rect 37976 8984 37982 8996
rect 38286 8984 38292 8996
rect 38344 8984 38350 9036
rect 35805 8959 35863 8965
rect 34793 8919 34851 8925
rect 35805 8925 35817 8959
rect 35851 8956 35863 8959
rect 37550 8956 37556 8968
rect 35851 8928 37556 8956
rect 35851 8925 35863 8928
rect 35805 8919 35863 8925
rect 37550 8916 37556 8928
rect 37608 8956 37614 8968
rect 40512 8965 40540 9064
rect 45112 9064 45560 9092
rect 45112 9033 45140 9064
rect 45554 9052 45560 9064
rect 45612 9052 45618 9104
rect 46014 9092 46020 9104
rect 45664 9064 46020 9092
rect 45097 9027 45155 9033
rect 45097 8993 45109 9027
rect 45143 8993 45155 9027
rect 45664 9024 45692 9064
rect 46014 9052 46020 9064
rect 46072 9052 46078 9104
rect 45830 9024 45836 9036
rect 45097 8987 45155 8993
rect 45388 8996 45692 9024
rect 45791 8996 45836 9024
rect 37645 8959 37703 8965
rect 37645 8956 37657 8959
rect 37608 8928 37657 8956
rect 37608 8916 37614 8928
rect 37645 8925 37657 8928
rect 37691 8925 37703 8959
rect 37645 8919 37703 8925
rect 40497 8959 40555 8965
rect 40497 8925 40509 8959
rect 40543 8925 40555 8959
rect 41046 8956 41052 8968
rect 41007 8928 41052 8956
rect 40497 8919 40555 8925
rect 41046 8916 41052 8928
rect 41104 8916 41110 8968
rect 45388 8956 45416 8996
rect 45830 8984 45836 8996
rect 45888 8984 45894 9036
rect 49142 9024 49148 9036
rect 49103 8996 49148 9024
rect 49142 8984 49148 8996
rect 49200 8984 49206 9036
rect 51810 9024 51816 9036
rect 51771 8996 51816 9024
rect 51810 8984 51816 8996
rect 51868 8984 51874 9036
rect 52089 9027 52147 9033
rect 52089 8993 52101 9027
rect 52135 9024 52147 9027
rect 55582 9024 55588 9036
rect 52135 8996 55588 9024
rect 52135 8993 52147 8996
rect 52089 8987 52147 8993
rect 41984 8942 45416 8956
rect 41984 8928 45402 8942
rect 30561 8891 30619 8897
rect 30561 8857 30573 8891
rect 30607 8857 30619 8891
rect 30742 8888 30748 8900
rect 30703 8860 30748 8888
rect 30561 8851 30619 8857
rect 28966 8792 29960 8820
rect 30101 8823 30159 8829
rect 30101 8789 30113 8823
rect 30147 8820 30159 8823
rect 30576 8820 30604 8851
rect 30742 8848 30748 8860
rect 30800 8848 30806 8900
rect 41984 8874 42012 8928
rect 48682 8916 48688 8968
rect 48740 8956 48746 8968
rect 48958 8956 48964 8968
rect 48740 8928 48964 8956
rect 48740 8916 48746 8928
rect 48958 8916 48964 8928
rect 49016 8956 49022 8968
rect 49237 8959 49295 8965
rect 49237 8956 49249 8959
rect 49016 8928 49249 8956
rect 49016 8916 49022 8928
rect 49237 8925 49249 8928
rect 49283 8925 49295 8959
rect 51442 8956 51448 8968
rect 49237 8919 49295 8925
rect 51046 8928 51448 8956
rect 30147 8792 30604 8820
rect 38933 8823 38991 8829
rect 30147 8789 30159 8792
rect 30101 8783 30159 8789
rect 38933 8789 38945 8823
rect 38979 8820 38991 8823
rect 39666 8820 39672 8832
rect 38979 8792 39672 8820
rect 38979 8789 38991 8792
rect 38933 8783 38991 8789
rect 39666 8780 39672 8792
rect 39724 8780 39730 8832
rect 49605 8823 49663 8829
rect 49605 8789 49617 8823
rect 49651 8820 49663 8823
rect 51046 8820 51074 8928
rect 51442 8916 51448 8928
rect 51500 8956 51506 8968
rect 54312 8965 54340 8996
rect 55582 8984 55588 8996
rect 55640 8984 55646 9036
rect 56134 8984 56140 9036
rect 56192 9024 56198 9036
rect 56192 8996 56456 9024
rect 56192 8984 56198 8996
rect 51721 8959 51779 8965
rect 51721 8956 51733 8959
rect 51500 8928 51733 8956
rect 51500 8916 51506 8928
rect 51721 8925 51733 8928
rect 51767 8925 51779 8959
rect 51721 8919 51779 8925
rect 54297 8959 54355 8965
rect 54297 8925 54309 8959
rect 54343 8925 54355 8959
rect 54297 8919 54355 8925
rect 54481 8959 54539 8965
rect 54481 8925 54493 8959
rect 54527 8956 54539 8959
rect 55306 8956 55312 8968
rect 54527 8928 55312 8956
rect 54527 8925 54539 8928
rect 54481 8919 54539 8925
rect 55306 8916 55312 8928
rect 55364 8916 55370 8968
rect 56226 8956 56232 8968
rect 56187 8928 56232 8956
rect 56226 8916 56232 8928
rect 56284 8916 56290 8968
rect 56428 8965 56456 8996
rect 56778 8984 56784 9036
rect 56836 9024 56842 9036
rect 57149 9027 57207 9033
rect 57149 9024 57161 9027
rect 56836 8996 57161 9024
rect 56836 8984 56842 8996
rect 57149 8993 57161 8996
rect 57195 8993 57207 9027
rect 57149 8987 57207 8993
rect 56413 8959 56471 8965
rect 56413 8925 56425 8959
rect 56459 8925 56471 8959
rect 56413 8919 56471 8925
rect 49651 8792 51074 8820
rect 49651 8789 49663 8792
rect 49605 8783 49663 8789
rect 1104 8730 58880 8752
rect 1104 8678 19574 8730
rect 19626 8678 19638 8730
rect 19690 8678 19702 8730
rect 19754 8678 19766 8730
rect 19818 8678 19830 8730
rect 19882 8678 50294 8730
rect 50346 8678 50358 8730
rect 50410 8678 50422 8730
rect 50474 8678 50486 8730
rect 50538 8678 50550 8730
rect 50602 8678 58880 8730
rect 1104 8656 58880 8678
rect 2225 8619 2283 8625
rect 2225 8585 2237 8619
rect 2271 8616 2283 8619
rect 2958 8616 2964 8628
rect 2271 8588 2964 8616
rect 2271 8585 2283 8588
rect 2225 8579 2283 8585
rect 1673 8483 1731 8489
rect 1673 8449 1685 8483
rect 1719 8480 1731 8483
rect 2240 8480 2268 8579
rect 2958 8576 2964 8588
rect 3016 8576 3022 8628
rect 4614 8616 4620 8628
rect 3436 8588 4620 8616
rect 1719 8452 2268 8480
rect 2869 8483 2927 8489
rect 1719 8449 1731 8452
rect 1673 8443 1731 8449
rect 2869 8449 2881 8483
rect 2915 8480 2927 8483
rect 3436 8480 3464 8588
rect 4614 8576 4620 8588
rect 4672 8576 4678 8628
rect 8570 8616 8576 8628
rect 8531 8588 8576 8616
rect 8570 8576 8576 8588
rect 8628 8576 8634 8628
rect 17681 8619 17739 8625
rect 17681 8585 17693 8619
rect 17727 8616 17739 8619
rect 17770 8616 17776 8628
rect 17727 8588 17776 8616
rect 17727 8585 17739 8588
rect 17681 8579 17739 8585
rect 17770 8576 17776 8588
rect 17828 8576 17834 8628
rect 18230 8576 18236 8628
rect 18288 8616 18294 8628
rect 18325 8619 18383 8625
rect 18325 8616 18337 8619
rect 18288 8588 18337 8616
rect 18288 8576 18294 8588
rect 18325 8585 18337 8588
rect 18371 8585 18383 8619
rect 18325 8579 18383 8585
rect 21085 8619 21143 8625
rect 21085 8585 21097 8619
rect 21131 8616 21143 8619
rect 21174 8616 21180 8628
rect 21131 8588 21180 8616
rect 21131 8585 21143 8588
rect 21085 8579 21143 8585
rect 21174 8576 21180 8588
rect 21232 8616 21238 8628
rect 22002 8616 22008 8628
rect 21232 8588 22008 8616
rect 21232 8576 21238 8588
rect 22002 8576 22008 8588
rect 22060 8576 22066 8628
rect 28258 8576 28264 8628
rect 28316 8616 28322 8628
rect 28316 8588 29132 8616
rect 28316 8576 28322 8588
rect 3896 8520 4660 8548
rect 3896 8492 3924 8520
rect 3878 8480 3884 8492
rect 2915 8452 3464 8480
rect 3528 8452 3884 8480
rect 2915 8449 2927 8452
rect 2869 8443 2927 8449
rect 3528 8421 3556 8452
rect 3878 8440 3884 8452
rect 3936 8440 3942 8492
rect 4433 8483 4491 8489
rect 4433 8449 4445 8483
rect 4479 8480 4491 8483
rect 4522 8480 4528 8492
rect 4479 8452 4528 8480
rect 4479 8449 4491 8452
rect 4433 8443 4491 8449
rect 4522 8440 4528 8452
rect 4580 8440 4586 8492
rect 4632 8489 4660 8520
rect 17126 8508 17132 8560
rect 17184 8548 17190 8560
rect 22922 8548 22928 8560
rect 17184 8520 22928 8548
rect 17184 8508 17190 8520
rect 22922 8508 22928 8520
rect 22980 8508 22986 8560
rect 25038 8548 25044 8560
rect 24999 8520 25044 8548
rect 25038 8508 25044 8520
rect 25096 8548 25102 8560
rect 28166 8548 28172 8560
rect 25096 8520 28172 8548
rect 25096 8508 25102 8520
rect 28166 8508 28172 8520
rect 28224 8548 28230 8560
rect 28629 8551 28687 8557
rect 28629 8548 28641 8551
rect 28224 8520 28641 8548
rect 28224 8508 28230 8520
rect 28629 8517 28641 8520
rect 28675 8517 28687 8551
rect 28629 8511 28687 8517
rect 28721 8551 28779 8557
rect 28721 8517 28733 8551
rect 28767 8548 28779 8551
rect 28994 8548 29000 8560
rect 28767 8520 29000 8548
rect 28767 8517 28779 8520
rect 28721 8511 28779 8517
rect 28994 8508 29000 8520
rect 29052 8508 29058 8560
rect 29104 8548 29132 8588
rect 29362 8576 29368 8628
rect 29420 8616 29426 8628
rect 29457 8619 29515 8625
rect 29457 8616 29469 8619
rect 29420 8588 29469 8616
rect 29420 8576 29426 8588
rect 29457 8585 29469 8588
rect 29503 8585 29515 8619
rect 29457 8579 29515 8585
rect 30374 8576 30380 8628
rect 30432 8616 30438 8628
rect 31389 8619 31447 8625
rect 31389 8616 31401 8619
rect 30432 8588 31401 8616
rect 30432 8576 30438 8588
rect 31389 8585 31401 8588
rect 31435 8585 31447 8619
rect 31389 8579 31447 8585
rect 34793 8619 34851 8625
rect 34793 8585 34805 8619
rect 34839 8616 34851 8619
rect 36538 8616 36544 8628
rect 34839 8588 36544 8616
rect 34839 8585 34851 8588
rect 34793 8579 34851 8585
rect 36538 8576 36544 8588
rect 36596 8576 36602 8628
rect 39114 8616 39120 8628
rect 39075 8588 39120 8616
rect 39114 8576 39120 8588
rect 39172 8576 39178 8628
rect 48314 8576 48320 8628
rect 48372 8616 48378 8628
rect 48593 8619 48651 8625
rect 48593 8616 48605 8619
rect 48372 8588 48605 8616
rect 48372 8576 48378 8588
rect 48593 8585 48605 8588
rect 48639 8585 48651 8619
rect 51534 8616 51540 8628
rect 51495 8588 51540 8616
rect 48593 8579 48651 8585
rect 51534 8576 51540 8588
rect 51592 8576 51598 8628
rect 53837 8619 53895 8625
rect 53837 8585 53849 8619
rect 53883 8616 53895 8619
rect 56226 8616 56232 8628
rect 53883 8588 56232 8616
rect 53883 8585 53895 8588
rect 53837 8579 53895 8585
rect 56226 8576 56232 8588
rect 56284 8576 56290 8628
rect 29730 8548 29736 8560
rect 29104 8520 29736 8548
rect 29730 8508 29736 8520
rect 29788 8508 29794 8560
rect 36262 8548 36268 8560
rect 36223 8520 36268 8548
rect 36262 8508 36268 8520
rect 36320 8508 36326 8560
rect 40221 8551 40279 8557
rect 40221 8548 40233 8551
rect 39592 8520 40233 8548
rect 4617 8483 4675 8489
rect 4617 8449 4629 8483
rect 4663 8449 4675 8483
rect 6546 8480 6552 8492
rect 6507 8452 6552 8480
rect 4617 8443 4675 8449
rect 6546 8440 6552 8452
rect 6604 8440 6610 8492
rect 6825 8483 6883 8489
rect 6825 8449 6837 8483
rect 6871 8449 6883 8483
rect 7006 8480 7012 8492
rect 6967 8452 7012 8480
rect 6825 8443 6883 8449
rect 2685 8415 2743 8421
rect 2685 8381 2697 8415
rect 2731 8412 2743 8415
rect 3513 8415 3571 8421
rect 3513 8412 3525 8415
rect 2731 8384 3525 8412
rect 2731 8381 2743 8384
rect 2685 8375 2743 8381
rect 3513 8381 3525 8384
rect 3559 8381 3571 8415
rect 3970 8412 3976 8424
rect 3883 8384 3976 8412
rect 3513 8375 3571 8381
rect 3970 8372 3976 8384
rect 4028 8412 4034 8424
rect 6365 8415 6423 8421
rect 6365 8412 6377 8415
rect 4028 8384 6377 8412
rect 4028 8372 4034 8384
rect 6365 8381 6377 8384
rect 6411 8381 6423 8415
rect 6840 8412 6868 8443
rect 7006 8440 7012 8452
rect 7064 8440 7070 8492
rect 15562 8440 15568 8492
rect 15620 8480 15626 8492
rect 19153 8483 19211 8489
rect 19153 8480 19165 8483
rect 15620 8452 19165 8480
rect 15620 8440 15626 8452
rect 19153 8449 19165 8452
rect 19199 8480 19211 8483
rect 19426 8480 19432 8492
rect 19199 8452 19432 8480
rect 19199 8449 19211 8452
rect 19153 8443 19211 8449
rect 19426 8440 19432 8452
rect 19484 8440 19490 8492
rect 24762 8480 24768 8492
rect 24504 8452 24768 8480
rect 6914 8412 6920 8424
rect 6827 8384 6920 8412
rect 6365 8375 6423 8381
rect 6914 8372 6920 8384
rect 6972 8412 6978 8424
rect 7650 8412 7656 8424
rect 6972 8384 7656 8412
rect 6972 8372 6978 8384
rect 7650 8372 7656 8384
rect 7708 8372 7714 8424
rect 19444 8412 19472 8440
rect 24504 8421 24532 8452
rect 24762 8440 24768 8452
rect 24820 8480 24826 8492
rect 24820 8452 25268 8480
rect 24820 8440 24826 8452
rect 24489 8415 24547 8421
rect 24489 8412 24501 8415
rect 19444 8384 24501 8412
rect 24489 8381 24501 8384
rect 24535 8381 24547 8415
rect 24489 8375 24547 8381
rect 25133 8415 25191 8421
rect 25133 8381 25145 8415
rect 25179 8381 25191 8415
rect 25240 8412 25268 8452
rect 25314 8440 25320 8492
rect 25372 8480 25378 8492
rect 25409 8483 25467 8489
rect 25409 8480 25421 8483
rect 25372 8452 25421 8480
rect 25372 8440 25378 8452
rect 25409 8449 25421 8452
rect 25455 8449 25467 8483
rect 25409 8443 25467 8449
rect 28445 8483 28503 8489
rect 28445 8449 28457 8483
rect 28491 8480 28503 8483
rect 28534 8480 28540 8492
rect 28491 8452 28540 8480
rect 28491 8449 28503 8452
rect 28445 8443 28503 8449
rect 28534 8440 28540 8452
rect 28592 8440 28598 8492
rect 28810 8480 28816 8492
rect 28771 8452 28816 8480
rect 28810 8440 28816 8452
rect 28868 8440 28874 8492
rect 30282 8480 30288 8492
rect 28920 8452 30288 8480
rect 25501 8415 25559 8421
rect 25501 8412 25513 8415
rect 25240 8384 25513 8412
rect 25133 8375 25191 8381
rect 25501 8381 25513 8384
rect 25547 8381 25559 8415
rect 25501 8375 25559 8381
rect 1486 8344 1492 8356
rect 1447 8316 1492 8344
rect 1486 8304 1492 8316
rect 1544 8304 1550 8356
rect 3050 8344 3056 8356
rect 3011 8316 3056 8344
rect 3050 8304 3056 8316
rect 3108 8304 3114 8356
rect 3697 8347 3755 8353
rect 3697 8313 3709 8347
rect 3743 8344 3755 8347
rect 4062 8344 4068 8356
rect 3743 8316 4068 8344
rect 3743 8313 3755 8316
rect 3697 8307 3755 8313
rect 4062 8304 4068 8316
rect 4120 8304 4126 8356
rect 4433 8347 4491 8353
rect 4433 8344 4445 8347
rect 4172 8316 4445 8344
rect 3602 8236 3608 8288
rect 3660 8276 3666 8288
rect 3878 8276 3884 8288
rect 3660 8248 3884 8276
rect 3660 8236 3666 8248
rect 3878 8236 3884 8248
rect 3936 8276 3942 8288
rect 4172 8276 4200 8316
rect 4433 8313 4445 8316
rect 4479 8313 4491 8347
rect 4433 8307 4491 8313
rect 23382 8304 23388 8356
rect 23440 8344 23446 8356
rect 25148 8344 25176 8375
rect 25590 8372 25596 8424
rect 25648 8412 25654 8424
rect 28920 8412 28948 8452
rect 30282 8440 30288 8452
rect 30340 8440 30346 8492
rect 34422 8480 34428 8492
rect 34383 8452 34428 8480
rect 34422 8440 34428 8452
rect 34480 8440 34486 8492
rect 34606 8480 34612 8492
rect 34567 8452 34612 8480
rect 34606 8440 34612 8452
rect 34664 8440 34670 8492
rect 37550 8480 37556 8492
rect 37511 8452 37556 8480
rect 37550 8440 37556 8452
rect 37608 8440 37614 8492
rect 37918 8480 37924 8492
rect 37879 8452 37924 8480
rect 37918 8440 37924 8452
rect 37976 8440 37982 8492
rect 38102 8440 38108 8492
rect 38160 8480 38166 8492
rect 39592 8489 39620 8520
rect 40221 8517 40233 8520
rect 40267 8517 40279 8551
rect 40221 8511 40279 8517
rect 52546 8508 52552 8560
rect 52604 8548 52610 8560
rect 52604 8520 53052 8548
rect 52604 8508 52610 8520
rect 39301 8483 39359 8489
rect 39301 8480 39313 8483
rect 38160 8452 39313 8480
rect 38160 8440 38166 8452
rect 39301 8449 39313 8452
rect 39347 8449 39359 8483
rect 39301 8443 39359 8449
rect 39393 8483 39451 8489
rect 39393 8449 39405 8483
rect 39439 8449 39451 8483
rect 39393 8443 39451 8449
rect 39577 8483 39635 8489
rect 39577 8449 39589 8483
rect 39623 8449 39635 8483
rect 40126 8480 40132 8492
rect 40087 8452 40132 8480
rect 39577 8443 39635 8449
rect 25648 8384 28948 8412
rect 38565 8415 38623 8421
rect 25648 8372 25654 8384
rect 38565 8381 38577 8415
rect 38611 8412 38623 8415
rect 39114 8412 39120 8424
rect 38611 8384 39120 8412
rect 38611 8381 38623 8384
rect 38565 8375 38623 8381
rect 39114 8372 39120 8384
rect 39172 8412 39178 8424
rect 39408 8412 39436 8443
rect 40126 8440 40132 8452
rect 40184 8440 40190 8492
rect 40313 8483 40371 8489
rect 40313 8449 40325 8483
rect 40359 8480 40371 8483
rect 41046 8480 41052 8492
rect 40359 8452 41052 8480
rect 40359 8449 40371 8452
rect 40313 8443 40371 8449
rect 41046 8440 41052 8452
rect 41104 8440 41110 8492
rect 42334 8440 42340 8492
rect 42392 8480 42398 8492
rect 42613 8483 42671 8489
rect 42613 8480 42625 8483
rect 42392 8452 42625 8480
rect 42392 8440 42398 8452
rect 42613 8449 42625 8452
rect 42659 8449 42671 8483
rect 46014 8480 46020 8492
rect 45975 8452 46020 8480
rect 42613 8443 42671 8449
rect 46014 8440 46020 8452
rect 46072 8440 46078 8492
rect 48590 8483 48648 8489
rect 48590 8449 48602 8483
rect 48636 8480 48648 8483
rect 48682 8480 48688 8492
rect 48636 8452 48688 8480
rect 48636 8449 48648 8452
rect 48590 8443 48648 8449
rect 48682 8440 48688 8452
rect 48740 8440 48746 8492
rect 48958 8480 48964 8492
rect 48919 8452 48964 8480
rect 48958 8440 48964 8452
rect 49016 8440 49022 8492
rect 49053 8483 49111 8489
rect 49053 8449 49065 8483
rect 49099 8480 49111 8483
rect 49142 8480 49148 8492
rect 49099 8452 49148 8480
rect 49099 8449 49111 8452
rect 49053 8443 49111 8449
rect 49142 8440 49148 8452
rect 49200 8440 49206 8492
rect 51442 8480 51448 8492
rect 51403 8452 51448 8480
rect 51442 8440 51448 8452
rect 51500 8440 51506 8492
rect 51629 8483 51687 8489
rect 51629 8449 51641 8483
rect 51675 8480 51687 8483
rect 51810 8480 51816 8492
rect 51675 8452 51816 8480
rect 51675 8449 51687 8452
rect 51629 8443 51687 8449
rect 51810 8440 51816 8452
rect 51868 8480 51874 8492
rect 52086 8480 52092 8492
rect 51868 8452 52092 8480
rect 51868 8440 51874 8452
rect 52086 8440 52092 8452
rect 52144 8440 52150 8492
rect 52822 8480 52828 8492
rect 52783 8452 52828 8480
rect 52822 8440 52828 8452
rect 52880 8440 52886 8492
rect 53024 8489 53052 8520
rect 53009 8483 53067 8489
rect 53009 8449 53021 8483
rect 53055 8449 53067 8483
rect 54478 8480 54484 8492
rect 54439 8452 54484 8480
rect 53009 8443 53067 8449
rect 54478 8440 54484 8452
rect 54536 8440 54542 8492
rect 57054 8480 57060 8492
rect 57015 8452 57060 8480
rect 57054 8440 57060 8452
rect 57112 8440 57118 8492
rect 42521 8415 42579 8421
rect 42521 8412 42533 8415
rect 39172 8384 42533 8412
rect 39172 8372 39178 8384
rect 42521 8381 42533 8384
rect 42567 8381 42579 8415
rect 45922 8412 45928 8424
rect 45883 8384 45928 8412
rect 42521 8375 42579 8381
rect 45922 8372 45928 8384
rect 45980 8372 45986 8424
rect 54570 8412 54576 8424
rect 54531 8384 54576 8412
rect 54570 8372 54576 8384
rect 54628 8372 54634 8424
rect 56134 8372 56140 8424
rect 56192 8412 56198 8424
rect 56229 8415 56287 8421
rect 56229 8412 56241 8415
rect 56192 8384 56241 8412
rect 56192 8372 56198 8384
rect 56229 8381 56241 8384
rect 56275 8381 56287 8415
rect 57146 8412 57152 8424
rect 57107 8384 57152 8412
rect 56229 8375 56287 8381
rect 57146 8372 57152 8384
rect 57204 8372 57210 8424
rect 27522 8344 27528 8356
rect 23440 8316 27528 8344
rect 23440 8304 23446 8316
rect 27522 8304 27528 8316
rect 27580 8304 27586 8356
rect 28997 8347 29055 8353
rect 28997 8313 29009 8347
rect 29043 8344 29055 8347
rect 31570 8344 31576 8356
rect 29043 8316 31576 8344
rect 29043 8313 29055 8316
rect 28997 8307 29055 8313
rect 31570 8304 31576 8316
rect 31628 8304 31634 8356
rect 39485 8347 39543 8353
rect 39485 8313 39497 8347
rect 39531 8344 39543 8347
rect 39666 8344 39672 8356
rect 39531 8316 39672 8344
rect 39531 8313 39543 8316
rect 39485 8307 39543 8313
rect 39666 8304 39672 8316
rect 39724 8304 39730 8356
rect 42981 8347 43039 8353
rect 42981 8313 42993 8347
rect 43027 8344 43039 8347
rect 45002 8344 45008 8356
rect 43027 8316 45008 8344
rect 43027 8313 43039 8316
rect 42981 8307 43039 8313
rect 45002 8304 45008 8316
rect 45060 8304 45066 8356
rect 46385 8347 46443 8353
rect 46385 8313 46397 8347
rect 46431 8344 46443 8347
rect 48314 8344 48320 8356
rect 46431 8316 48320 8344
rect 46431 8313 46443 8316
rect 46385 8307 46443 8313
rect 48314 8304 48320 8316
rect 48372 8304 48378 8356
rect 48406 8304 48412 8356
rect 48464 8344 48470 8356
rect 48464 8316 48509 8344
rect 48464 8304 48470 8316
rect 54662 8304 54668 8356
rect 54720 8344 54726 8356
rect 54849 8347 54907 8353
rect 54849 8344 54861 8347
rect 54720 8316 54861 8344
rect 54720 8304 54726 8316
rect 54849 8313 54861 8316
rect 54895 8313 54907 8347
rect 54849 8307 54907 8313
rect 3936 8248 4200 8276
rect 11793 8279 11851 8285
rect 3936 8236 3942 8248
rect 11793 8245 11805 8279
rect 11839 8276 11851 8279
rect 12434 8276 12440 8288
rect 11839 8248 12440 8276
rect 11839 8245 11851 8248
rect 11793 8239 11851 8245
rect 12434 8236 12440 8248
rect 12492 8236 12498 8288
rect 15010 8236 15016 8288
rect 15068 8276 15074 8288
rect 21358 8276 21364 8288
rect 15068 8248 21364 8276
rect 15068 8236 15074 8248
rect 21358 8236 21364 8248
rect 21416 8236 21422 8288
rect 25685 8279 25743 8285
rect 25685 8245 25697 8279
rect 25731 8276 25743 8279
rect 31662 8276 31668 8288
rect 25731 8248 31668 8276
rect 25731 8245 25743 8248
rect 25685 8239 25743 8245
rect 31662 8236 31668 8248
rect 31720 8236 31726 8288
rect 1104 8186 58880 8208
rect 1104 8134 4214 8186
rect 4266 8134 4278 8186
rect 4330 8134 4342 8186
rect 4394 8134 4406 8186
rect 4458 8134 4470 8186
rect 4522 8134 34934 8186
rect 34986 8134 34998 8186
rect 35050 8134 35062 8186
rect 35114 8134 35126 8186
rect 35178 8134 35190 8186
rect 35242 8134 58880 8186
rect 1104 8112 58880 8134
rect 3786 8072 3792 8084
rect 3747 8044 3792 8072
rect 3786 8032 3792 8044
rect 3844 8032 3850 8084
rect 6546 8032 6552 8084
rect 6604 8072 6610 8084
rect 6733 8075 6791 8081
rect 6733 8072 6745 8075
rect 6604 8044 6745 8072
rect 6604 8032 6610 8044
rect 6733 8041 6745 8044
rect 6779 8041 6791 8075
rect 7650 8072 7656 8084
rect 7611 8044 7656 8072
rect 6733 8035 6791 8041
rect 7650 8032 7656 8044
rect 7708 8032 7714 8084
rect 10870 8072 10876 8084
rect 10831 8044 10876 8072
rect 10870 8032 10876 8044
rect 10928 8032 10934 8084
rect 26510 8032 26516 8084
rect 26568 8072 26574 8084
rect 28258 8072 28264 8084
rect 26568 8044 28264 8072
rect 26568 8032 26574 8044
rect 28258 8032 28264 8044
rect 28316 8032 28322 8084
rect 28813 8075 28871 8081
rect 28813 8041 28825 8075
rect 28859 8072 28871 8075
rect 35618 8072 35624 8084
rect 28859 8044 35624 8072
rect 28859 8041 28871 8044
rect 28813 8035 28871 8041
rect 35618 8032 35624 8044
rect 35676 8072 35682 8084
rect 35713 8075 35771 8081
rect 35713 8072 35725 8075
rect 35676 8044 35725 8072
rect 35676 8032 35682 8044
rect 35713 8041 35725 8044
rect 35759 8041 35771 8075
rect 35713 8035 35771 8041
rect 3970 8004 3976 8016
rect 3931 7976 3976 8004
rect 3970 7964 3976 7976
rect 4028 7964 4034 8016
rect 6917 8007 6975 8013
rect 6917 7973 6929 8007
rect 6963 8004 6975 8007
rect 7837 8007 7895 8013
rect 7837 8004 7849 8007
rect 6963 7976 7144 8004
rect 6963 7973 6975 7976
rect 6917 7967 6975 7973
rect 7116 7868 7144 7976
rect 7208 7976 7849 8004
rect 7208 7945 7236 7976
rect 7837 7973 7849 7976
rect 7883 8004 7895 8007
rect 10321 8007 10379 8013
rect 10321 8004 10333 8007
rect 7883 7976 10333 8004
rect 7883 7973 7895 7976
rect 7837 7967 7895 7973
rect 10321 7973 10333 7976
rect 10367 7973 10379 8007
rect 10321 7967 10379 7973
rect 27801 8007 27859 8013
rect 27801 7973 27813 8007
rect 27847 8004 27859 8007
rect 45649 8007 45707 8013
rect 27847 7976 30972 8004
rect 27847 7973 27859 7976
rect 27801 7967 27859 7973
rect 7193 7939 7251 7945
rect 7193 7905 7205 7939
rect 7239 7905 7251 7939
rect 10962 7936 10968 7948
rect 10923 7908 10968 7936
rect 7193 7899 7251 7905
rect 10962 7896 10968 7908
rect 11020 7896 11026 7948
rect 14093 7939 14151 7945
rect 14093 7936 14105 7939
rect 12406 7908 14105 7936
rect 10502 7871 10560 7877
rect 7116 7840 8156 7868
rect 4246 7800 4252 7812
rect 4207 7772 4252 7800
rect 4246 7760 4252 7772
rect 4304 7760 4310 7812
rect 8128 7809 8156 7840
rect 10502 7837 10514 7871
rect 10548 7868 10560 7871
rect 11422 7868 11428 7880
rect 10548 7840 11428 7868
rect 10548 7837 10560 7840
rect 10502 7831 10560 7837
rect 11422 7828 11428 7840
rect 11480 7828 11486 7880
rect 11606 7828 11612 7880
rect 11664 7868 11670 7880
rect 12069 7871 12127 7877
rect 12069 7868 12081 7871
rect 11664 7840 12081 7868
rect 11664 7828 11670 7840
rect 12069 7837 12081 7840
rect 12115 7837 12127 7871
rect 12069 7831 12127 7837
rect 8113 7803 8171 7809
rect 8113 7769 8125 7803
rect 8159 7800 8171 7803
rect 9582 7800 9588 7812
rect 8159 7772 9588 7800
rect 8159 7769 8171 7772
rect 8113 7763 8171 7769
rect 9582 7760 9588 7772
rect 9640 7760 9646 7812
rect 10410 7760 10416 7812
rect 10468 7800 10474 7812
rect 12406 7800 12434 7908
rect 14093 7905 14105 7908
rect 14139 7905 14151 7939
rect 14093 7899 14151 7905
rect 17313 7939 17371 7945
rect 17313 7905 17325 7939
rect 17359 7936 17371 7939
rect 17402 7936 17408 7948
rect 17359 7908 17408 7936
rect 17359 7905 17371 7908
rect 17313 7899 17371 7905
rect 17402 7896 17408 7908
rect 17460 7936 17466 7948
rect 17770 7936 17776 7948
rect 17460 7908 17776 7936
rect 17460 7896 17466 7908
rect 17770 7896 17776 7908
rect 17828 7896 17834 7948
rect 20162 7936 20168 7948
rect 20123 7908 20168 7936
rect 20162 7896 20168 7908
rect 20220 7896 20226 7948
rect 21358 7936 21364 7948
rect 21319 7908 21364 7936
rect 21358 7896 21364 7908
rect 21416 7896 21422 7948
rect 22370 7936 22376 7948
rect 22331 7908 22376 7936
rect 22370 7896 22376 7908
rect 22428 7896 22434 7948
rect 23842 7936 23848 7948
rect 22664 7908 23848 7936
rect 14458 7868 14464 7880
rect 14419 7840 14464 7868
rect 14458 7828 14464 7840
rect 14516 7828 14522 7880
rect 14918 7868 14924 7880
rect 14831 7840 14924 7868
rect 14918 7828 14924 7840
rect 14976 7868 14982 7880
rect 16393 7871 16451 7877
rect 16393 7868 16405 7871
rect 14976 7840 16405 7868
rect 14976 7828 14982 7840
rect 16393 7837 16405 7840
rect 16439 7837 16451 7871
rect 16393 7831 16451 7837
rect 17221 7871 17279 7877
rect 17221 7837 17233 7871
rect 17267 7868 17279 7871
rect 18141 7871 18199 7877
rect 17267 7840 18092 7868
rect 17267 7837 17279 7840
rect 17221 7831 17279 7837
rect 10468 7772 12434 7800
rect 10468 7760 10474 7772
rect 18064 7744 18092 7840
rect 18141 7837 18153 7871
rect 18187 7868 18199 7871
rect 18230 7868 18236 7880
rect 18187 7840 18236 7868
rect 18187 7837 18199 7840
rect 18141 7831 18199 7837
rect 18230 7828 18236 7840
rect 18288 7828 18294 7880
rect 20254 7868 20260 7880
rect 20167 7840 20260 7868
rect 20254 7828 20260 7840
rect 20312 7868 20318 7880
rect 21174 7868 21180 7880
rect 20312 7840 20668 7868
rect 21135 7840 21180 7868
rect 20312 7828 20318 7840
rect 18248 7800 18276 7828
rect 20640 7812 20668 7840
rect 21174 7828 21180 7840
rect 21232 7828 21238 7880
rect 22664 7877 22692 7908
rect 23842 7896 23848 7908
rect 23900 7896 23906 7948
rect 28810 7936 28816 7948
rect 27356 7908 28816 7936
rect 27356 7880 27384 7908
rect 22649 7871 22707 7877
rect 22649 7868 22661 7871
rect 22066 7840 22661 7868
rect 18248 7772 20116 7800
rect 10502 7732 10508 7744
rect 10463 7704 10508 7732
rect 10502 7692 10508 7704
rect 10560 7692 10566 7744
rect 11514 7732 11520 7744
rect 11475 7704 11520 7732
rect 11514 7692 11520 7704
rect 11572 7692 11578 7744
rect 18046 7732 18052 7744
rect 18007 7704 18052 7732
rect 18046 7692 18052 7704
rect 18104 7692 18110 7744
rect 19889 7735 19947 7741
rect 19889 7701 19901 7735
rect 19935 7732 19947 7735
rect 19978 7732 19984 7744
rect 19935 7704 19984 7732
rect 19935 7701 19947 7704
rect 19889 7695 19947 7701
rect 19978 7692 19984 7704
rect 20036 7692 20042 7744
rect 20088 7732 20116 7772
rect 20622 7760 20628 7812
rect 20680 7800 20686 7812
rect 22066 7800 22094 7840
rect 22649 7837 22661 7840
rect 22695 7837 22707 7871
rect 27338 7868 27344 7880
rect 27299 7840 27344 7868
rect 22649 7831 22707 7837
rect 27338 7828 27344 7840
rect 27396 7828 27402 7880
rect 27617 7871 27675 7877
rect 27617 7837 27629 7871
rect 27663 7868 27675 7871
rect 27798 7868 27804 7880
rect 27663 7840 27804 7868
rect 27663 7837 27675 7840
rect 27617 7831 27675 7837
rect 27798 7828 27804 7840
rect 27856 7828 27862 7880
rect 28258 7868 28264 7880
rect 28219 7840 28264 7868
rect 28258 7828 28264 7840
rect 28316 7828 28322 7880
rect 28460 7877 28488 7908
rect 28810 7896 28816 7908
rect 28868 7896 28874 7948
rect 30193 7939 30251 7945
rect 30193 7905 30205 7939
rect 30239 7936 30251 7939
rect 30374 7936 30380 7948
rect 30239 7908 30380 7936
rect 30239 7905 30251 7908
rect 30193 7899 30251 7905
rect 30374 7896 30380 7908
rect 30432 7936 30438 7948
rect 30432 7908 30788 7936
rect 30432 7896 30438 7908
rect 28445 7871 28503 7877
rect 28445 7837 28457 7871
rect 28491 7837 28503 7871
rect 28445 7831 28503 7837
rect 28629 7871 28687 7877
rect 28629 7837 28641 7871
rect 28675 7837 28687 7871
rect 28629 7831 28687 7837
rect 20680 7772 22094 7800
rect 23293 7803 23351 7809
rect 20680 7760 20686 7772
rect 23293 7769 23305 7803
rect 23339 7800 23351 7803
rect 24210 7800 24216 7812
rect 23339 7772 24216 7800
rect 23339 7769 23351 7772
rect 23293 7763 23351 7769
rect 24210 7760 24216 7772
rect 24268 7760 24274 7812
rect 27433 7803 27491 7809
rect 27433 7769 27445 7803
rect 27479 7800 27491 7803
rect 28534 7800 28540 7812
rect 27479 7772 28540 7800
rect 27479 7769 27491 7772
rect 27433 7763 27491 7769
rect 28534 7760 28540 7772
rect 28592 7760 28598 7812
rect 23566 7732 23572 7744
rect 20088 7704 23572 7732
rect 23566 7692 23572 7704
rect 23624 7692 23630 7744
rect 23842 7732 23848 7744
rect 23755 7704 23848 7732
rect 23842 7692 23848 7704
rect 23900 7732 23906 7744
rect 27338 7732 27344 7744
rect 23900 7704 27344 7732
rect 23900 7692 23906 7704
rect 27338 7692 27344 7704
rect 27396 7692 27402 7744
rect 27982 7692 27988 7744
rect 28040 7732 28046 7744
rect 28644 7732 28672 7831
rect 29914 7828 29920 7880
rect 29972 7868 29978 7880
rect 30760 7877 30788 7908
rect 30944 7877 30972 7976
rect 45649 7973 45661 8007
rect 45695 8004 45707 8007
rect 45830 8004 45836 8016
rect 45695 7976 45836 8004
rect 45695 7973 45707 7976
rect 45649 7967 45707 7973
rect 45830 7964 45836 7976
rect 45888 7964 45894 8016
rect 48869 8007 48927 8013
rect 48869 7973 48881 8007
rect 48915 8004 48927 8007
rect 49142 8004 49148 8016
rect 48915 7976 49148 8004
rect 48915 7973 48927 7976
rect 48869 7967 48927 7973
rect 49142 7964 49148 7976
rect 49200 7964 49206 8016
rect 52086 8004 52092 8016
rect 52047 7976 52092 8004
rect 52086 7964 52092 7976
rect 52144 7964 52150 8016
rect 31570 7936 31576 7948
rect 31531 7908 31576 7936
rect 31570 7896 31576 7908
rect 31628 7896 31634 7948
rect 32122 7936 32128 7948
rect 32083 7908 32128 7936
rect 32122 7896 32128 7908
rect 32180 7896 32186 7948
rect 33134 7896 33140 7948
rect 33192 7936 33198 7948
rect 34701 7939 34759 7945
rect 34701 7936 34713 7939
rect 33192 7908 34713 7936
rect 33192 7896 33198 7908
rect 30653 7871 30711 7877
rect 30653 7868 30665 7871
rect 29972 7840 30665 7868
rect 29972 7828 29978 7840
rect 30653 7837 30665 7840
rect 30699 7837 30711 7871
rect 30653 7831 30711 7837
rect 30745 7871 30803 7877
rect 30745 7837 30757 7871
rect 30791 7837 30803 7871
rect 30745 7831 30803 7837
rect 30929 7871 30987 7877
rect 30929 7837 30941 7871
rect 30975 7837 30987 7871
rect 31941 7871 31999 7877
rect 31941 7868 31953 7871
rect 30929 7831 30987 7837
rect 31036 7840 31953 7868
rect 30760 7800 30788 7831
rect 31036 7800 31064 7840
rect 31941 7837 31953 7840
rect 31987 7837 31999 7871
rect 33410 7868 33416 7880
rect 33323 7840 33416 7868
rect 31941 7831 31999 7837
rect 33410 7828 33416 7840
rect 33468 7868 33474 7880
rect 34072 7877 34100 7908
rect 34701 7905 34713 7908
rect 34747 7905 34759 7939
rect 34701 7899 34759 7905
rect 38654 7896 38660 7948
rect 38712 7936 38718 7948
rect 39850 7936 39856 7948
rect 38712 7908 39856 7936
rect 38712 7896 38718 7908
rect 33873 7871 33931 7877
rect 33873 7868 33885 7871
rect 33468 7840 33885 7868
rect 33468 7828 33474 7840
rect 33873 7837 33885 7840
rect 33919 7837 33931 7871
rect 33873 7831 33931 7837
rect 34057 7871 34115 7877
rect 34057 7837 34069 7871
rect 34103 7837 34115 7871
rect 35710 7868 35716 7880
rect 35671 7840 35716 7868
rect 34057 7831 34115 7837
rect 35710 7828 35716 7840
rect 35768 7828 35774 7880
rect 35894 7868 35900 7880
rect 35855 7840 35900 7868
rect 35894 7828 35900 7840
rect 35952 7828 35958 7880
rect 39114 7868 39120 7880
rect 39075 7840 39120 7868
rect 39114 7828 39120 7840
rect 39172 7828 39178 7880
rect 39316 7877 39344 7908
rect 39850 7896 39856 7908
rect 39908 7896 39914 7948
rect 40957 7939 41015 7945
rect 40957 7905 40969 7939
rect 41003 7936 41015 7939
rect 41046 7936 41052 7948
rect 41003 7908 41052 7936
rect 41003 7905 41015 7908
rect 40957 7899 41015 7905
rect 41046 7896 41052 7908
rect 41104 7896 41110 7948
rect 41892 7908 42840 7936
rect 41892 7880 41920 7908
rect 39301 7871 39359 7877
rect 39301 7837 39313 7871
rect 39347 7837 39359 7871
rect 39301 7831 39359 7837
rect 39666 7828 39672 7880
rect 39724 7868 39730 7880
rect 39945 7871 40003 7877
rect 39945 7868 39957 7871
rect 39724 7840 39957 7868
rect 39724 7828 39730 7840
rect 39945 7837 39957 7840
rect 39991 7837 40003 7871
rect 39945 7831 40003 7837
rect 40129 7871 40187 7877
rect 40129 7837 40141 7871
rect 40175 7837 40187 7871
rect 40129 7831 40187 7837
rect 41693 7871 41751 7877
rect 41693 7837 41705 7871
rect 41739 7837 41751 7871
rect 41874 7868 41880 7880
rect 41835 7840 41880 7868
rect 41693 7831 41751 7837
rect 30760 7772 31064 7800
rect 31113 7803 31171 7809
rect 31113 7769 31125 7803
rect 31159 7800 31171 7803
rect 37734 7800 37740 7812
rect 31159 7772 37740 7800
rect 31159 7769 31171 7772
rect 31113 7763 31171 7769
rect 37734 7760 37740 7772
rect 37792 7760 37798 7812
rect 39209 7803 39267 7809
rect 39209 7769 39221 7803
rect 39255 7800 39267 7803
rect 40144 7800 40172 7831
rect 41708 7800 41736 7831
rect 41874 7828 41880 7840
rect 41932 7828 41938 7880
rect 42334 7868 42340 7880
rect 42295 7840 42340 7868
rect 42334 7828 42340 7840
rect 42392 7828 42398 7880
rect 42518 7868 42524 7880
rect 42479 7840 42524 7868
rect 42518 7828 42524 7840
rect 42576 7828 42582 7880
rect 42812 7877 42840 7908
rect 48314 7896 48320 7948
rect 48372 7936 48378 7948
rect 48409 7939 48467 7945
rect 48409 7936 48421 7939
rect 48372 7908 48421 7936
rect 48372 7896 48378 7908
rect 48409 7905 48421 7908
rect 48455 7905 48467 7939
rect 52822 7936 52828 7948
rect 48409 7899 48467 7905
rect 52288 7908 52828 7936
rect 42797 7871 42855 7877
rect 42797 7837 42809 7871
rect 42843 7837 42855 7871
rect 45554 7868 45560 7880
rect 45515 7840 45560 7868
rect 42797 7831 42855 7837
rect 45554 7828 45560 7840
rect 45612 7828 45618 7880
rect 45922 7868 45928 7880
rect 45883 7840 45928 7868
rect 45922 7828 45928 7840
rect 45980 7828 45986 7880
rect 46014 7828 46020 7880
rect 46072 7868 46078 7880
rect 46293 7871 46351 7877
rect 46293 7868 46305 7871
rect 46072 7840 46305 7868
rect 46072 7828 46078 7840
rect 46293 7837 46305 7840
rect 46339 7837 46351 7871
rect 46293 7831 46351 7837
rect 48501 7871 48559 7877
rect 48501 7837 48513 7871
rect 48547 7868 48559 7871
rect 48682 7868 48688 7880
rect 48547 7840 48688 7868
rect 48547 7837 48559 7840
rect 48501 7831 48559 7837
rect 48682 7828 48688 7840
rect 48740 7828 48746 7880
rect 51626 7868 51632 7880
rect 51587 7840 51632 7868
rect 51626 7828 51632 7840
rect 51684 7828 51690 7880
rect 51902 7868 51908 7880
rect 51863 7840 51908 7868
rect 51902 7828 51908 7840
rect 51960 7828 51966 7880
rect 52288 7877 52316 7908
rect 52822 7896 52828 7908
rect 52880 7896 52886 7948
rect 52273 7871 52331 7877
rect 52273 7837 52285 7871
rect 52319 7837 52331 7871
rect 52273 7831 52331 7837
rect 52365 7871 52423 7877
rect 52365 7837 52377 7871
rect 52411 7868 52423 7871
rect 52546 7868 52552 7880
rect 52411 7840 52552 7868
rect 52411 7837 52423 7840
rect 52365 7831 52423 7837
rect 52546 7828 52552 7840
rect 52604 7828 52610 7880
rect 58066 7868 58072 7880
rect 58027 7840 58072 7868
rect 58066 7828 58072 7840
rect 58124 7828 58130 7880
rect 42352 7800 42380 7828
rect 57514 7800 57520 7812
rect 39255 7772 40172 7800
rect 41386 7772 42380 7800
rect 57475 7772 57520 7800
rect 39255 7769 39267 7772
rect 39209 7763 39267 7769
rect 31938 7732 31944 7744
rect 28040 7704 28672 7732
rect 31899 7704 31944 7732
rect 28040 7692 28046 7704
rect 31938 7692 31944 7704
rect 31996 7692 32002 7744
rect 33962 7732 33968 7744
rect 33923 7704 33968 7732
rect 33962 7692 33968 7704
rect 34020 7692 34026 7744
rect 34882 7692 34888 7744
rect 34940 7732 34946 7744
rect 35802 7732 35808 7744
rect 34940 7704 35808 7732
rect 34940 7692 34946 7704
rect 35802 7692 35808 7704
rect 35860 7692 35866 7744
rect 36081 7735 36139 7741
rect 36081 7701 36093 7735
rect 36127 7732 36139 7735
rect 36446 7732 36452 7744
rect 36127 7704 36452 7732
rect 36127 7701 36139 7704
rect 36081 7695 36139 7701
rect 36446 7692 36452 7704
rect 36504 7692 36510 7744
rect 38930 7692 38936 7744
rect 38988 7732 38994 7744
rect 41386 7732 41414 7772
rect 57514 7760 57520 7772
rect 57572 7760 57578 7812
rect 38988 7704 41414 7732
rect 41785 7735 41843 7741
rect 38988 7692 38994 7704
rect 41785 7701 41797 7735
rect 41831 7732 41843 7735
rect 42610 7732 42616 7744
rect 41831 7704 42616 7732
rect 41831 7701 41843 7704
rect 41785 7695 41843 7701
rect 42610 7692 42616 7704
rect 42668 7692 42674 7744
rect 42981 7735 43039 7741
rect 42981 7701 42993 7735
rect 43027 7732 43039 7735
rect 45186 7732 45192 7744
rect 43027 7704 45192 7732
rect 43027 7701 43039 7704
rect 42981 7695 43039 7701
rect 45186 7692 45192 7704
rect 45244 7692 45250 7744
rect 1104 7642 58880 7664
rect 1104 7590 19574 7642
rect 19626 7590 19638 7642
rect 19690 7590 19702 7642
rect 19754 7590 19766 7642
rect 19818 7590 19830 7642
rect 19882 7590 50294 7642
rect 50346 7590 50358 7642
rect 50410 7590 50422 7642
rect 50474 7590 50486 7642
rect 50538 7590 50550 7642
rect 50602 7590 58880 7642
rect 1104 7568 58880 7590
rect 10781 7531 10839 7537
rect 10781 7497 10793 7531
rect 10827 7528 10839 7531
rect 10962 7528 10968 7540
rect 10827 7500 10968 7528
rect 10827 7497 10839 7500
rect 10781 7491 10839 7497
rect 10962 7488 10968 7500
rect 11020 7488 11026 7540
rect 11422 7488 11428 7540
rect 11480 7528 11486 7540
rect 11517 7531 11575 7537
rect 11517 7528 11529 7531
rect 11480 7500 11529 7528
rect 11480 7488 11486 7500
rect 11517 7497 11529 7500
rect 11563 7528 11575 7531
rect 12434 7528 12440 7540
rect 11563 7500 12440 7528
rect 11563 7497 11575 7500
rect 11517 7491 11575 7497
rect 12434 7488 12440 7500
rect 12492 7528 12498 7540
rect 13722 7528 13728 7540
rect 12492 7500 13728 7528
rect 12492 7488 12498 7500
rect 13722 7488 13728 7500
rect 13780 7488 13786 7540
rect 20622 7528 20628 7540
rect 20583 7500 20628 7528
rect 20622 7488 20628 7500
rect 20680 7488 20686 7540
rect 27798 7528 27804 7540
rect 27759 7500 27804 7528
rect 27798 7488 27804 7500
rect 27856 7488 27862 7540
rect 28166 7488 28172 7540
rect 28224 7528 28230 7540
rect 31478 7528 31484 7540
rect 28224 7500 28856 7528
rect 31439 7500 31484 7528
rect 28224 7488 28230 7500
rect 14277 7463 14335 7469
rect 14277 7429 14289 7463
rect 14323 7460 14335 7463
rect 14918 7460 14924 7472
rect 14323 7432 14924 7460
rect 14323 7429 14335 7432
rect 14277 7423 14335 7429
rect 14918 7420 14924 7432
rect 14976 7420 14982 7472
rect 22833 7463 22891 7469
rect 22833 7460 22845 7463
rect 22066 7432 22845 7460
rect 6730 7392 6736 7404
rect 6691 7364 6736 7392
rect 6730 7352 6736 7364
rect 6788 7352 6794 7404
rect 10410 7392 10416 7404
rect 10371 7364 10416 7392
rect 10410 7352 10416 7364
rect 10468 7352 10474 7404
rect 13081 7395 13139 7401
rect 13081 7361 13093 7395
rect 13127 7392 13139 7395
rect 14182 7392 14188 7404
rect 13127 7364 14188 7392
rect 13127 7361 13139 7364
rect 13081 7355 13139 7361
rect 14182 7352 14188 7364
rect 14240 7352 14246 7404
rect 16853 7395 16911 7401
rect 16853 7361 16865 7395
rect 16899 7392 16911 7395
rect 17402 7392 17408 7404
rect 16899 7364 17408 7392
rect 16899 7361 16911 7364
rect 16853 7355 16911 7361
rect 17402 7352 17408 7364
rect 17460 7352 17466 7404
rect 17678 7392 17684 7404
rect 17639 7364 17684 7392
rect 17678 7352 17684 7364
rect 17736 7392 17742 7404
rect 18693 7395 18751 7401
rect 17736 7364 18644 7392
rect 17736 7352 17742 7364
rect 4246 7284 4252 7336
rect 4304 7324 4310 7336
rect 6365 7327 6423 7333
rect 6365 7324 6377 7327
rect 4304 7296 6377 7324
rect 4304 7284 4310 7296
rect 6365 7293 6377 7296
rect 6411 7293 6423 7327
rect 6822 7324 6828 7336
rect 6783 7296 6828 7324
rect 6365 7287 6423 7293
rect 6822 7284 6828 7296
rect 6880 7284 6886 7336
rect 10505 7327 10563 7333
rect 10505 7293 10517 7327
rect 10551 7324 10563 7327
rect 11514 7324 11520 7336
rect 10551 7296 11520 7324
rect 10551 7293 10563 7296
rect 10505 7287 10563 7293
rect 11514 7284 11520 7296
rect 11572 7284 11578 7336
rect 13357 7327 13415 7333
rect 13357 7293 13369 7327
rect 13403 7324 13415 7327
rect 14366 7324 14372 7336
rect 13403 7296 14372 7324
rect 13403 7293 13415 7296
rect 13357 7287 13415 7293
rect 14366 7284 14372 7296
rect 14424 7284 14430 7336
rect 18616 7333 18644 7364
rect 18693 7361 18705 7395
rect 18739 7392 18751 7395
rect 22066 7392 22094 7432
rect 22833 7429 22845 7432
rect 22879 7429 22891 7463
rect 22833 7423 22891 7429
rect 23566 7420 23572 7472
rect 23624 7460 23630 7472
rect 23624 7432 24716 7460
rect 23624 7420 23630 7432
rect 18739 7364 22094 7392
rect 22741 7395 22799 7401
rect 18739 7361 18751 7364
rect 18693 7355 18751 7361
rect 22741 7361 22753 7395
rect 22787 7361 22799 7395
rect 22741 7355 22799 7361
rect 23017 7395 23075 7401
rect 23017 7361 23029 7395
rect 23063 7392 23075 7395
rect 23658 7392 23664 7404
rect 23063 7364 23664 7392
rect 23063 7361 23075 7364
rect 23017 7355 23075 7361
rect 17037 7327 17095 7333
rect 17037 7293 17049 7327
rect 17083 7324 17095 7327
rect 17865 7327 17923 7333
rect 17865 7324 17877 7327
rect 17083 7296 17877 7324
rect 17083 7293 17095 7296
rect 17037 7287 17095 7293
rect 17865 7293 17877 7296
rect 17911 7293 17923 7327
rect 17865 7287 17923 7293
rect 18601 7327 18659 7333
rect 18601 7293 18613 7327
rect 18647 7293 18659 7327
rect 18601 7287 18659 7293
rect 14001 7259 14059 7265
rect 14001 7225 14013 7259
rect 14047 7256 14059 7259
rect 14458 7256 14464 7268
rect 14047 7228 14464 7256
rect 14047 7225 14059 7228
rect 14001 7219 14059 7225
rect 14458 7216 14464 7228
rect 14516 7216 14522 7268
rect 17880 7256 17908 7287
rect 18046 7256 18052 7268
rect 17880 7228 18052 7256
rect 18046 7216 18052 7228
rect 18104 7256 18110 7268
rect 18708 7256 18736 7355
rect 22756 7324 22784 7355
rect 23658 7352 23664 7364
rect 23716 7352 23722 7404
rect 23750 7352 23756 7404
rect 23808 7392 23814 7404
rect 24688 7401 24716 7432
rect 26326 7420 26332 7472
rect 26384 7460 26390 7472
rect 26384 7432 27476 7460
rect 26384 7420 26390 7432
rect 24673 7395 24731 7401
rect 23808 7364 23853 7392
rect 23808 7352 23814 7364
rect 24673 7361 24685 7395
rect 24719 7392 24731 7395
rect 27154 7392 27160 7404
rect 24719 7364 26188 7392
rect 27115 7364 27160 7392
rect 24719 7361 24731 7364
rect 24673 7355 24731 7361
rect 23768 7324 23796 7352
rect 22756 7296 23796 7324
rect 18104 7228 18736 7256
rect 19061 7259 19119 7265
rect 18104 7216 18110 7228
rect 19061 7225 19073 7259
rect 19107 7256 19119 7259
rect 20254 7256 20260 7268
rect 19107 7228 20260 7256
rect 19107 7225 19119 7228
rect 19061 7219 19119 7225
rect 20254 7216 20260 7228
rect 20312 7216 20318 7268
rect 26160 7265 26188 7364
rect 27154 7352 27160 7364
rect 27212 7352 27218 7404
rect 27341 7395 27399 7401
rect 27341 7361 27353 7395
rect 27387 7361 27399 7395
rect 27448 7392 27476 7432
rect 28258 7420 28264 7472
rect 28316 7460 28322 7472
rect 28316 7432 28396 7460
rect 28316 7420 28322 7432
rect 27982 7392 27988 7404
rect 27448 7364 27988 7392
rect 27908 7362 27988 7364
rect 27341 7355 27399 7361
rect 27356 7324 27384 7355
rect 27982 7352 27988 7362
rect 28040 7352 28046 7404
rect 28077 7395 28135 7401
rect 28077 7361 28089 7395
rect 28123 7361 28135 7395
rect 28077 7355 28135 7361
rect 28092 7324 28120 7355
rect 28166 7352 28172 7404
rect 28224 7392 28230 7404
rect 28368 7401 28396 7432
rect 28828 7401 28856 7500
rect 31478 7488 31484 7500
rect 31536 7488 31542 7540
rect 31662 7488 31668 7540
rect 31720 7528 31726 7540
rect 33965 7531 34023 7537
rect 31720 7500 31892 7528
rect 31720 7488 31726 7500
rect 28353 7395 28411 7401
rect 28224 7364 28269 7392
rect 28224 7352 28230 7364
rect 28353 7361 28365 7395
rect 28399 7361 28411 7395
rect 28353 7355 28411 7361
rect 28813 7395 28871 7401
rect 28813 7361 28825 7395
rect 28859 7361 28871 7395
rect 28994 7392 29000 7404
rect 28813 7355 28871 7361
rect 28966 7352 29000 7392
rect 29052 7392 29058 7404
rect 30653 7395 30711 7401
rect 29052 7364 29097 7392
rect 29052 7352 29058 7364
rect 30653 7361 30665 7395
rect 30699 7392 30711 7395
rect 31478 7392 31484 7404
rect 30699 7364 31484 7392
rect 30699 7361 30711 7364
rect 30653 7355 30711 7361
rect 28966 7324 28994 7352
rect 30558 7324 30564 7336
rect 27356 7296 28994 7324
rect 30519 7296 30564 7324
rect 30558 7284 30564 7296
rect 30616 7284 30622 7336
rect 26145 7259 26203 7265
rect 26145 7225 26157 7259
rect 26191 7256 26203 7259
rect 27338 7256 27344 7268
rect 26191 7228 27344 7256
rect 26191 7225 26203 7228
rect 26145 7219 26203 7225
rect 27338 7216 27344 7228
rect 27396 7216 27402 7268
rect 27430 7216 27436 7268
rect 27488 7256 27494 7268
rect 30668 7256 30696 7355
rect 31478 7352 31484 7364
rect 31536 7352 31542 7404
rect 31018 7256 31024 7268
rect 27488 7228 30696 7256
rect 30979 7228 31024 7256
rect 27488 7216 27494 7228
rect 31018 7216 31024 7228
rect 31076 7216 31082 7268
rect 31864 7256 31892 7500
rect 33965 7497 33977 7531
rect 34011 7528 34023 7531
rect 35526 7528 35532 7540
rect 34011 7500 35532 7528
rect 34011 7497 34023 7500
rect 33965 7491 34023 7497
rect 35526 7488 35532 7500
rect 35584 7488 35590 7540
rect 43530 7528 43536 7540
rect 35636 7500 43536 7528
rect 31938 7420 31944 7472
rect 31996 7460 32002 7472
rect 35636 7460 35664 7500
rect 43530 7488 43536 7500
rect 43588 7488 43594 7540
rect 46014 7528 46020 7540
rect 45975 7500 46020 7528
rect 46014 7488 46020 7500
rect 46072 7488 46078 7540
rect 58066 7528 58072 7540
rect 58027 7500 58072 7528
rect 58066 7488 58072 7500
rect 58124 7488 58130 7540
rect 31996 7432 35664 7460
rect 31996 7420 32002 7432
rect 35894 7420 35900 7472
rect 35952 7460 35958 7472
rect 36081 7463 36139 7469
rect 36081 7460 36093 7463
rect 35952 7432 36093 7460
rect 35952 7420 35958 7432
rect 36081 7429 36093 7432
rect 36127 7429 36139 7463
rect 36081 7423 36139 7429
rect 42518 7420 42524 7472
rect 42576 7460 42582 7472
rect 52181 7463 52239 7469
rect 42576 7432 42748 7460
rect 42576 7420 42582 7432
rect 32306 7352 32312 7404
rect 32364 7392 32370 7404
rect 33137 7395 33195 7401
rect 33137 7392 33149 7395
rect 32364 7364 33149 7392
rect 32364 7352 32370 7364
rect 33137 7361 33149 7364
rect 33183 7361 33195 7395
rect 33137 7355 33195 7361
rect 33962 7352 33968 7404
rect 34020 7392 34026 7404
rect 34701 7395 34759 7401
rect 34701 7392 34713 7395
rect 34020 7364 34713 7392
rect 34020 7352 34026 7364
rect 34701 7361 34713 7364
rect 34747 7361 34759 7395
rect 34882 7392 34888 7404
rect 34843 7364 34888 7392
rect 34701 7355 34759 7361
rect 34882 7352 34888 7364
rect 34940 7352 34946 7404
rect 35710 7392 35716 7404
rect 34992 7364 35716 7392
rect 33226 7324 33232 7336
rect 33187 7296 33232 7324
rect 33226 7284 33232 7296
rect 33284 7284 33290 7336
rect 34992 7324 35020 7364
rect 35710 7352 35716 7364
rect 35768 7352 35774 7404
rect 38657 7395 38715 7401
rect 38657 7361 38669 7395
rect 38703 7392 38715 7395
rect 38930 7392 38936 7404
rect 38703 7364 38936 7392
rect 38703 7361 38715 7364
rect 38657 7355 38715 7361
rect 38930 7352 38936 7364
rect 38988 7352 38994 7404
rect 42610 7392 42616 7404
rect 42571 7364 42616 7392
rect 42610 7352 42616 7364
rect 42668 7352 42674 7404
rect 42720 7378 42748 7432
rect 52181 7429 52193 7463
rect 52227 7460 52239 7463
rect 52822 7460 52828 7472
rect 52227 7432 52828 7460
rect 52227 7429 52239 7432
rect 52181 7423 52239 7429
rect 52822 7420 52828 7432
rect 52880 7420 52886 7472
rect 45002 7392 45008 7404
rect 44963 7364 45008 7392
rect 45002 7352 45008 7364
rect 45060 7352 45066 7404
rect 45186 7392 45192 7404
rect 45147 7364 45192 7392
rect 45186 7352 45192 7364
rect 45244 7352 45250 7404
rect 51626 7352 51632 7404
rect 51684 7352 51690 7404
rect 56226 7352 56232 7404
rect 56284 7392 56290 7404
rect 56965 7395 57023 7401
rect 56965 7392 56977 7395
rect 56284 7364 56977 7392
rect 56284 7352 56290 7364
rect 56965 7361 56977 7364
rect 57011 7361 57023 7395
rect 56965 7355 57023 7361
rect 35618 7324 35624 7336
rect 34624 7296 35020 7324
rect 35579 7296 35624 7324
rect 34624 7256 34652 7296
rect 35618 7284 35624 7296
rect 35676 7284 35682 7336
rect 39666 7324 39672 7336
rect 39627 7296 39672 7324
rect 39666 7284 39672 7296
rect 39724 7284 39730 7336
rect 43625 7327 43683 7333
rect 43625 7293 43637 7327
rect 43671 7324 43683 7327
rect 45462 7324 45468 7336
rect 43671 7296 45468 7324
rect 43671 7293 43683 7296
rect 43625 7287 43683 7293
rect 45462 7284 45468 7296
rect 45520 7284 45526 7336
rect 51353 7327 51411 7333
rect 51353 7293 51365 7327
rect 51399 7324 51411 7327
rect 51902 7324 51908 7336
rect 51399 7296 51908 7324
rect 51399 7293 51411 7296
rect 51353 7287 51411 7293
rect 51902 7284 51908 7296
rect 51960 7284 51966 7336
rect 57054 7324 57060 7336
rect 57015 7296 57060 7324
rect 57054 7284 57060 7296
rect 57112 7284 57118 7336
rect 57330 7324 57336 7336
rect 57291 7296 57336 7324
rect 57330 7284 57336 7296
rect 57388 7284 57394 7336
rect 31864 7228 34652 7256
rect 34698 7216 34704 7268
rect 34756 7256 34762 7268
rect 35713 7259 35771 7265
rect 34756 7228 34801 7256
rect 34756 7216 34762 7228
rect 35713 7225 35725 7259
rect 35759 7225 35771 7259
rect 35713 7219 35771 7225
rect 12894 7188 12900 7200
rect 12855 7160 12900 7188
rect 12894 7148 12900 7160
rect 12952 7148 12958 7200
rect 13265 7191 13323 7197
rect 13265 7157 13277 7191
rect 13311 7188 13323 7191
rect 13817 7191 13875 7197
rect 13817 7188 13829 7191
rect 13311 7160 13829 7188
rect 13311 7157 13323 7160
rect 13265 7151 13323 7157
rect 13817 7157 13829 7160
rect 13863 7188 13875 7191
rect 14182 7188 14188 7200
rect 13863 7160 14188 7188
rect 13863 7157 13875 7160
rect 13817 7151 13875 7157
rect 14182 7148 14188 7160
rect 14240 7148 14246 7200
rect 14366 7148 14372 7200
rect 14424 7188 14430 7200
rect 16669 7191 16727 7197
rect 16669 7188 16681 7191
rect 14424 7160 16681 7188
rect 14424 7148 14430 7160
rect 16669 7157 16681 7160
rect 16715 7157 16727 7191
rect 16669 7151 16727 7157
rect 16850 7148 16856 7200
rect 16908 7188 16914 7200
rect 17497 7191 17555 7197
rect 17497 7188 17509 7191
rect 16908 7160 17509 7188
rect 16908 7148 16914 7160
rect 17497 7157 17509 7160
rect 17543 7157 17555 7191
rect 17497 7151 17555 7157
rect 23201 7191 23259 7197
rect 23201 7157 23213 7191
rect 23247 7188 23259 7191
rect 23290 7188 23296 7200
rect 23247 7160 23296 7188
rect 23247 7157 23259 7160
rect 23201 7151 23259 7157
rect 23290 7148 23296 7160
rect 23348 7148 23354 7200
rect 25222 7188 25228 7200
rect 25183 7160 25228 7188
rect 25222 7148 25228 7160
rect 25280 7148 25286 7200
rect 27249 7191 27307 7197
rect 27249 7157 27261 7191
rect 27295 7188 27307 7191
rect 27614 7188 27620 7200
rect 27295 7160 27620 7188
rect 27295 7157 27307 7160
rect 27249 7151 27307 7157
rect 27614 7148 27620 7160
rect 27672 7148 27678 7200
rect 28902 7188 28908 7200
rect 28863 7160 28908 7188
rect 28902 7148 28908 7160
rect 28960 7148 28966 7200
rect 32306 7188 32312 7200
rect 32267 7160 32312 7188
rect 32306 7148 32312 7160
rect 32364 7148 32370 7200
rect 35618 7148 35624 7200
rect 35676 7188 35682 7200
rect 35728 7188 35756 7219
rect 38470 7188 38476 7200
rect 35676 7160 35756 7188
rect 38431 7160 38476 7188
rect 35676 7148 35682 7160
rect 38470 7148 38476 7160
rect 38528 7148 38534 7200
rect 55766 7188 55772 7200
rect 55727 7160 55772 7188
rect 55766 7148 55772 7160
rect 55824 7148 55830 7200
rect 1104 7098 58880 7120
rect 1104 7046 4214 7098
rect 4266 7046 4278 7098
rect 4330 7046 4342 7098
rect 4394 7046 4406 7098
rect 4458 7046 4470 7098
rect 4522 7046 34934 7098
rect 34986 7046 34998 7098
rect 35050 7046 35062 7098
rect 35114 7046 35126 7098
rect 35178 7046 35190 7098
rect 35242 7046 58880 7098
rect 1104 7024 58880 7046
rect 9582 6984 9588 6996
rect 9543 6956 9588 6984
rect 9582 6944 9588 6956
rect 9640 6944 9646 6996
rect 10502 6944 10508 6996
rect 10560 6984 10566 6996
rect 10597 6987 10655 6993
rect 10597 6984 10609 6987
rect 10560 6956 10609 6984
rect 10560 6944 10566 6956
rect 10597 6953 10609 6956
rect 10643 6953 10655 6987
rect 10597 6947 10655 6953
rect 11333 6987 11391 6993
rect 11333 6953 11345 6987
rect 11379 6984 11391 6987
rect 11606 6984 11612 6996
rect 11379 6956 11612 6984
rect 11379 6953 11391 6956
rect 11333 6947 11391 6953
rect 11606 6944 11612 6956
rect 11664 6944 11670 6996
rect 17402 6984 17408 6996
rect 17363 6956 17408 6984
rect 17402 6944 17408 6956
rect 17460 6944 17466 6996
rect 18322 6944 18328 6996
rect 18380 6984 18386 6996
rect 26973 6987 27031 6993
rect 26973 6984 26985 6987
rect 18380 6956 26985 6984
rect 18380 6944 18386 6956
rect 26973 6953 26985 6956
rect 27019 6984 27031 6987
rect 27154 6984 27160 6996
rect 27019 6956 27160 6984
rect 27019 6953 27031 6956
rect 26973 6947 27031 6953
rect 27154 6944 27160 6956
rect 27212 6944 27218 6996
rect 27338 6944 27344 6996
rect 27396 6984 27402 6996
rect 33134 6984 33140 6996
rect 27396 6956 33140 6984
rect 27396 6944 27402 6956
rect 33134 6944 33140 6956
rect 33192 6944 33198 6996
rect 35894 6944 35900 6996
rect 35952 6984 35958 6996
rect 35989 6987 36047 6993
rect 35989 6984 36001 6987
rect 35952 6956 36001 6984
rect 35952 6944 35958 6956
rect 35989 6953 36001 6956
rect 36035 6953 36047 6987
rect 45554 6984 45560 6996
rect 45515 6956 45560 6984
rect 35989 6947 36047 6953
rect 45554 6944 45560 6956
rect 45612 6944 45618 6996
rect 48682 6984 48688 6996
rect 48643 6956 48688 6984
rect 48682 6944 48688 6956
rect 48740 6944 48746 6996
rect 51258 6944 51264 6996
rect 51316 6984 51322 6996
rect 51626 6984 51632 6996
rect 51316 6956 51632 6984
rect 51316 6944 51322 6956
rect 51626 6944 51632 6956
rect 51684 6944 51690 6996
rect 6730 6876 6736 6928
rect 6788 6916 6794 6928
rect 12894 6916 12900 6928
rect 6788 6888 12900 6916
rect 6788 6876 6794 6888
rect 12894 6876 12900 6888
rect 12952 6876 12958 6928
rect 14182 6916 14188 6928
rect 14143 6888 14188 6916
rect 14182 6876 14188 6888
rect 14240 6876 14246 6928
rect 19978 6916 19984 6928
rect 19939 6888 19984 6916
rect 19978 6876 19984 6888
rect 20036 6876 20042 6928
rect 38838 6916 38844 6928
rect 32324 6888 38844 6916
rect 32324 6860 32352 6888
rect 38838 6876 38844 6888
rect 38896 6916 38902 6928
rect 40126 6916 40132 6928
rect 38896 6888 39252 6916
rect 40087 6888 40132 6916
rect 38896 6876 38902 6888
rect 10042 6848 10048 6860
rect 10003 6820 10048 6848
rect 10042 6808 10048 6820
rect 10100 6808 10106 6860
rect 12802 6808 12808 6860
rect 12860 6848 12866 6860
rect 14366 6848 14372 6860
rect 12860 6820 13676 6848
rect 14327 6820 14372 6848
rect 12860 6808 12866 6820
rect 9953 6783 10011 6789
rect 9953 6749 9965 6783
rect 9999 6749 10011 6783
rect 9953 6743 10011 6749
rect 9968 6712 9996 6743
rect 10410 6740 10416 6792
rect 10468 6780 10474 6792
rect 10597 6783 10655 6789
rect 10597 6780 10609 6783
rect 10468 6752 10609 6780
rect 10468 6740 10474 6752
rect 10597 6749 10609 6752
rect 10643 6749 10655 6783
rect 10597 6743 10655 6749
rect 10781 6783 10839 6789
rect 10781 6749 10793 6783
rect 10827 6780 10839 6783
rect 11606 6780 11612 6792
rect 10827 6752 11612 6780
rect 10827 6749 10839 6752
rect 10781 6743 10839 6749
rect 11606 6740 11612 6752
rect 11664 6740 11670 6792
rect 12894 6740 12900 6792
rect 12952 6780 12958 6792
rect 13265 6783 13323 6789
rect 13265 6780 13277 6783
rect 12952 6752 13277 6780
rect 12952 6740 12958 6752
rect 13265 6749 13277 6752
rect 13311 6749 13323 6783
rect 13265 6743 13323 6749
rect 10134 6712 10140 6724
rect 9968 6684 10140 6712
rect 10134 6672 10140 6684
rect 10192 6712 10198 6724
rect 13081 6715 13139 6721
rect 13081 6712 13093 6715
rect 10192 6684 13093 6712
rect 10192 6672 10198 6684
rect 13081 6681 13093 6684
rect 13127 6681 13139 6715
rect 13081 6675 13139 6681
rect 13449 6715 13507 6721
rect 13449 6681 13461 6715
rect 13495 6681 13507 6715
rect 13648 6712 13676 6820
rect 14366 6808 14372 6820
rect 14424 6808 14430 6860
rect 16574 6848 16580 6860
rect 16535 6820 16580 6848
rect 16574 6808 16580 6820
rect 16632 6808 16638 6860
rect 16758 6808 16764 6860
rect 16816 6848 16822 6860
rect 19797 6851 19855 6857
rect 19797 6848 19809 6851
rect 16816 6820 19809 6848
rect 16816 6808 16822 6820
rect 19797 6817 19809 6820
rect 19843 6817 19855 6851
rect 20254 6848 20260 6860
rect 20215 6820 20260 6848
rect 19797 6811 19855 6817
rect 20254 6808 20260 6820
rect 20312 6808 20318 6860
rect 32306 6848 32312 6860
rect 27816 6820 32312 6848
rect 14093 6783 14151 6789
rect 14093 6749 14105 6783
rect 14139 6780 14151 6783
rect 14274 6780 14280 6792
rect 14139 6752 14280 6780
rect 14139 6749 14151 6752
rect 14093 6743 14151 6749
rect 14274 6740 14280 6752
rect 14332 6740 14338 6792
rect 16850 6740 16856 6792
rect 16908 6780 16914 6792
rect 16908 6752 16953 6780
rect 16908 6740 16914 6752
rect 24210 6740 24216 6792
rect 24268 6780 24274 6792
rect 24581 6783 24639 6789
rect 24581 6780 24593 6783
rect 24268 6752 24593 6780
rect 24268 6740 24274 6752
rect 24581 6749 24593 6752
rect 24627 6749 24639 6783
rect 25222 6780 25228 6792
rect 25183 6752 25228 6780
rect 24581 6743 24639 6749
rect 25222 6740 25228 6752
rect 25280 6740 25286 6792
rect 20438 6712 20444 6724
rect 13648 6684 20444 6712
rect 13449 6675 13507 6681
rect 13464 6644 13492 6675
rect 20438 6672 20444 6684
rect 20496 6672 20502 6724
rect 21082 6672 21088 6724
rect 21140 6712 21146 6724
rect 26421 6715 26479 6721
rect 26421 6712 26433 6715
rect 21140 6684 26433 6712
rect 21140 6672 21146 6684
rect 26421 6681 26433 6684
rect 26467 6712 26479 6715
rect 27338 6712 27344 6724
rect 26467 6684 27344 6712
rect 26467 6681 26479 6684
rect 26421 6675 26479 6681
rect 27338 6672 27344 6684
rect 27396 6672 27402 6724
rect 27816 6656 27844 6820
rect 32306 6808 32312 6820
rect 32364 6808 32370 6860
rect 39224 6857 39252 6888
rect 40126 6876 40132 6888
rect 40184 6876 40190 6928
rect 48041 6919 48099 6925
rect 48041 6885 48053 6919
rect 48087 6885 48099 6919
rect 48041 6879 48099 6885
rect 39209 6851 39267 6857
rect 39209 6817 39221 6851
rect 39255 6817 39267 6851
rect 39209 6811 39267 6817
rect 31018 6740 31024 6792
rect 31076 6780 31082 6792
rect 31113 6783 31171 6789
rect 31113 6780 31125 6783
rect 31076 6752 31125 6780
rect 31076 6740 31082 6752
rect 31113 6749 31125 6752
rect 31159 6749 31171 6783
rect 31113 6743 31171 6749
rect 31297 6783 31355 6789
rect 31297 6749 31309 6783
rect 31343 6780 31355 6783
rect 31478 6780 31484 6792
rect 31343 6752 31484 6780
rect 31343 6749 31355 6752
rect 31297 6743 31355 6749
rect 31478 6740 31484 6752
rect 31536 6780 31542 6792
rect 34698 6780 34704 6792
rect 31536 6752 34704 6780
rect 31536 6740 31542 6752
rect 34698 6740 34704 6752
rect 34756 6740 34762 6792
rect 35526 6780 35532 6792
rect 35487 6752 35532 6780
rect 35526 6740 35532 6752
rect 35584 6740 35590 6792
rect 35802 6780 35808 6792
rect 35763 6752 35808 6780
rect 35802 6740 35808 6752
rect 35860 6740 35866 6792
rect 27982 6672 27988 6724
rect 28040 6712 28046 6724
rect 38013 6715 38071 6721
rect 38013 6712 38025 6715
rect 28040 6684 38025 6712
rect 28040 6672 28046 6684
rect 38013 6681 38025 6684
rect 38059 6712 38071 6715
rect 38470 6712 38476 6724
rect 38059 6684 38476 6712
rect 38059 6681 38071 6684
rect 38013 6675 38071 6681
rect 38470 6672 38476 6684
rect 38528 6712 38534 6724
rect 38657 6715 38715 6721
rect 38657 6712 38669 6715
rect 38528 6684 38669 6712
rect 38528 6672 38534 6684
rect 38657 6681 38669 6684
rect 38703 6681 38715 6715
rect 38657 6675 38715 6681
rect 14093 6647 14151 6653
rect 14093 6644 14105 6647
rect 13464 6616 14105 6644
rect 14093 6613 14105 6616
rect 14139 6613 14151 6647
rect 14093 6607 14151 6613
rect 16577 6647 16635 6653
rect 16577 6613 16589 6647
rect 16623 6644 16635 6647
rect 17218 6644 17224 6656
rect 16623 6616 17224 6644
rect 16623 6613 16635 6616
rect 16577 6607 16635 6613
rect 17218 6604 17224 6616
rect 17276 6604 17282 6656
rect 21358 6604 21364 6656
rect 21416 6644 21422 6656
rect 27617 6647 27675 6653
rect 27617 6644 27629 6647
rect 21416 6616 27629 6644
rect 21416 6604 21422 6616
rect 27617 6613 27629 6616
rect 27663 6644 27675 6647
rect 27798 6644 27804 6656
rect 27663 6616 27804 6644
rect 27663 6613 27675 6616
rect 27617 6607 27675 6613
rect 27798 6604 27804 6616
rect 27856 6604 27862 6656
rect 31202 6644 31208 6656
rect 31163 6616 31208 6644
rect 31202 6604 31208 6616
rect 31260 6604 31266 6656
rect 35621 6647 35679 6653
rect 35621 6613 35633 6647
rect 35667 6644 35679 6647
rect 36998 6644 37004 6656
rect 35667 6616 37004 6644
rect 35667 6613 35679 6616
rect 35621 6607 35679 6613
rect 36998 6604 37004 6616
rect 37056 6604 37062 6656
rect 38102 6644 38108 6656
rect 38063 6616 38108 6644
rect 38102 6604 38108 6616
rect 38160 6604 38166 6656
rect 39224 6644 39252 6811
rect 45186 6808 45192 6860
rect 45244 6848 45250 6860
rect 45244 6820 45416 6848
rect 45244 6808 45250 6820
rect 39853 6783 39911 6789
rect 39853 6749 39865 6783
rect 39899 6780 39911 6783
rect 39942 6780 39948 6792
rect 39899 6752 39948 6780
rect 39899 6749 39911 6752
rect 39853 6743 39911 6749
rect 39942 6740 39948 6752
rect 40000 6740 40006 6792
rect 45388 6789 45416 6820
rect 45462 6808 45468 6860
rect 45520 6848 45526 6860
rect 47670 6848 47676 6860
rect 45520 6820 47676 6848
rect 45520 6808 45526 6820
rect 47670 6808 47676 6820
rect 47728 6848 47734 6860
rect 47765 6851 47823 6857
rect 47765 6848 47777 6851
rect 47728 6820 47777 6848
rect 47728 6808 47734 6820
rect 47765 6817 47777 6820
rect 47811 6817 47823 6851
rect 47765 6811 47823 6817
rect 47946 6808 47952 6860
rect 48004 6848 48010 6860
rect 48056 6848 48084 6879
rect 48004 6820 48084 6848
rect 48225 6851 48283 6857
rect 48004 6808 48010 6820
rect 48225 6817 48237 6851
rect 48271 6848 48283 6851
rect 54665 6851 54723 6857
rect 48271 6820 48912 6848
rect 48271 6817 48283 6820
rect 48225 6811 48283 6817
rect 48884 6789 48912 6820
rect 54665 6817 54677 6851
rect 54711 6848 54723 6851
rect 55401 6851 55459 6857
rect 55401 6848 55413 6851
rect 54711 6820 55413 6848
rect 54711 6817 54723 6820
rect 54665 6811 54723 6817
rect 55401 6817 55413 6820
rect 55447 6817 55459 6851
rect 56686 6848 56692 6860
rect 55401 6811 55459 6817
rect 55876 6820 56692 6848
rect 45373 6783 45431 6789
rect 45373 6749 45385 6783
rect 45419 6749 45431 6783
rect 45373 6743 45431 6749
rect 48869 6783 48927 6789
rect 48869 6749 48881 6783
rect 48915 6749 48927 6783
rect 48869 6743 48927 6749
rect 49145 6783 49203 6789
rect 49145 6749 49157 6783
rect 49191 6780 49203 6783
rect 49510 6780 49516 6792
rect 49191 6752 49516 6780
rect 49191 6749 49203 6752
rect 49145 6743 49203 6749
rect 49510 6740 49516 6752
rect 49568 6740 49574 6792
rect 54570 6780 54576 6792
rect 54531 6752 54576 6780
rect 54570 6740 54576 6752
rect 54628 6740 54634 6792
rect 54757 6783 54815 6789
rect 54757 6749 54769 6783
rect 54803 6780 54815 6783
rect 54938 6780 54944 6792
rect 54803 6752 54944 6780
rect 54803 6749 54815 6752
rect 54757 6743 54815 6749
rect 54938 6740 54944 6752
rect 54996 6740 55002 6792
rect 55490 6780 55496 6792
rect 55451 6752 55496 6780
rect 55490 6740 55496 6752
rect 55548 6740 55554 6792
rect 40034 6672 40040 6724
rect 40092 6712 40098 6724
rect 40129 6715 40187 6721
rect 40129 6712 40141 6715
rect 40092 6684 40141 6712
rect 40092 6672 40098 6684
rect 40129 6681 40141 6684
rect 40175 6681 40187 6715
rect 40129 6675 40187 6681
rect 45002 6672 45008 6724
rect 45060 6712 45066 6724
rect 45189 6715 45247 6721
rect 45189 6712 45201 6715
rect 45060 6684 45201 6712
rect 45060 6672 45066 6684
rect 45189 6681 45201 6684
rect 45235 6681 45247 6715
rect 45189 6675 45247 6681
rect 55398 6672 55404 6724
rect 55456 6712 55462 6724
rect 55876 6712 55904 6820
rect 56060 6789 56088 6820
rect 56686 6808 56692 6820
rect 56744 6848 56750 6860
rect 57241 6851 57299 6857
rect 57241 6848 57253 6851
rect 56744 6820 57253 6848
rect 56744 6808 56750 6820
rect 57241 6817 57253 6820
rect 57287 6848 57299 6851
rect 57793 6851 57851 6857
rect 57793 6848 57805 6851
rect 57287 6820 57805 6848
rect 57287 6817 57299 6820
rect 57241 6811 57299 6817
rect 57793 6817 57805 6820
rect 57839 6817 57851 6851
rect 57793 6811 57851 6817
rect 55953 6783 56011 6789
rect 55953 6749 55965 6783
rect 55999 6749 56011 6783
rect 55953 6743 56011 6749
rect 56045 6783 56103 6789
rect 56045 6749 56057 6783
rect 56091 6749 56103 6783
rect 56226 6780 56232 6792
rect 56187 6752 56232 6780
rect 56045 6743 56103 6749
rect 55456 6684 55904 6712
rect 55968 6712 55996 6743
rect 56226 6740 56232 6752
rect 56284 6740 56290 6792
rect 56778 6780 56784 6792
rect 56739 6752 56784 6780
rect 56778 6740 56784 6752
rect 56836 6740 56842 6792
rect 56870 6712 56876 6724
rect 55968 6684 56876 6712
rect 55456 6672 55462 6684
rect 56870 6672 56876 6684
rect 56928 6672 56934 6724
rect 39945 6647 40003 6653
rect 39945 6644 39957 6647
rect 39224 6616 39957 6644
rect 39945 6613 39957 6616
rect 39991 6613 40003 6647
rect 49050 6644 49056 6656
rect 49011 6616 49056 6644
rect 39945 6607 40003 6613
rect 49050 6604 49056 6616
rect 49108 6604 49114 6656
rect 1104 6554 58880 6576
rect 1104 6502 19574 6554
rect 19626 6502 19638 6554
rect 19690 6502 19702 6554
rect 19754 6502 19766 6554
rect 19818 6502 19830 6554
rect 19882 6502 50294 6554
rect 50346 6502 50358 6554
rect 50410 6502 50422 6554
rect 50474 6502 50486 6554
rect 50538 6502 50550 6554
rect 50602 6502 58880 6554
rect 1104 6480 58880 6502
rect 6822 6440 6828 6452
rect 6783 6412 6828 6440
rect 6822 6400 6828 6412
rect 6880 6400 6886 6452
rect 10505 6443 10563 6449
rect 10505 6409 10517 6443
rect 10551 6440 10563 6443
rect 12802 6440 12808 6452
rect 10551 6412 12808 6440
rect 10551 6409 10563 6412
rect 10505 6403 10563 6409
rect 12802 6400 12808 6412
rect 12860 6400 12866 6452
rect 20990 6440 20996 6452
rect 13924 6412 20996 6440
rect 3510 6332 3516 6384
rect 3568 6332 3574 6384
rect 4706 6372 4712 6384
rect 4080 6344 4712 6372
rect 1578 6264 1584 6316
rect 1636 6304 1642 6316
rect 1857 6307 1915 6313
rect 1857 6304 1869 6307
rect 1636 6276 1869 6304
rect 1636 6264 1642 6276
rect 1857 6273 1869 6276
rect 1903 6273 1915 6307
rect 3418 6304 3424 6316
rect 3379 6276 3424 6304
rect 1857 6267 1915 6273
rect 3418 6264 3424 6276
rect 3476 6264 3482 6316
rect 4080 6313 4108 6344
rect 4706 6332 4712 6344
rect 4764 6372 4770 6384
rect 10226 6372 10232 6384
rect 4764 6344 10232 6372
rect 4764 6332 4770 6344
rect 10226 6332 10232 6344
rect 10284 6332 10290 6384
rect 10410 6332 10416 6384
rect 10468 6332 10474 6384
rect 11606 6332 11612 6384
rect 11664 6372 11670 6384
rect 12161 6375 12219 6381
rect 12161 6372 12173 6375
rect 11664 6344 12173 6372
rect 11664 6332 11670 6344
rect 12161 6341 12173 6344
rect 12207 6372 12219 6375
rect 13924 6372 13952 6412
rect 20990 6400 20996 6412
rect 21048 6400 21054 6452
rect 23658 6400 23664 6452
rect 23716 6440 23722 6452
rect 24029 6443 24087 6449
rect 24029 6440 24041 6443
rect 23716 6412 24041 6440
rect 23716 6400 23722 6412
rect 24029 6409 24041 6412
rect 24075 6409 24087 6443
rect 27709 6443 27767 6449
rect 27709 6440 27721 6443
rect 24029 6403 24087 6409
rect 26344 6412 27721 6440
rect 12207 6344 12434 6372
rect 12207 6341 12219 6344
rect 12161 6335 12219 6341
rect 4065 6307 4123 6313
rect 4065 6273 4077 6307
rect 4111 6273 4123 6307
rect 4065 6267 4123 6273
rect 7193 6307 7251 6313
rect 7193 6273 7205 6307
rect 7239 6273 7251 6307
rect 10042 6304 10048 6316
rect 10003 6276 10048 6304
rect 7193 6267 7251 6273
rect 2038 6168 2044 6180
rect 1999 6140 2044 6168
rect 2038 6128 2044 6140
rect 2096 6128 2102 6180
rect 7208 6168 7236 6267
rect 10042 6264 10048 6276
rect 10100 6264 10106 6316
rect 10134 6264 10140 6316
rect 10192 6304 10198 6316
rect 10428 6304 10456 6332
rect 10508 6307 10566 6313
rect 10508 6304 10520 6307
rect 10192 6276 10237 6304
rect 10428 6276 10520 6304
rect 10192 6264 10198 6276
rect 10508 6273 10520 6276
rect 10554 6273 10566 6307
rect 12406 6304 12434 6344
rect 12728 6344 13952 6372
rect 12728 6313 12756 6344
rect 13998 6332 14004 6384
rect 14056 6372 14062 6384
rect 21082 6372 21088 6384
rect 14056 6344 21088 6372
rect 14056 6332 14062 6344
rect 21082 6332 21088 6344
rect 21140 6332 21146 6384
rect 24489 6375 24547 6381
rect 24489 6341 24501 6375
rect 24535 6372 24547 6375
rect 25222 6372 25228 6384
rect 24535 6344 25228 6372
rect 24535 6341 24547 6344
rect 24489 6335 24547 6341
rect 25222 6332 25228 6344
rect 25280 6332 25286 6384
rect 12713 6307 12771 6313
rect 12713 6304 12725 6307
rect 12406 6276 12725 6304
rect 10508 6267 10566 6273
rect 12713 6273 12725 6276
rect 12759 6273 12771 6307
rect 12713 6267 12771 6273
rect 12897 6307 12955 6313
rect 12897 6273 12909 6307
rect 12943 6273 12955 6307
rect 12897 6267 12955 6273
rect 13449 6307 13507 6313
rect 13449 6273 13461 6307
rect 13495 6304 13507 6307
rect 13538 6304 13544 6316
rect 13495 6276 13544 6304
rect 13495 6273 13507 6276
rect 13449 6267 13507 6273
rect 7285 6239 7343 6245
rect 7285 6205 7297 6239
rect 7331 6236 7343 6239
rect 8297 6239 8355 6245
rect 8297 6236 8309 6239
rect 7331 6208 8309 6236
rect 7331 6205 7343 6208
rect 7285 6199 7343 6205
rect 8297 6205 8309 6208
rect 8343 6205 8355 6239
rect 8297 6199 8355 6205
rect 8021 6171 8079 6177
rect 8021 6168 8033 6171
rect 7208 6140 8033 6168
rect 8021 6137 8033 6140
rect 8067 6137 8079 6171
rect 8312 6168 8340 6199
rect 10410 6196 10416 6248
rect 10468 6236 10474 6248
rect 12912 6236 12940 6267
rect 13538 6264 13544 6276
rect 13596 6264 13602 6316
rect 13630 6264 13636 6316
rect 13688 6304 13694 6316
rect 13688 6276 13733 6304
rect 13688 6264 13694 6276
rect 16574 6264 16580 6316
rect 16632 6304 16638 6316
rect 16669 6307 16727 6313
rect 16669 6304 16681 6307
rect 16632 6276 16681 6304
rect 16632 6264 16638 6276
rect 16669 6273 16681 6276
rect 16715 6273 16727 6307
rect 16850 6304 16856 6316
rect 16811 6276 16856 6304
rect 16669 6267 16727 6273
rect 16850 6264 16856 6276
rect 16908 6264 16914 6316
rect 17218 6264 17224 6316
rect 17276 6304 17282 6316
rect 17497 6307 17555 6313
rect 17497 6304 17509 6307
rect 17276 6276 17509 6304
rect 17276 6264 17282 6276
rect 17497 6273 17509 6276
rect 17543 6273 17555 6307
rect 17497 6267 17555 6273
rect 17681 6307 17739 6313
rect 17681 6273 17693 6307
rect 17727 6304 17739 6307
rect 17954 6304 17960 6316
rect 17727 6276 17960 6304
rect 17727 6273 17739 6276
rect 17681 6267 17739 6273
rect 17954 6264 17960 6276
rect 18012 6264 18018 6316
rect 20254 6304 20260 6316
rect 20215 6276 20260 6304
rect 20254 6264 20260 6276
rect 20312 6264 20318 6316
rect 20438 6264 20444 6316
rect 20496 6304 20502 6316
rect 26234 6304 26240 6316
rect 20496 6276 26240 6304
rect 20496 6264 20502 6276
rect 26234 6264 26240 6276
rect 26292 6304 26298 6316
rect 26344 6313 26372 6412
rect 27709 6409 27721 6412
rect 27755 6409 27767 6443
rect 27709 6403 27767 6409
rect 33594 6400 33600 6452
rect 33652 6440 33658 6452
rect 38654 6440 38660 6452
rect 33652 6412 38660 6440
rect 33652 6400 33658 6412
rect 38654 6400 38660 6412
rect 38712 6400 38718 6452
rect 38838 6440 38844 6452
rect 38799 6412 38844 6440
rect 38838 6400 38844 6412
rect 38896 6400 38902 6452
rect 54757 6443 54815 6449
rect 54757 6409 54769 6443
rect 54803 6440 54815 6443
rect 55490 6440 55496 6452
rect 54803 6412 55496 6440
rect 54803 6409 54815 6412
rect 54757 6403 54815 6409
rect 55490 6400 55496 6412
rect 55548 6400 55554 6452
rect 56870 6440 56876 6452
rect 56831 6412 56876 6440
rect 56870 6400 56876 6412
rect 56928 6400 56934 6452
rect 57054 6400 57060 6452
rect 57112 6440 57118 6452
rect 57241 6443 57299 6449
rect 57241 6440 57253 6443
rect 57112 6412 57253 6440
rect 57112 6400 57118 6412
rect 57241 6409 57253 6412
rect 57287 6409 57299 6443
rect 57241 6403 57299 6409
rect 27614 6332 27620 6384
rect 27672 6332 27678 6384
rect 35529 6375 35587 6381
rect 35529 6341 35541 6375
rect 35575 6372 35587 6375
rect 35802 6372 35808 6384
rect 35575 6344 35808 6372
rect 35575 6341 35587 6344
rect 35529 6335 35587 6341
rect 35802 6332 35808 6344
rect 35860 6332 35866 6384
rect 43530 6372 43536 6384
rect 37384 6344 39988 6372
rect 43491 6344 43536 6372
rect 26329 6307 26387 6313
rect 26329 6304 26341 6307
rect 26292 6276 26341 6304
rect 26292 6264 26298 6276
rect 26329 6273 26341 6276
rect 26375 6273 26387 6307
rect 27632 6304 27660 6332
rect 26329 6267 26387 6273
rect 27540 6276 27660 6304
rect 19978 6236 19984 6248
rect 10468 6208 12940 6236
rect 19939 6208 19984 6236
rect 10468 6196 10474 6208
rect 10689 6171 10747 6177
rect 10689 6168 10701 6171
rect 8312 6140 10701 6168
rect 8021 6131 8079 6137
rect 10689 6137 10701 6140
rect 10735 6137 10747 6171
rect 12912 6168 12940 6208
rect 19978 6196 19984 6208
rect 20036 6196 20042 6248
rect 20346 6196 20352 6248
rect 20404 6236 20410 6248
rect 27540 6245 27568 6276
rect 31018 6264 31024 6316
rect 31076 6304 31082 6316
rect 31389 6307 31447 6313
rect 31389 6304 31401 6307
rect 31076 6276 31401 6304
rect 31076 6264 31082 6276
rect 31389 6273 31401 6276
rect 31435 6273 31447 6307
rect 31389 6267 31447 6273
rect 31478 6264 31484 6316
rect 31536 6304 31542 6316
rect 31536 6276 31581 6304
rect 31536 6264 31542 6276
rect 34698 6264 34704 6316
rect 34756 6304 34762 6316
rect 35710 6304 35716 6316
rect 34756 6276 35716 6304
rect 34756 6264 34762 6276
rect 35710 6264 35716 6276
rect 35768 6304 35774 6316
rect 36173 6307 36231 6313
rect 36173 6304 36185 6307
rect 35768 6276 36185 6304
rect 35768 6264 35774 6276
rect 36173 6273 36185 6276
rect 36219 6273 36231 6307
rect 36173 6267 36231 6273
rect 36357 6307 36415 6313
rect 36357 6273 36369 6307
rect 36403 6304 36415 6307
rect 36998 6304 37004 6316
rect 36403 6276 37004 6304
rect 36403 6273 36415 6276
rect 36357 6267 36415 6273
rect 36998 6264 37004 6276
rect 37056 6304 37062 6316
rect 37384 6313 37412 6344
rect 39960 6316 39988 6344
rect 43530 6332 43536 6344
rect 43588 6332 43594 6384
rect 44634 6332 44640 6384
rect 44692 6372 44698 6384
rect 44692 6344 57928 6372
rect 44692 6332 44698 6344
rect 37369 6307 37427 6313
rect 37369 6304 37381 6307
rect 37056 6276 37381 6304
rect 37056 6264 37062 6276
rect 37369 6273 37381 6276
rect 37415 6273 37427 6307
rect 37369 6267 37427 6273
rect 37458 6264 37464 6316
rect 37516 6304 37522 6316
rect 37516 6276 37561 6304
rect 37516 6264 37522 6276
rect 38838 6264 38844 6316
rect 38896 6304 38902 6316
rect 39669 6307 39727 6313
rect 39669 6304 39681 6307
rect 38896 6276 39681 6304
rect 38896 6264 38902 6276
rect 39669 6273 39681 6276
rect 39715 6273 39727 6307
rect 39942 6304 39948 6316
rect 39903 6276 39948 6304
rect 39669 6267 39727 6273
rect 39942 6264 39948 6276
rect 40000 6264 40006 6316
rect 47670 6304 47676 6316
rect 47631 6276 47676 6304
rect 47670 6264 47676 6276
rect 47728 6264 47734 6316
rect 47946 6304 47952 6316
rect 47907 6276 47952 6304
rect 47946 6264 47952 6276
rect 48004 6264 48010 6316
rect 48685 6307 48743 6313
rect 48685 6273 48697 6307
rect 48731 6304 48743 6307
rect 49050 6304 49056 6316
rect 48731 6276 49056 6304
rect 48731 6273 48743 6276
rect 48685 6267 48743 6273
rect 49050 6264 49056 6276
rect 49108 6304 49114 6316
rect 49329 6307 49387 6313
rect 49329 6304 49341 6307
rect 49108 6276 49341 6304
rect 49108 6264 49114 6276
rect 49329 6273 49341 6276
rect 49375 6273 49387 6307
rect 49329 6267 49387 6273
rect 49510 6264 49516 6316
rect 49568 6264 49574 6316
rect 50341 6307 50399 6313
rect 50341 6273 50353 6307
rect 50387 6304 50399 6307
rect 51258 6304 51264 6316
rect 50387 6276 51264 6304
rect 50387 6273 50399 6276
rect 50341 6267 50399 6273
rect 51258 6264 51264 6276
rect 51316 6264 51322 6316
rect 53558 6264 53564 6316
rect 53616 6304 53622 6316
rect 53929 6307 53987 6313
rect 53929 6304 53941 6307
rect 53616 6276 53941 6304
rect 53616 6264 53622 6276
rect 53929 6273 53941 6276
rect 53975 6273 53987 6307
rect 54570 6304 54576 6316
rect 53929 6267 53987 6273
rect 54036 6276 54576 6304
rect 20809 6239 20867 6245
rect 20809 6236 20821 6239
rect 20404 6208 20821 6236
rect 20404 6196 20410 6208
rect 20809 6205 20821 6208
rect 20855 6205 20867 6239
rect 20809 6199 20867 6205
rect 27525 6239 27583 6245
rect 27525 6205 27537 6239
rect 27571 6205 27583 6239
rect 27525 6199 27583 6205
rect 27617 6239 27675 6245
rect 27617 6205 27629 6239
rect 27663 6236 27675 6239
rect 27798 6236 27804 6248
rect 27663 6208 27804 6236
rect 27663 6205 27675 6208
rect 27617 6199 27675 6205
rect 27798 6196 27804 6208
rect 27856 6196 27862 6248
rect 37734 6196 37740 6248
rect 37792 6236 37798 6248
rect 40218 6236 40224 6248
rect 37792 6208 40224 6236
rect 37792 6196 37798 6208
rect 40218 6196 40224 6208
rect 40276 6196 40282 6248
rect 40402 6236 40408 6248
rect 40363 6208 40408 6236
rect 40402 6196 40408 6208
rect 40460 6196 40466 6248
rect 54036 6245 54064 6276
rect 54570 6264 54576 6276
rect 54628 6304 54634 6316
rect 55033 6307 55091 6313
rect 55033 6304 55045 6307
rect 54628 6276 55045 6304
rect 54628 6264 54634 6276
rect 55033 6273 55045 6276
rect 55079 6273 55091 6307
rect 55033 6267 55091 6273
rect 55401 6307 55459 6313
rect 55401 6273 55413 6307
rect 55447 6304 55459 6307
rect 56134 6304 56140 6316
rect 55447 6276 56140 6304
rect 55447 6273 55459 6276
rect 55401 6267 55459 6273
rect 56134 6264 56140 6276
rect 56192 6264 56198 6316
rect 56686 6264 56692 6316
rect 56744 6304 56750 6316
rect 56781 6307 56839 6313
rect 56781 6304 56793 6307
rect 56744 6276 56793 6304
rect 56744 6264 56750 6276
rect 56781 6273 56793 6276
rect 56827 6273 56839 6307
rect 56781 6267 56839 6273
rect 57057 6307 57115 6313
rect 57057 6273 57069 6307
rect 57103 6273 57115 6307
rect 57057 6267 57115 6273
rect 54021 6239 54079 6245
rect 54021 6205 54033 6239
rect 54067 6205 54079 6239
rect 54938 6236 54944 6248
rect 54899 6208 54944 6236
rect 54021 6199 54079 6205
rect 54938 6196 54944 6208
rect 54996 6196 55002 6248
rect 55309 6239 55367 6245
rect 55309 6205 55321 6239
rect 55355 6236 55367 6239
rect 55766 6236 55772 6248
rect 55355 6208 55772 6236
rect 55355 6205 55367 6208
rect 55309 6199 55367 6205
rect 55766 6196 55772 6208
rect 55824 6236 55830 6248
rect 55953 6239 56011 6245
rect 55953 6236 55965 6239
rect 55824 6208 55965 6236
rect 55824 6196 55830 6208
rect 55953 6205 55965 6208
rect 55999 6205 56011 6239
rect 55953 6199 56011 6205
rect 56321 6239 56379 6245
rect 56321 6205 56333 6239
rect 56367 6236 56379 6239
rect 57072 6236 57100 6267
rect 57790 6264 57796 6316
rect 57848 6304 57854 6316
rect 57900 6313 57928 6344
rect 57885 6307 57943 6313
rect 57885 6304 57897 6307
rect 57848 6276 57897 6304
rect 57848 6264 57854 6276
rect 57885 6273 57897 6276
rect 57931 6273 57943 6307
rect 57885 6267 57943 6273
rect 56367 6208 57100 6236
rect 56367 6205 56379 6208
rect 56321 6199 56379 6205
rect 20364 6168 20392 6196
rect 24210 6168 24216 6180
rect 12912 6140 20392 6168
rect 24171 6140 24216 6168
rect 10689 6131 10747 6137
rect 7190 6060 7196 6112
rect 7248 6100 7254 6112
rect 7837 6103 7895 6109
rect 7837 6100 7849 6103
rect 7248 6072 7849 6100
rect 7248 6060 7254 6072
rect 7837 6069 7849 6072
rect 7883 6069 7895 6103
rect 8036 6100 8064 6131
rect 24210 6128 24216 6140
rect 24268 6128 24274 6180
rect 28077 6171 28135 6177
rect 28077 6137 28089 6171
rect 28123 6168 28135 6171
rect 37458 6168 37464 6180
rect 28123 6140 37464 6168
rect 28123 6137 28135 6140
rect 28077 6131 28135 6137
rect 37458 6128 37464 6140
rect 37516 6128 37522 6180
rect 40126 6128 40132 6180
rect 40184 6168 40190 6180
rect 43809 6171 43867 6177
rect 43809 6168 43821 6171
rect 40184 6140 43821 6168
rect 40184 6128 40190 6140
rect 43548 6112 43576 6140
rect 43809 6137 43821 6140
rect 43855 6137 43867 6171
rect 43809 6131 43867 6137
rect 54297 6171 54355 6177
rect 54297 6137 54309 6171
rect 54343 6168 54355 6171
rect 56226 6168 56232 6180
rect 54343 6140 56232 6168
rect 54343 6137 54355 6140
rect 54297 6131 54355 6137
rect 56226 6128 56232 6140
rect 56284 6128 56290 6180
rect 58066 6168 58072 6180
rect 58027 6140 58072 6168
rect 58066 6128 58072 6140
rect 58124 6128 58130 6180
rect 9674 6100 9680 6112
rect 8036 6072 9680 6100
rect 7837 6063 7895 6069
rect 9674 6060 9680 6072
rect 9732 6060 9738 6112
rect 13446 6060 13452 6112
rect 13504 6100 13510 6112
rect 13541 6103 13599 6109
rect 13541 6100 13553 6103
rect 13504 6072 13553 6100
rect 13504 6060 13510 6072
rect 13541 6069 13553 6072
rect 13587 6069 13599 6103
rect 16758 6100 16764 6112
rect 16719 6072 16764 6100
rect 13541 6063 13599 6069
rect 16758 6060 16764 6072
rect 16816 6060 16822 6112
rect 17037 6103 17095 6109
rect 17037 6069 17049 6103
rect 17083 6100 17095 6103
rect 17586 6100 17592 6112
rect 17083 6072 17592 6100
rect 17083 6069 17095 6072
rect 17037 6063 17095 6069
rect 17586 6060 17592 6072
rect 17644 6060 17650 6112
rect 17678 6060 17684 6112
rect 17736 6100 17742 6112
rect 31205 6103 31263 6109
rect 17736 6072 17781 6100
rect 17736 6060 17742 6072
rect 31205 6069 31217 6103
rect 31251 6100 31263 6103
rect 31386 6100 31392 6112
rect 31251 6072 31392 6100
rect 31251 6069 31263 6072
rect 31205 6063 31263 6069
rect 31386 6060 31392 6072
rect 31444 6100 31450 6112
rect 32030 6100 32036 6112
rect 31444 6072 32036 6100
rect 31444 6060 31450 6072
rect 32030 6060 32036 6072
rect 32088 6060 32094 6112
rect 35434 6100 35440 6112
rect 35395 6072 35440 6100
rect 35434 6060 35440 6072
rect 35492 6060 35498 6112
rect 37645 6103 37703 6109
rect 37645 6069 37657 6103
rect 37691 6100 37703 6103
rect 37826 6100 37832 6112
rect 37691 6072 37832 6100
rect 37691 6069 37703 6072
rect 37645 6063 37703 6069
rect 37826 6060 37832 6072
rect 37884 6060 37890 6112
rect 43530 6060 43536 6112
rect 43588 6060 43594 6112
rect 43993 6103 44051 6109
rect 43993 6069 44005 6103
rect 44039 6100 44051 6103
rect 44450 6100 44456 6112
rect 44039 6072 44456 6100
rect 44039 6069 44051 6072
rect 43993 6063 44051 6069
rect 44450 6060 44456 6072
rect 44508 6060 44514 6112
rect 53285 6103 53343 6109
rect 53285 6069 53297 6103
rect 53331 6100 53343 6103
rect 53558 6100 53564 6112
rect 53331 6072 53564 6100
rect 53331 6069 53343 6072
rect 53285 6063 53343 6069
rect 53558 6060 53564 6072
rect 53616 6060 53622 6112
rect 1104 6010 58880 6032
rect 1104 5958 4214 6010
rect 4266 5958 4278 6010
rect 4330 5958 4342 6010
rect 4394 5958 4406 6010
rect 4458 5958 4470 6010
rect 4522 5958 34934 6010
rect 34986 5958 34998 6010
rect 35050 5958 35062 6010
rect 35114 5958 35126 6010
rect 35178 5958 35190 6010
rect 35242 5958 58880 6010
rect 1104 5936 58880 5958
rect 1578 5896 1584 5908
rect 1539 5868 1584 5896
rect 1578 5856 1584 5868
rect 1636 5856 1642 5908
rect 10042 5856 10048 5908
rect 10100 5896 10106 5908
rect 10137 5899 10195 5905
rect 10137 5896 10149 5899
rect 10100 5868 10149 5896
rect 10100 5856 10106 5868
rect 10137 5865 10149 5868
rect 10183 5865 10195 5899
rect 17681 5899 17739 5905
rect 17681 5896 17693 5899
rect 10137 5859 10195 5865
rect 16132 5868 17693 5896
rect 6822 5828 6828 5840
rect 6656 5800 6828 5828
rect 4341 5763 4399 5769
rect 4341 5729 4353 5763
rect 4387 5760 4399 5763
rect 4614 5760 4620 5772
rect 4387 5732 4620 5760
rect 4387 5729 4399 5732
rect 4341 5723 4399 5729
rect 4614 5720 4620 5732
rect 4672 5720 4678 5772
rect 6656 5769 6684 5800
rect 6822 5788 6828 5800
rect 6880 5788 6886 5840
rect 16025 5831 16083 5837
rect 16025 5828 16037 5831
rect 12406 5800 16037 5828
rect 6641 5763 6699 5769
rect 6641 5729 6653 5763
rect 6687 5729 6699 5763
rect 6641 5723 6699 5729
rect 6730 5720 6736 5772
rect 6788 5720 6794 5772
rect 7190 5760 7196 5772
rect 7151 5732 7196 5760
rect 7190 5720 7196 5732
rect 7248 5720 7254 5772
rect 10502 5760 10508 5772
rect 10463 5732 10508 5760
rect 10502 5720 10508 5732
rect 10560 5720 10566 5772
rect 5077 5695 5135 5701
rect 5077 5661 5089 5695
rect 5123 5661 5135 5695
rect 5077 5655 5135 5661
rect 5261 5695 5319 5701
rect 5261 5661 5273 5695
rect 5307 5661 5319 5695
rect 6748 5692 6776 5720
rect 6825 5695 6883 5701
rect 6825 5692 6837 5695
rect 6748 5664 6837 5692
rect 5261 5655 5319 5661
rect 6825 5661 6837 5664
rect 6871 5661 6883 5695
rect 10410 5692 10416 5704
rect 10371 5664 10416 5692
rect 6825 5655 6883 5661
rect 5092 5556 5120 5655
rect 5276 5624 5304 5655
rect 10410 5652 10416 5664
rect 10468 5652 10474 5704
rect 6730 5624 6736 5636
rect 5276 5596 6736 5624
rect 6730 5584 6736 5596
rect 6788 5624 6794 5636
rect 7101 5627 7159 5633
rect 7101 5624 7113 5627
rect 6788 5596 7113 5624
rect 6788 5584 6794 5596
rect 7101 5593 7113 5596
rect 7147 5593 7159 5627
rect 7101 5587 7159 5593
rect 6822 5556 6828 5568
rect 5092 5528 6828 5556
rect 6822 5516 6828 5528
rect 6880 5556 6886 5568
rect 12406 5556 12434 5800
rect 16025 5797 16037 5800
rect 16071 5797 16083 5831
rect 16025 5791 16083 5797
rect 12802 5760 12808 5772
rect 12763 5732 12808 5760
rect 12802 5720 12808 5732
rect 12860 5720 12866 5772
rect 13630 5720 13636 5772
rect 13688 5760 13694 5772
rect 16132 5760 16160 5868
rect 17681 5865 17693 5868
rect 17727 5865 17739 5899
rect 17681 5859 17739 5865
rect 20990 5856 20996 5908
rect 21048 5896 21054 5908
rect 27982 5896 27988 5908
rect 21048 5868 27988 5896
rect 21048 5856 21054 5868
rect 27982 5856 27988 5868
rect 28040 5856 28046 5908
rect 30653 5899 30711 5905
rect 30653 5865 30665 5899
rect 30699 5896 30711 5899
rect 31386 5896 31392 5908
rect 30699 5868 31392 5896
rect 30699 5865 30711 5868
rect 30653 5859 30711 5865
rect 31386 5856 31392 5868
rect 31444 5856 31450 5908
rect 32030 5896 32036 5908
rect 31991 5868 32036 5896
rect 32030 5856 32036 5868
rect 32088 5856 32094 5908
rect 54205 5899 54263 5905
rect 40144 5868 40356 5896
rect 17954 5828 17960 5840
rect 13688 5732 16160 5760
rect 16960 5800 17960 5828
rect 13688 5720 13694 5732
rect 12897 5695 12955 5701
rect 12897 5661 12909 5695
rect 12943 5692 12955 5695
rect 13998 5692 14004 5704
rect 12943 5664 14004 5692
rect 12943 5661 12955 5664
rect 12897 5655 12955 5661
rect 13998 5652 14004 5664
rect 14056 5652 14062 5704
rect 14292 5701 14320 5732
rect 14277 5695 14335 5701
rect 14277 5661 14289 5695
rect 14323 5661 14335 5695
rect 14277 5655 14335 5661
rect 16117 5695 16175 5701
rect 16117 5661 16129 5695
rect 16163 5661 16175 5695
rect 16117 5655 16175 5661
rect 16301 5695 16359 5701
rect 16301 5661 16313 5695
rect 16347 5692 16359 5695
rect 16574 5692 16580 5704
rect 16347 5664 16580 5692
rect 16347 5661 16359 5664
rect 16301 5655 16359 5661
rect 13538 5624 13544 5636
rect 13280 5596 13544 5624
rect 13280 5565 13308 5596
rect 13538 5584 13544 5596
rect 13596 5624 13602 5636
rect 14093 5627 14151 5633
rect 14093 5624 14105 5627
rect 13596 5596 14105 5624
rect 13596 5584 13602 5596
rect 14093 5593 14105 5596
rect 14139 5593 14151 5627
rect 16132 5624 16160 5655
rect 16574 5652 16580 5664
rect 16632 5652 16638 5704
rect 16960 5701 16988 5800
rect 17954 5788 17960 5800
rect 18012 5788 18018 5840
rect 19613 5831 19671 5837
rect 19613 5797 19625 5831
rect 19659 5828 19671 5831
rect 20162 5828 20168 5840
rect 19659 5800 20168 5828
rect 19659 5797 19671 5800
rect 19613 5791 19671 5797
rect 20162 5788 20168 5800
rect 20220 5788 20226 5840
rect 21177 5831 21235 5837
rect 21177 5797 21189 5831
rect 21223 5828 21235 5831
rect 27614 5828 27620 5840
rect 21223 5800 27620 5828
rect 21223 5797 21235 5800
rect 21177 5791 21235 5797
rect 17129 5763 17187 5769
rect 17129 5729 17141 5763
rect 17175 5760 17187 5763
rect 17218 5760 17224 5772
rect 17175 5732 17224 5760
rect 17175 5729 17187 5732
rect 17129 5723 17187 5729
rect 17218 5720 17224 5732
rect 17276 5760 17282 5772
rect 19978 5760 19984 5772
rect 17276 5732 17816 5760
rect 19891 5732 19984 5760
rect 17276 5720 17282 5732
rect 16945 5695 17003 5701
rect 16945 5661 16957 5695
rect 16991 5661 17003 5695
rect 17586 5692 17592 5704
rect 17547 5664 17592 5692
rect 16945 5655 17003 5661
rect 17586 5652 17592 5664
rect 17644 5652 17650 5704
rect 17788 5701 17816 5732
rect 19904 5701 19932 5732
rect 19978 5720 19984 5732
rect 20036 5760 20042 5772
rect 20441 5763 20499 5769
rect 20441 5760 20453 5763
rect 20036 5732 20453 5760
rect 20036 5720 20042 5732
rect 20441 5729 20453 5732
rect 20487 5729 20499 5763
rect 21192 5760 21220 5791
rect 27614 5788 27620 5800
rect 27672 5788 27678 5840
rect 31938 5828 31944 5840
rect 30484 5800 31944 5828
rect 20441 5723 20499 5729
rect 20548 5732 21220 5760
rect 17773 5695 17831 5701
rect 17773 5661 17785 5695
rect 17819 5661 17831 5695
rect 17773 5655 17831 5661
rect 19889 5695 19947 5701
rect 19889 5661 19901 5695
rect 19935 5661 19947 5695
rect 20346 5692 20352 5704
rect 20307 5664 20352 5692
rect 19889 5655 19947 5661
rect 20346 5652 20352 5664
rect 20404 5652 20410 5704
rect 20548 5701 20576 5732
rect 23014 5720 23020 5772
rect 23072 5760 23078 5772
rect 23072 5732 23513 5760
rect 23072 5720 23078 5732
rect 20533 5695 20591 5701
rect 20533 5661 20545 5695
rect 20579 5661 20591 5695
rect 20990 5692 20996 5704
rect 20951 5664 20996 5692
rect 20533 5655 20591 5661
rect 20990 5652 20996 5664
rect 21048 5652 21054 5704
rect 21082 5652 21088 5704
rect 21140 5692 21146 5704
rect 21177 5695 21235 5701
rect 21177 5692 21189 5695
rect 21140 5664 21189 5692
rect 21140 5652 21146 5664
rect 21177 5661 21189 5664
rect 21223 5661 21235 5695
rect 23290 5692 23296 5704
rect 23251 5664 23296 5692
rect 21177 5655 21235 5661
rect 23290 5652 23296 5664
rect 23348 5652 23354 5704
rect 23485 5701 23513 5732
rect 29638 5720 29644 5772
rect 29696 5760 29702 5772
rect 30484 5769 30512 5800
rect 31938 5788 31944 5800
rect 31996 5788 32002 5840
rect 35452 5800 36860 5828
rect 35452 5772 35480 5800
rect 30469 5763 30527 5769
rect 30469 5760 30481 5763
rect 29696 5732 30481 5760
rect 29696 5720 29702 5732
rect 30469 5729 30481 5732
rect 30515 5729 30527 5763
rect 32125 5763 32183 5769
rect 32125 5760 32137 5763
rect 30469 5723 30527 5729
rect 30760 5732 32137 5760
rect 23477 5695 23535 5701
rect 23477 5661 23489 5695
rect 23523 5692 23535 5695
rect 24026 5692 24032 5704
rect 23523 5664 24032 5692
rect 23523 5661 23535 5664
rect 23477 5655 23535 5661
rect 24026 5652 24032 5664
rect 24084 5692 24090 5704
rect 24397 5695 24455 5701
rect 24397 5692 24409 5695
rect 24084 5664 24409 5692
rect 24084 5652 24090 5664
rect 24397 5661 24409 5664
rect 24443 5661 24455 5695
rect 26970 5692 26976 5704
rect 26931 5664 26976 5692
rect 24397 5655 24455 5661
rect 26970 5652 26976 5664
rect 27028 5652 27034 5704
rect 27338 5692 27344 5704
rect 27299 5664 27344 5692
rect 27338 5652 27344 5664
rect 27396 5652 27402 5704
rect 30760 5701 30788 5732
rect 32125 5729 32137 5732
rect 32171 5760 32183 5763
rect 35434 5760 35440 5772
rect 32171 5732 35440 5760
rect 32171 5729 32183 5732
rect 32125 5723 32183 5729
rect 35434 5720 35440 5732
rect 35492 5720 35498 5772
rect 35710 5720 35716 5772
rect 35768 5760 35774 5772
rect 35989 5763 36047 5769
rect 35989 5760 36001 5763
rect 35768 5732 36001 5760
rect 35768 5720 35774 5732
rect 35989 5729 36001 5732
rect 36035 5729 36047 5763
rect 35989 5723 36047 5729
rect 35532 5704 35584 5710
rect 30745 5695 30803 5701
rect 30745 5661 30757 5695
rect 30791 5661 30803 5695
rect 31202 5692 31208 5704
rect 31163 5664 31208 5692
rect 30745 5655 30803 5661
rect 31202 5652 31208 5664
rect 31260 5652 31266 5704
rect 31386 5692 31392 5704
rect 31347 5664 31392 5692
rect 31386 5652 31392 5664
rect 31444 5652 31450 5704
rect 31938 5652 31944 5704
rect 31996 5692 32002 5704
rect 32033 5695 32091 5701
rect 32033 5692 32045 5695
rect 31996 5664 32045 5692
rect 31996 5652 32002 5664
rect 32033 5661 32045 5664
rect 32079 5661 32091 5695
rect 32033 5655 32091 5661
rect 33134 5652 33140 5704
rect 33192 5692 33198 5704
rect 33413 5695 33471 5701
rect 33413 5692 33425 5695
rect 33192 5664 33425 5692
rect 33192 5652 33198 5664
rect 33413 5661 33425 5664
rect 33459 5661 33471 5695
rect 33594 5692 33600 5704
rect 33555 5664 33600 5692
rect 33413 5655 33471 5661
rect 33594 5652 33600 5664
rect 33652 5652 33658 5704
rect 16761 5627 16819 5633
rect 16761 5624 16773 5627
rect 16132 5596 16773 5624
rect 14093 5587 14151 5593
rect 16761 5593 16773 5596
rect 16807 5593 16819 5627
rect 16761 5587 16819 5593
rect 17604 5596 19380 5624
rect 6880 5528 12434 5556
rect 13265 5559 13323 5565
rect 6880 5516 6886 5528
rect 13265 5525 13277 5559
rect 13311 5525 13323 5559
rect 14458 5556 14464 5568
rect 14419 5528 14464 5556
rect 13265 5519 13323 5525
rect 14458 5516 14464 5528
rect 14516 5556 14522 5568
rect 17604 5556 17632 5596
rect 19352 5568 19380 5596
rect 19426 5584 19432 5636
rect 19484 5624 19490 5636
rect 19613 5627 19671 5633
rect 19613 5624 19625 5627
rect 19484 5596 19625 5624
rect 19484 5584 19490 5596
rect 19613 5593 19625 5596
rect 19659 5593 19671 5627
rect 21008 5624 21036 5652
rect 35532 5646 35584 5652
rect 21637 5627 21695 5633
rect 21637 5624 21649 5627
rect 21008 5596 21649 5624
rect 19613 5587 19671 5593
rect 21637 5593 21649 5596
rect 21683 5593 21695 5627
rect 24578 5624 24584 5636
rect 24539 5596 24584 5624
rect 21637 5587 21695 5593
rect 24578 5584 24584 5596
rect 24636 5584 24642 5636
rect 26878 5584 26884 5636
rect 26936 5624 26942 5636
rect 27065 5627 27123 5633
rect 27065 5624 27077 5627
rect 26936 5596 27077 5624
rect 26936 5584 26942 5596
rect 27065 5593 27077 5596
rect 27111 5593 27123 5627
rect 27065 5587 27123 5593
rect 27157 5627 27215 5633
rect 27157 5593 27169 5627
rect 27203 5624 27215 5627
rect 35437 5627 35495 5633
rect 27203 5596 31248 5624
rect 27203 5593 27215 5596
rect 27157 5587 27215 5593
rect 19334 5556 19340 5568
rect 14516 5528 17632 5556
rect 19247 5528 19340 5556
rect 14516 5516 14522 5528
rect 19334 5516 19340 5528
rect 19392 5556 19398 5568
rect 19797 5559 19855 5565
rect 19797 5556 19809 5559
rect 19392 5528 19809 5556
rect 19392 5516 19398 5528
rect 19797 5525 19809 5528
rect 19843 5525 19855 5559
rect 23382 5556 23388 5568
rect 23343 5528 23388 5556
rect 19797 5519 19855 5525
rect 23382 5516 23388 5528
rect 23440 5516 23446 5568
rect 24762 5556 24768 5568
rect 24723 5528 24768 5556
rect 24762 5516 24768 5528
rect 24820 5516 24826 5568
rect 25314 5516 25320 5568
rect 25372 5556 25378 5568
rect 26789 5559 26847 5565
rect 26789 5556 26801 5559
rect 25372 5528 26801 5556
rect 25372 5516 25378 5528
rect 26789 5525 26801 5528
rect 26835 5525 26847 5559
rect 30466 5556 30472 5568
rect 30427 5528 30472 5556
rect 26789 5519 26847 5525
rect 30466 5516 30472 5528
rect 30524 5516 30530 5568
rect 31220 5556 31248 5596
rect 31496 5596 33272 5624
rect 31496 5556 31524 5596
rect 33244 5568 33272 5596
rect 35437 5593 35449 5627
rect 35483 5593 35495 5627
rect 36832 5624 36860 5800
rect 40144 5769 40172 5868
rect 40328 5828 40356 5868
rect 54205 5865 54217 5899
rect 54251 5896 54263 5899
rect 54938 5896 54944 5908
rect 54251 5868 54944 5896
rect 54251 5865 54263 5868
rect 54205 5859 54263 5865
rect 54938 5856 54944 5868
rect 54996 5856 55002 5908
rect 55493 5899 55551 5905
rect 55493 5865 55505 5899
rect 55539 5896 55551 5899
rect 55766 5896 55772 5908
rect 55539 5868 55772 5896
rect 55539 5865 55551 5868
rect 55493 5859 55551 5865
rect 55766 5856 55772 5868
rect 55824 5856 55830 5908
rect 57790 5896 57796 5908
rect 57751 5868 57796 5896
rect 57790 5856 57796 5868
rect 57848 5856 57854 5908
rect 40328 5800 41092 5828
rect 41064 5769 41092 5800
rect 37093 5763 37151 5769
rect 37093 5729 37105 5763
rect 37139 5760 37151 5763
rect 40129 5763 40187 5769
rect 40129 5760 40141 5763
rect 37139 5732 37688 5760
rect 37139 5729 37151 5732
rect 37093 5723 37151 5729
rect 36998 5692 37004 5704
rect 36959 5664 37004 5692
rect 36998 5652 37004 5664
rect 37056 5652 37062 5704
rect 37185 5695 37243 5701
rect 37185 5661 37197 5695
rect 37231 5692 37243 5695
rect 37458 5692 37464 5704
rect 37231 5664 37464 5692
rect 37231 5661 37243 5664
rect 37185 5655 37243 5661
rect 37458 5652 37464 5664
rect 37516 5652 37522 5704
rect 37660 5701 37688 5732
rect 37844 5732 40141 5760
rect 37844 5704 37872 5732
rect 40129 5729 40141 5732
rect 40175 5729 40187 5763
rect 40129 5723 40187 5729
rect 41049 5763 41107 5769
rect 41049 5729 41061 5763
rect 41095 5729 41107 5763
rect 43438 5760 43444 5772
rect 43399 5732 43444 5760
rect 41049 5723 41107 5729
rect 43438 5720 43444 5732
rect 43496 5720 43502 5772
rect 56870 5720 56876 5772
rect 56928 5760 56934 5772
rect 56965 5763 57023 5769
rect 56965 5760 56977 5763
rect 56928 5732 56977 5760
rect 56928 5720 56934 5732
rect 56965 5729 56977 5732
rect 57011 5729 57023 5763
rect 56965 5723 57023 5729
rect 56140 5704 56192 5710
rect 37645 5695 37703 5701
rect 37645 5661 37657 5695
rect 37691 5661 37703 5695
rect 37826 5692 37832 5704
rect 37787 5664 37832 5692
rect 37645 5655 37703 5661
rect 37826 5652 37832 5664
rect 37884 5652 37890 5704
rect 40034 5692 40040 5704
rect 39947 5664 40040 5692
rect 40034 5652 40040 5664
rect 40092 5652 40098 5704
rect 40218 5652 40224 5704
rect 40276 5692 40282 5704
rect 40313 5695 40371 5701
rect 40313 5692 40325 5695
rect 40276 5664 40325 5692
rect 40276 5652 40282 5664
rect 40313 5661 40325 5664
rect 40359 5692 40371 5695
rect 40957 5695 41015 5701
rect 40957 5692 40969 5695
rect 40359 5664 40969 5692
rect 40359 5661 40371 5664
rect 40313 5655 40371 5661
rect 40957 5661 40969 5664
rect 41003 5661 41015 5695
rect 43530 5692 43536 5704
rect 43491 5664 43536 5692
rect 40957 5655 41015 5661
rect 43530 5652 43536 5664
rect 43588 5652 43594 5704
rect 53558 5652 53564 5704
rect 53616 5692 53622 5704
rect 54113 5695 54171 5701
rect 54113 5692 54125 5695
rect 53616 5664 54125 5692
rect 53616 5652 53622 5664
rect 54113 5661 54125 5664
rect 54159 5661 54171 5695
rect 54113 5655 54171 5661
rect 55766 5652 55772 5704
rect 55824 5692 55830 5704
rect 56045 5695 56103 5701
rect 56045 5692 56057 5695
rect 55824 5664 56057 5692
rect 55824 5652 55830 5664
rect 56045 5661 56057 5664
rect 56091 5661 56103 5695
rect 56045 5655 56103 5661
rect 40052 5624 40080 5652
rect 56140 5646 56192 5652
rect 41233 5627 41291 5633
rect 41233 5624 41245 5627
rect 36832 5596 41245 5624
rect 35437 5587 35495 5593
rect 41233 5593 41245 5596
rect 41279 5593 41291 5627
rect 41233 5587 41291 5593
rect 31220 5528 31524 5556
rect 31570 5516 31576 5568
rect 31628 5556 31634 5568
rect 32398 5556 32404 5568
rect 31628 5528 31673 5556
rect 32359 5528 32404 5556
rect 31628 5516 31634 5528
rect 32398 5516 32404 5528
rect 32456 5516 32462 5568
rect 33226 5556 33232 5568
rect 33187 5528 33232 5556
rect 33226 5516 33232 5528
rect 33284 5516 33290 5568
rect 35452 5556 35480 5587
rect 35894 5556 35900 5568
rect 35452 5528 35900 5556
rect 35894 5516 35900 5528
rect 35952 5556 35958 5568
rect 37090 5556 37096 5568
rect 35952 5528 37096 5556
rect 35952 5516 35958 5528
rect 37090 5516 37096 5528
rect 37148 5516 37154 5568
rect 37737 5559 37795 5565
rect 37737 5525 37749 5559
rect 37783 5556 37795 5559
rect 37826 5556 37832 5568
rect 37783 5528 37832 5556
rect 37783 5525 37795 5528
rect 37737 5519 37795 5525
rect 37826 5516 37832 5528
rect 37884 5516 37890 5568
rect 40494 5556 40500 5568
rect 40455 5528 40500 5556
rect 40494 5516 40500 5528
rect 40552 5516 40558 5568
rect 40862 5516 40868 5568
rect 40920 5556 40926 5568
rect 40957 5559 41015 5565
rect 40957 5556 40969 5559
rect 40920 5528 40969 5556
rect 40920 5516 40926 5528
rect 40957 5525 40969 5528
rect 41003 5525 41015 5559
rect 40957 5519 41015 5525
rect 43901 5559 43959 5565
rect 43901 5525 43913 5559
rect 43947 5556 43959 5559
rect 44174 5556 44180 5568
rect 43947 5528 44180 5556
rect 43947 5525 43959 5528
rect 43901 5519 43959 5525
rect 44174 5516 44180 5528
rect 44232 5516 44238 5568
rect 53558 5556 53564 5568
rect 53519 5528 53564 5556
rect 53558 5516 53564 5528
rect 53616 5516 53622 5568
rect 1104 5466 58880 5488
rect 1104 5414 19574 5466
rect 19626 5414 19638 5466
rect 19690 5414 19702 5466
rect 19754 5414 19766 5466
rect 19818 5414 19830 5466
rect 19882 5414 50294 5466
rect 50346 5414 50358 5466
rect 50410 5414 50422 5466
rect 50474 5414 50486 5466
rect 50538 5414 50550 5466
rect 50602 5414 58880 5466
rect 1104 5392 58880 5414
rect 3145 5355 3203 5361
rect 3145 5321 3157 5355
rect 3191 5352 3203 5355
rect 3418 5352 3424 5364
rect 3191 5324 3424 5352
rect 3191 5321 3203 5324
rect 3145 5315 3203 5321
rect 3418 5312 3424 5324
rect 3476 5312 3482 5364
rect 9674 5312 9680 5364
rect 9732 5352 9738 5364
rect 13265 5355 13323 5361
rect 13265 5352 13277 5355
rect 9732 5324 13277 5352
rect 9732 5312 9738 5324
rect 13265 5321 13277 5324
rect 13311 5321 13323 5355
rect 22557 5355 22615 5361
rect 22557 5352 22569 5355
rect 13265 5315 13323 5321
rect 22066 5324 22569 5352
rect 3050 5244 3056 5296
rect 3108 5284 3114 5296
rect 4065 5287 4123 5293
rect 4065 5284 4077 5287
rect 3108 5256 4077 5284
rect 3108 5244 3114 5256
rect 4065 5253 4077 5256
rect 4111 5253 4123 5287
rect 4065 5247 4123 5253
rect 6730 5244 6736 5296
rect 6788 5284 6794 5296
rect 6825 5287 6883 5293
rect 6825 5284 6837 5287
rect 6788 5256 6837 5284
rect 6788 5244 6794 5256
rect 6825 5253 6837 5256
rect 6871 5253 6883 5287
rect 6825 5247 6883 5253
rect 19334 5244 19340 5296
rect 19392 5284 19398 5296
rect 19978 5293 19984 5296
rect 19705 5287 19763 5293
rect 19705 5284 19717 5287
rect 19392 5256 19717 5284
rect 19392 5244 19398 5256
rect 19705 5253 19717 5256
rect 19751 5253 19763 5287
rect 19705 5247 19763 5253
rect 19921 5287 19984 5293
rect 19921 5253 19933 5287
rect 19967 5253 19984 5287
rect 19921 5247 19984 5253
rect 19978 5244 19984 5247
rect 20036 5244 20042 5296
rect 2961 5219 3019 5225
rect 2961 5185 2973 5219
rect 3007 5185 3019 5219
rect 3234 5216 3240 5228
rect 3195 5188 3240 5216
rect 2961 5179 3019 5185
rect 2976 5148 3004 5179
rect 3234 5176 3240 5188
rect 3292 5176 3298 5228
rect 3697 5219 3755 5225
rect 3697 5185 3709 5219
rect 3743 5185 3755 5219
rect 3697 5179 3755 5185
rect 3712 5148 3740 5179
rect 3786 5176 3792 5228
rect 3844 5216 3850 5228
rect 3970 5216 3976 5228
rect 3844 5188 3889 5216
rect 3931 5188 3976 5216
rect 3844 5176 3850 5188
rect 3970 5176 3976 5188
rect 4028 5176 4034 5228
rect 4203 5219 4261 5225
rect 4203 5185 4215 5219
rect 4249 5216 4261 5219
rect 6454 5216 6460 5228
rect 4249 5188 6460 5216
rect 4249 5185 4261 5188
rect 4203 5179 4261 5185
rect 6454 5176 6460 5188
rect 6512 5176 6518 5228
rect 7282 5176 7288 5228
rect 7340 5216 7346 5228
rect 9309 5219 9367 5225
rect 9309 5216 9321 5219
rect 7340 5188 9321 5216
rect 7340 5176 7346 5188
rect 9309 5185 9321 5188
rect 9355 5185 9367 5219
rect 9309 5179 9367 5185
rect 9493 5219 9551 5225
rect 9493 5185 9505 5219
rect 9539 5216 9551 5219
rect 10042 5216 10048 5228
rect 9539 5188 10048 5216
rect 9539 5185 9551 5188
rect 9493 5179 9551 5185
rect 10042 5176 10048 5188
rect 10100 5176 10106 5228
rect 13446 5216 13452 5228
rect 13407 5188 13452 5216
rect 13446 5176 13452 5188
rect 13504 5176 13510 5228
rect 13633 5219 13691 5225
rect 13633 5185 13645 5219
rect 13679 5216 13691 5219
rect 14458 5216 14464 5228
rect 13679 5188 14464 5216
rect 13679 5185 13691 5188
rect 13633 5179 13691 5185
rect 14458 5176 14464 5188
rect 14516 5176 14522 5228
rect 16853 5219 16911 5225
rect 16853 5185 16865 5219
rect 16899 5216 16911 5219
rect 17589 5219 17647 5225
rect 17589 5216 17601 5219
rect 16899 5188 17601 5216
rect 16899 5185 16911 5188
rect 16853 5179 16911 5185
rect 17589 5185 17601 5188
rect 17635 5216 17647 5219
rect 22066 5216 22094 5324
rect 22557 5321 22569 5324
rect 22603 5321 22615 5355
rect 22557 5315 22615 5321
rect 26970 5312 26976 5364
rect 27028 5352 27034 5364
rect 27341 5355 27399 5361
rect 27341 5352 27353 5355
rect 27028 5324 27353 5352
rect 27028 5312 27034 5324
rect 27341 5321 27353 5324
rect 27387 5321 27399 5355
rect 56321 5355 56379 5361
rect 27341 5315 27399 5321
rect 27448 5324 41414 5352
rect 23474 5244 23480 5296
rect 23532 5284 23538 5296
rect 24121 5287 24179 5293
rect 24121 5284 24133 5287
rect 23532 5256 24133 5284
rect 23532 5244 23538 5256
rect 24121 5253 24133 5256
rect 24167 5284 24179 5287
rect 24578 5284 24584 5296
rect 24167 5256 24584 5284
rect 24167 5253 24179 5256
rect 24121 5247 24179 5253
rect 24578 5244 24584 5256
rect 24636 5244 24642 5296
rect 26142 5244 26148 5296
rect 26200 5284 26206 5296
rect 27448 5284 27476 5324
rect 31570 5284 31576 5296
rect 26200 5256 27476 5284
rect 27724 5256 31576 5284
rect 26200 5244 26206 5256
rect 17635 5188 22094 5216
rect 22925 5219 22983 5225
rect 17635 5185 17647 5188
rect 17589 5179 17647 5185
rect 22925 5185 22937 5219
rect 22971 5216 22983 5219
rect 23382 5216 23388 5228
rect 22971 5188 23388 5216
rect 22971 5185 22983 5188
rect 22925 5179 22983 5185
rect 23382 5176 23388 5188
rect 23440 5176 23446 5228
rect 23937 5219 23995 5225
rect 23937 5185 23949 5219
rect 23983 5185 23995 5219
rect 23937 5179 23995 5185
rect 6638 5148 6644 5160
rect 2976 5120 6644 5148
rect 6638 5108 6644 5120
rect 6696 5108 6702 5160
rect 17129 5151 17187 5157
rect 17129 5117 17141 5151
rect 17175 5148 17187 5151
rect 17865 5151 17923 5157
rect 17865 5148 17877 5151
rect 17175 5120 17877 5148
rect 17175 5117 17187 5120
rect 17129 5111 17187 5117
rect 17865 5117 17877 5120
rect 17911 5148 17923 5151
rect 20162 5148 20168 5160
rect 17911 5120 20168 5148
rect 17911 5117 17923 5120
rect 17865 5111 17923 5117
rect 20162 5108 20168 5120
rect 20220 5108 20226 5160
rect 23017 5151 23075 5157
rect 23017 5117 23029 5151
rect 23063 5148 23075 5151
rect 23952 5148 23980 5179
rect 24026 5176 24032 5228
rect 24084 5216 24090 5228
rect 24259 5219 24317 5225
rect 24084 5188 24129 5216
rect 24084 5176 24090 5188
rect 24259 5185 24271 5219
rect 24305 5216 24317 5219
rect 25225 5219 25283 5225
rect 24305 5188 25176 5216
rect 24305 5185 24317 5188
rect 24259 5179 24317 5185
rect 23063 5120 23980 5148
rect 23063 5117 23075 5120
rect 23017 5111 23075 5117
rect 4341 5083 4399 5089
rect 4341 5049 4353 5083
rect 4387 5080 4399 5083
rect 6549 5083 6607 5089
rect 4387 5052 6500 5080
rect 4387 5049 4399 5052
rect 4341 5043 4399 5049
rect 6270 4972 6276 5024
rect 6328 5012 6334 5024
rect 6365 5015 6423 5021
rect 6365 5012 6377 5015
rect 6328 4984 6377 5012
rect 6328 4972 6334 4984
rect 6365 4981 6377 4984
rect 6411 4981 6423 5015
rect 6472 5012 6500 5052
rect 6549 5049 6561 5083
rect 6595 5080 6607 5083
rect 6822 5080 6828 5092
rect 6595 5052 6828 5080
rect 6595 5049 6607 5052
rect 6549 5043 6607 5049
rect 6822 5040 6828 5052
rect 6880 5040 6886 5092
rect 9674 5080 9680 5092
rect 9416 5052 9680 5080
rect 9416 5012 9444 5052
rect 9674 5040 9680 5052
rect 9732 5040 9738 5092
rect 16574 5040 16580 5092
rect 16632 5080 16638 5092
rect 17037 5083 17095 5089
rect 17037 5080 17049 5083
rect 16632 5052 17049 5080
rect 16632 5040 16638 5052
rect 17037 5049 17049 5052
rect 17083 5080 17095 5083
rect 17678 5080 17684 5092
rect 17083 5052 17684 5080
rect 17083 5049 17095 5052
rect 17037 5043 17095 5049
rect 17678 5040 17684 5052
rect 17736 5040 17742 5092
rect 23952 5080 23980 5120
rect 24397 5151 24455 5157
rect 24397 5117 24409 5151
rect 24443 5148 24455 5151
rect 25148 5148 25176 5188
rect 25225 5185 25237 5219
rect 25271 5216 25283 5219
rect 27430 5216 27436 5228
rect 25271 5188 27436 5216
rect 25271 5185 25283 5188
rect 25225 5179 25283 5185
rect 25314 5148 25320 5160
rect 24443 5120 25084 5148
rect 25148 5120 25320 5148
rect 24443 5117 24455 5120
rect 24397 5111 24455 5117
rect 24857 5083 24915 5089
rect 24857 5080 24869 5083
rect 23952 5052 24869 5080
rect 24857 5049 24869 5052
rect 24903 5049 24915 5083
rect 25056 5080 25084 5120
rect 25314 5108 25320 5120
rect 25372 5108 25378 5160
rect 25424 5080 25452 5188
rect 27430 5176 27436 5188
rect 27488 5176 27494 5228
rect 27724 5225 27752 5256
rect 31570 5244 31576 5256
rect 31628 5284 31634 5296
rect 33134 5284 33140 5296
rect 31628 5256 33140 5284
rect 31628 5244 31634 5256
rect 33134 5244 33140 5256
rect 33192 5244 33198 5296
rect 41386 5284 41414 5324
rect 56321 5321 56333 5355
rect 56367 5352 56379 5355
rect 56686 5352 56692 5364
rect 56367 5324 56692 5352
rect 56367 5321 56379 5324
rect 56321 5315 56379 5321
rect 56686 5312 56692 5324
rect 56744 5312 56750 5364
rect 57698 5284 57704 5296
rect 41386 5256 57704 5284
rect 57698 5244 57704 5256
rect 57756 5244 57762 5296
rect 33232 5228 33284 5234
rect 27709 5219 27767 5225
rect 27709 5185 27721 5219
rect 27755 5185 27767 5219
rect 27709 5179 27767 5185
rect 30466 5176 30472 5228
rect 30524 5216 30530 5228
rect 31205 5219 31263 5225
rect 31205 5216 31217 5219
rect 30524 5188 31217 5216
rect 30524 5176 30530 5188
rect 31205 5185 31217 5188
rect 31251 5185 31263 5219
rect 31205 5179 31263 5185
rect 31389 5219 31447 5225
rect 31389 5185 31401 5219
rect 31435 5216 31447 5219
rect 32398 5216 32404 5228
rect 31435 5188 32404 5216
rect 31435 5185 31447 5188
rect 31389 5179 31447 5185
rect 27614 5148 27620 5160
rect 27575 5120 27620 5148
rect 27614 5108 27620 5120
rect 27672 5108 27678 5160
rect 31220 5148 31248 5179
rect 32398 5176 32404 5188
rect 32456 5176 32462 5228
rect 33873 5219 33931 5225
rect 33873 5185 33885 5219
rect 33919 5216 33931 5219
rect 35894 5216 35900 5228
rect 33919 5188 35900 5216
rect 33919 5185 33931 5188
rect 33873 5179 33931 5185
rect 35894 5176 35900 5188
rect 35952 5176 35958 5228
rect 40494 5176 40500 5228
rect 40552 5216 40558 5228
rect 40681 5219 40739 5225
rect 40681 5216 40693 5219
rect 40552 5188 40693 5216
rect 40552 5176 40558 5188
rect 40681 5185 40693 5188
rect 40727 5185 40739 5219
rect 40862 5216 40868 5228
rect 40823 5188 40868 5216
rect 40681 5179 40739 5185
rect 33232 5170 33284 5176
rect 32214 5148 32220 5160
rect 31220 5120 32220 5148
rect 32214 5108 32220 5120
rect 32272 5108 32278 5160
rect 32858 5148 32864 5160
rect 32819 5120 32864 5148
rect 32858 5108 32864 5120
rect 32916 5108 32922 5160
rect 40696 5148 40724 5179
rect 40862 5176 40868 5188
rect 40920 5176 40926 5228
rect 44174 5216 44180 5228
rect 44135 5188 44180 5216
rect 44174 5176 44180 5188
rect 44232 5176 44238 5228
rect 44266 5176 44272 5228
rect 44324 5216 44330 5228
rect 44450 5216 44456 5228
rect 44324 5188 44369 5216
rect 44411 5188 44456 5216
rect 44324 5176 44330 5188
rect 44450 5176 44456 5188
rect 44508 5176 44514 5228
rect 45186 5216 45192 5228
rect 45147 5188 45192 5216
rect 45186 5176 45192 5188
rect 45244 5176 45250 5228
rect 56870 5176 56876 5228
rect 56928 5216 56934 5228
rect 56965 5219 57023 5225
rect 56965 5216 56977 5219
rect 56928 5188 56977 5216
rect 56928 5176 56934 5188
rect 56965 5185 56977 5188
rect 57011 5185 57023 5219
rect 56965 5179 57023 5185
rect 41230 5148 41236 5160
rect 40696 5120 41236 5148
rect 41230 5108 41236 5120
rect 41288 5108 41294 5160
rect 25056 5052 25452 5080
rect 24857 5043 24915 5049
rect 38654 5040 38660 5092
rect 38712 5080 38718 5092
rect 40494 5080 40500 5092
rect 38712 5052 40500 5080
rect 38712 5040 38718 5052
rect 40494 5040 40500 5052
rect 40552 5040 40558 5092
rect 44192 5080 44220 5176
rect 44358 5148 44364 5160
rect 44319 5120 44364 5148
rect 44358 5108 44364 5120
rect 44416 5108 44422 5160
rect 45097 5151 45155 5157
rect 45097 5117 45109 5151
rect 45143 5117 45155 5151
rect 45097 5111 45155 5117
rect 45112 5080 45140 5111
rect 56686 5108 56692 5160
rect 56744 5148 56750 5160
rect 57057 5151 57115 5157
rect 57057 5148 57069 5151
rect 56744 5120 57069 5148
rect 56744 5108 56750 5120
rect 57057 5117 57069 5120
rect 57103 5117 57115 5151
rect 57057 5111 57115 5117
rect 45554 5080 45560 5092
rect 44192 5052 45140 5080
rect 45515 5052 45560 5080
rect 45554 5040 45560 5052
rect 45612 5040 45618 5092
rect 6472 4984 9444 5012
rect 9493 5015 9551 5021
rect 6365 4975 6423 4981
rect 9493 4981 9505 5015
rect 9539 5012 9551 5015
rect 10318 5012 10324 5024
rect 9539 4984 10324 5012
rect 9539 4981 9551 4984
rect 9493 4975 9551 4981
rect 10318 4972 10324 4984
rect 10376 4972 10382 5024
rect 16666 5012 16672 5024
rect 16627 4984 16672 5012
rect 16666 4972 16672 4984
rect 16724 4972 16730 5024
rect 17586 5012 17592 5024
rect 17547 4984 17592 5012
rect 17586 4972 17592 4984
rect 17644 4972 17650 5024
rect 19426 4972 19432 5024
rect 19484 5012 19490 5024
rect 19886 5012 19892 5024
rect 19484 4984 19892 5012
rect 19484 4972 19490 4984
rect 19886 4972 19892 4984
rect 19944 4972 19950 5024
rect 20070 5012 20076 5024
rect 20031 4984 20076 5012
rect 20070 4972 20076 4984
rect 20128 4972 20134 5024
rect 23750 5012 23756 5024
rect 23711 4984 23756 5012
rect 23750 4972 23756 4984
rect 23808 4972 23814 5024
rect 31570 5012 31576 5024
rect 31531 4984 31576 5012
rect 31570 4972 31576 4984
rect 31628 4972 31634 5024
rect 40865 5015 40923 5021
rect 40865 4981 40877 5015
rect 40911 5012 40923 5015
rect 41506 5012 41512 5024
rect 40911 4984 41512 5012
rect 40911 4981 40923 4984
rect 40865 4975 40923 4981
rect 41506 4972 41512 4984
rect 41564 4972 41570 5024
rect 43806 4972 43812 5024
rect 43864 5012 43870 5024
rect 43993 5015 44051 5021
rect 43993 5012 44005 5015
rect 43864 4984 44005 5012
rect 43864 4972 43870 4984
rect 43993 4981 44005 4984
rect 44039 4981 44051 5015
rect 54570 5012 54576 5024
rect 54531 4984 54576 5012
rect 43993 4975 44051 4981
rect 54570 4972 54576 4984
rect 54628 5012 54634 5024
rect 55766 5012 55772 5024
rect 54628 4984 55772 5012
rect 54628 4972 54634 4984
rect 55766 4972 55772 4984
rect 55824 4972 55830 5024
rect 57333 5015 57391 5021
rect 57333 4981 57345 5015
rect 57379 5012 57391 5015
rect 57882 5012 57888 5024
rect 57379 4984 57888 5012
rect 57379 4981 57391 4984
rect 57333 4975 57391 4981
rect 57882 4972 57888 4984
rect 57940 4972 57946 5024
rect 1104 4922 58880 4944
rect 1104 4870 4214 4922
rect 4266 4870 4278 4922
rect 4330 4870 4342 4922
rect 4394 4870 4406 4922
rect 4458 4870 4470 4922
rect 4522 4870 34934 4922
rect 34986 4870 34998 4922
rect 35050 4870 35062 4922
rect 35114 4870 35126 4922
rect 35178 4870 35190 4922
rect 35242 4870 58880 4922
rect 1104 4848 58880 4870
rect 3970 4808 3976 4820
rect 3931 4780 3976 4808
rect 3970 4768 3976 4780
rect 4028 4768 4034 4820
rect 6638 4808 6644 4820
rect 6551 4780 6644 4808
rect 6638 4768 6644 4780
rect 6696 4808 6702 4820
rect 7098 4808 7104 4820
rect 6696 4780 7104 4808
rect 6696 4768 6702 4780
rect 7098 4768 7104 4780
rect 7156 4768 7162 4820
rect 7282 4808 7288 4820
rect 7243 4780 7288 4808
rect 7282 4768 7288 4780
rect 7340 4768 7346 4820
rect 15838 4808 15844 4820
rect 10060 4780 15844 4808
rect 2225 4743 2283 4749
rect 2225 4709 2237 4743
rect 2271 4709 2283 4743
rect 2225 4703 2283 4709
rect 1673 4607 1731 4613
rect 1673 4573 1685 4607
rect 1719 4604 1731 4607
rect 2240 4604 2268 4703
rect 3234 4700 3240 4752
rect 3292 4740 3298 4752
rect 7300 4740 7328 4768
rect 3292 4712 7328 4740
rect 3292 4700 3298 4712
rect 1719 4576 2268 4604
rect 2409 4607 2467 4613
rect 1719 4573 1731 4576
rect 1673 4567 1731 4573
rect 2409 4573 2421 4607
rect 2455 4604 2467 4607
rect 3789 4607 3847 4613
rect 2455 4576 3004 4604
rect 2455 4573 2467 4576
rect 2409 4567 2467 4573
rect 2976 4545 3004 4576
rect 3789 4573 3801 4607
rect 3835 4604 3847 4607
rect 3878 4604 3884 4616
rect 3835 4576 3884 4604
rect 3835 4573 3847 4576
rect 3789 4567 3847 4573
rect 3878 4564 3884 4576
rect 3936 4564 3942 4616
rect 3988 4613 4016 4712
rect 6270 4672 6276 4684
rect 6231 4644 6276 4672
rect 6270 4632 6276 4644
rect 6328 4632 6334 4684
rect 7374 4632 7380 4684
rect 7432 4672 7438 4684
rect 10060 4681 10088 4780
rect 15838 4768 15844 4780
rect 15896 4768 15902 4820
rect 16022 4768 16028 4820
rect 16080 4808 16086 4820
rect 16209 4811 16267 4817
rect 16209 4808 16221 4811
rect 16080 4780 16221 4808
rect 16080 4768 16086 4780
rect 16209 4777 16221 4780
rect 16255 4777 16267 4811
rect 16209 4771 16267 4777
rect 17954 4768 17960 4820
rect 18012 4808 18018 4820
rect 19429 4811 19487 4817
rect 19429 4808 19441 4811
rect 18012 4780 19441 4808
rect 18012 4768 18018 4780
rect 19429 4777 19441 4780
rect 19475 4777 19487 4811
rect 19429 4771 19487 4777
rect 19886 4768 19892 4820
rect 19944 4808 19950 4820
rect 27065 4811 27123 4817
rect 27065 4808 27077 4811
rect 19944 4780 27077 4808
rect 19944 4768 19950 4780
rect 27065 4777 27077 4780
rect 27111 4777 27123 4811
rect 27065 4771 27123 4777
rect 33134 4768 33140 4820
rect 33192 4808 33198 4820
rect 33597 4811 33655 4817
rect 33597 4808 33609 4811
rect 33192 4780 33609 4808
rect 33192 4768 33198 4780
rect 33597 4777 33609 4780
rect 33643 4777 33655 4811
rect 33597 4771 33655 4777
rect 37642 4768 37648 4820
rect 37700 4808 37706 4820
rect 38102 4808 38108 4820
rect 37700 4780 38108 4808
rect 37700 4768 37706 4780
rect 38102 4768 38108 4780
rect 38160 4808 38166 4820
rect 44358 4808 44364 4820
rect 38160 4780 44364 4808
rect 38160 4768 38166 4780
rect 44358 4768 44364 4780
rect 44416 4768 44422 4820
rect 45097 4811 45155 4817
rect 45097 4777 45109 4811
rect 45143 4808 45155 4811
rect 45186 4808 45192 4820
rect 45143 4780 45192 4808
rect 45143 4777 45155 4780
rect 45097 4771 45155 4777
rect 45186 4768 45192 4780
rect 45244 4768 45250 4820
rect 53558 4740 53564 4752
rect 10152 4712 53564 4740
rect 10045 4675 10103 4681
rect 7432 4644 9904 4672
rect 7432 4632 7438 4644
rect 7185 4617 7243 4623
rect 3973 4607 4031 4613
rect 3973 4573 3985 4607
rect 4019 4573 4031 4607
rect 6454 4604 6460 4616
rect 6415 4576 6460 4604
rect 3973 4567 4031 4573
rect 6454 4564 6460 4576
rect 6512 4564 6518 4616
rect 6730 4564 6736 4616
rect 6788 4604 6794 4616
rect 7185 4614 7197 4617
rect 7024 4604 7197 4614
rect 6788 4586 7197 4604
rect 6788 4576 7052 4586
rect 7185 4583 7197 4586
rect 7231 4583 7243 4617
rect 7185 4577 7243 4583
rect 6788 4564 6794 4576
rect 7282 4564 7288 4616
rect 7340 4604 7346 4616
rect 9769 4607 9827 4613
rect 9769 4604 9781 4607
rect 7340 4576 9781 4604
rect 7340 4564 7346 4576
rect 9769 4573 9781 4576
rect 9815 4573 9827 4607
rect 9876 4604 9904 4644
rect 10045 4641 10057 4675
rect 10091 4641 10103 4675
rect 10045 4635 10103 4641
rect 10152 4604 10180 4712
rect 53558 4700 53564 4712
rect 53616 4700 53622 4752
rect 10226 4632 10232 4684
rect 10284 4672 10290 4684
rect 10284 4644 10329 4672
rect 12406 4644 22094 4672
rect 10284 4632 10290 4644
rect 10318 4604 10324 4616
rect 9876 4576 10180 4604
rect 10279 4576 10324 4604
rect 9769 4567 9827 4573
rect 10318 4564 10324 4576
rect 10376 4564 10382 4616
rect 11054 4604 11060 4616
rect 11015 4576 11060 4604
rect 11054 4564 11060 4576
rect 11112 4564 11118 4616
rect 2961 4539 3019 4545
rect 2961 4505 2973 4539
rect 3007 4536 3019 4539
rect 12406 4536 12434 4644
rect 16025 4607 16083 4613
rect 16025 4573 16037 4607
rect 16071 4573 16083 4607
rect 16025 4567 16083 4573
rect 16209 4607 16267 4613
rect 16209 4573 16221 4607
rect 16255 4604 16267 4607
rect 17586 4604 17592 4616
rect 16255 4576 17592 4604
rect 16255 4573 16267 4576
rect 16209 4567 16267 4573
rect 3007 4508 6684 4536
rect 3007 4505 3019 4508
rect 2961 4499 3019 4505
rect 1486 4468 1492 4480
rect 1447 4440 1492 4468
rect 1486 4428 1492 4440
rect 1544 4428 1550 4480
rect 6656 4468 6684 4508
rect 9876 4508 12434 4536
rect 16040 4536 16068 4567
rect 17586 4564 17592 4576
rect 17644 4564 17650 4616
rect 19797 4607 19855 4613
rect 19797 4573 19809 4607
rect 19843 4604 19855 4607
rect 20070 4604 20076 4616
rect 19843 4576 20076 4604
rect 19843 4573 19855 4576
rect 19797 4567 19855 4573
rect 20070 4564 20076 4576
rect 20128 4564 20134 4616
rect 22066 4604 22094 4644
rect 23382 4632 23388 4684
rect 23440 4672 23446 4684
rect 24397 4675 24455 4681
rect 24397 4672 24409 4675
rect 23440 4644 24409 4672
rect 23440 4632 23446 4644
rect 24397 4641 24409 4644
rect 24443 4641 24455 4675
rect 26694 4672 26700 4684
rect 24397 4635 24455 4641
rect 24504 4644 26700 4672
rect 24504 4604 24532 4644
rect 26694 4632 26700 4644
rect 26752 4632 26758 4684
rect 26970 4632 26976 4684
rect 27028 4672 27034 4684
rect 27249 4675 27307 4681
rect 27249 4672 27261 4675
rect 27028 4644 27261 4672
rect 27028 4632 27034 4644
rect 27249 4641 27261 4644
rect 27295 4641 27307 4675
rect 27249 4635 27307 4641
rect 27430 4632 27436 4684
rect 27488 4672 27494 4684
rect 29733 4675 29791 4681
rect 29733 4672 29745 4675
rect 27488 4644 29745 4672
rect 27488 4632 27494 4644
rect 29733 4641 29745 4644
rect 29779 4641 29791 4675
rect 29733 4635 29791 4641
rect 37274 4632 37280 4684
rect 37332 4672 37338 4684
rect 37737 4675 37795 4681
rect 37737 4672 37749 4675
rect 37332 4644 37749 4672
rect 37332 4632 37338 4644
rect 37737 4641 37749 4644
rect 37783 4672 37795 4675
rect 40313 4675 40371 4681
rect 40313 4672 40325 4675
rect 37783 4644 40325 4672
rect 37783 4641 37795 4644
rect 37737 4635 37795 4641
rect 40313 4641 40325 4644
rect 40359 4641 40371 4675
rect 44266 4672 44272 4684
rect 40313 4635 40371 4641
rect 40696 4644 44272 4672
rect 40696 4616 40724 4644
rect 44266 4632 44272 4644
rect 44324 4672 44330 4684
rect 46201 4675 46259 4681
rect 44324 4644 44956 4672
rect 44324 4632 44330 4644
rect 22066 4576 24532 4604
rect 24581 4607 24639 4613
rect 24581 4573 24593 4607
rect 24627 4604 24639 4607
rect 24762 4604 24768 4616
rect 24627 4576 24768 4604
rect 24627 4573 24639 4576
rect 24581 4567 24639 4573
rect 24762 4564 24768 4576
rect 24820 4564 24826 4616
rect 27341 4607 27399 4613
rect 27341 4573 27353 4607
rect 27387 4573 27399 4607
rect 30745 4607 30803 4613
rect 27341 4567 27399 4573
rect 16666 4536 16672 4548
rect 16040 4508 16672 4536
rect 9876 4468 9904 4508
rect 16666 4496 16672 4508
rect 16724 4496 16730 4548
rect 19613 4539 19671 4545
rect 19613 4505 19625 4539
rect 19659 4536 19671 4539
rect 20162 4536 20168 4548
rect 19659 4508 20168 4536
rect 19659 4505 19671 4508
rect 19613 4499 19671 4505
rect 20162 4496 20168 4508
rect 20220 4496 20226 4548
rect 26878 4536 26884 4548
rect 24780 4508 26884 4536
rect 11146 4468 11152 4480
rect 6656 4440 9904 4468
rect 11107 4440 11152 4468
rect 11146 4428 11152 4440
rect 11204 4428 11210 4480
rect 12710 4428 12716 4480
rect 12768 4468 12774 4480
rect 16942 4468 16948 4480
rect 12768 4440 16948 4468
rect 12768 4428 12774 4440
rect 16942 4428 16948 4440
rect 17000 4428 17006 4480
rect 24780 4477 24808 4508
rect 26878 4496 26884 4508
rect 26936 4536 26942 4548
rect 27356 4536 27384 4567
rect 26936 4508 27384 4536
rect 30668 4536 30696 4590
rect 30745 4573 30757 4607
rect 30791 4604 30803 4607
rect 31570 4604 31576 4616
rect 30791 4576 31576 4604
rect 30791 4573 30803 4576
rect 30745 4567 30803 4573
rect 31570 4564 31576 4576
rect 31628 4604 31634 4616
rect 33170 4607 33228 4613
rect 33170 4604 33182 4607
rect 31628 4576 33182 4604
rect 31628 4564 31634 4576
rect 33170 4573 33182 4576
rect 33216 4573 33228 4607
rect 33170 4567 33228 4573
rect 33689 4607 33747 4613
rect 33689 4573 33701 4607
rect 33735 4604 33747 4607
rect 36725 4607 36783 4613
rect 36725 4604 36737 4607
rect 33735 4576 36737 4604
rect 33735 4573 33747 4576
rect 33689 4567 33747 4573
rect 36725 4573 36737 4576
rect 36771 4604 36783 4607
rect 37550 4604 37556 4616
rect 36771 4576 37556 4604
rect 36771 4573 36783 4576
rect 36725 4567 36783 4573
rect 37550 4564 37556 4576
rect 37608 4564 37614 4616
rect 37642 4564 37648 4616
rect 37700 4604 37706 4616
rect 37700 4576 37745 4604
rect 37700 4564 37706 4576
rect 37826 4564 37832 4616
rect 37884 4604 37890 4616
rect 40402 4604 40408 4616
rect 37884 4576 37929 4604
rect 40363 4576 40408 4604
rect 37884 4564 37890 4576
rect 40402 4564 40408 4576
rect 40460 4604 40466 4616
rect 40678 4604 40684 4616
rect 40460 4576 40684 4604
rect 40460 4564 40466 4576
rect 40678 4564 40684 4576
rect 40736 4564 40742 4616
rect 41322 4604 41328 4616
rect 40788 4576 41328 4604
rect 32858 4536 32864 4548
rect 30668 4508 32864 4536
rect 26936 4496 26942 4508
rect 32858 4496 32864 4508
rect 32916 4536 32922 4548
rect 36909 4539 36967 4545
rect 32916 4508 33272 4536
rect 32916 4496 32922 4508
rect 24765 4471 24823 4477
rect 24765 4437 24777 4471
rect 24811 4437 24823 4471
rect 24765 4431 24823 4437
rect 33045 4471 33103 4477
rect 33045 4437 33057 4471
rect 33091 4468 33103 4471
rect 33134 4468 33140 4480
rect 33091 4440 33140 4468
rect 33091 4437 33103 4440
rect 33045 4431 33103 4437
rect 33134 4428 33140 4440
rect 33192 4428 33198 4480
rect 33244 4477 33272 4508
rect 36909 4505 36921 4539
rect 36955 4505 36967 4539
rect 37090 4536 37096 4548
rect 37051 4508 37096 4536
rect 36909 4499 36967 4505
rect 33229 4471 33287 4477
rect 33229 4437 33241 4471
rect 33275 4437 33287 4471
rect 36924 4468 36952 4499
rect 37090 4496 37096 4508
rect 37148 4496 37154 4548
rect 37660 4468 37688 4564
rect 40788 4477 40816 4576
rect 41322 4564 41328 4576
rect 41380 4604 41386 4616
rect 41417 4607 41475 4613
rect 41417 4604 41429 4607
rect 41380 4576 41429 4604
rect 41380 4564 41386 4576
rect 41417 4573 41429 4576
rect 41463 4573 41475 4607
rect 41417 4567 41475 4573
rect 41506 4564 41512 4616
rect 41564 4604 41570 4616
rect 44928 4604 44956 4644
rect 46201 4641 46213 4675
rect 46247 4672 46259 4675
rect 46290 4672 46296 4684
rect 46247 4644 46296 4672
rect 46247 4641 46259 4644
rect 46201 4635 46259 4641
rect 46290 4632 46296 4644
rect 46348 4632 46354 4684
rect 46382 4632 46388 4684
rect 46440 4672 46446 4684
rect 46477 4675 46535 4681
rect 46477 4672 46489 4675
rect 46440 4644 46489 4672
rect 46440 4632 46446 4644
rect 46477 4641 46489 4644
rect 46523 4641 46535 4675
rect 46477 4635 46535 4641
rect 45005 4607 45063 4613
rect 45005 4604 45017 4607
rect 41564 4576 41609 4604
rect 44928 4576 45017 4604
rect 41564 4564 41570 4576
rect 45005 4573 45017 4576
rect 45051 4573 45063 4607
rect 45005 4567 45063 4573
rect 45189 4607 45247 4613
rect 45189 4573 45201 4607
rect 45235 4573 45247 4607
rect 45189 4567 45247 4573
rect 44358 4496 44364 4548
rect 44416 4536 44422 4548
rect 45204 4536 45232 4567
rect 45554 4564 45560 4616
rect 45612 4604 45618 4616
rect 46569 4607 46627 4613
rect 46569 4604 46581 4607
rect 45612 4576 46581 4604
rect 45612 4564 45618 4576
rect 46216 4548 46244 4576
rect 46569 4573 46581 4576
rect 46615 4573 46627 4607
rect 46569 4567 46627 4573
rect 44416 4508 45232 4536
rect 44416 4496 44422 4508
rect 46198 4496 46204 4548
rect 46256 4496 46262 4548
rect 36924 4440 37688 4468
rect 40773 4471 40831 4477
rect 33229 4431 33287 4437
rect 40773 4437 40785 4471
rect 40819 4437 40831 4471
rect 40773 4431 40831 4437
rect 40862 4428 40868 4480
rect 40920 4468 40926 4480
rect 41233 4471 41291 4477
rect 41233 4468 41245 4471
rect 40920 4440 41245 4468
rect 40920 4428 40926 4440
rect 41233 4437 41245 4440
rect 41279 4437 41291 4471
rect 41233 4431 41291 4437
rect 1104 4378 58880 4400
rect 1104 4326 19574 4378
rect 19626 4326 19638 4378
rect 19690 4326 19702 4378
rect 19754 4326 19766 4378
rect 19818 4326 19830 4378
rect 19882 4326 50294 4378
rect 50346 4326 50358 4378
rect 50410 4326 50422 4378
rect 50474 4326 50486 4378
rect 50538 4326 50550 4378
rect 50602 4326 58880 4378
rect 1104 4304 58880 4326
rect 6454 4224 6460 4276
rect 6512 4264 6518 4276
rect 16022 4264 16028 4276
rect 6512 4236 16028 4264
rect 6512 4224 6518 4236
rect 6270 4156 6276 4208
rect 6328 4196 6334 4208
rect 6549 4199 6607 4205
rect 6549 4196 6561 4199
rect 6328 4168 6561 4196
rect 6328 4156 6334 4168
rect 6549 4165 6561 4168
rect 6595 4165 6607 4199
rect 6549 4159 6607 4165
rect 6365 4131 6423 4137
rect 6365 4097 6377 4131
rect 6411 4128 6423 4131
rect 6656 4128 6684 4236
rect 16022 4224 16028 4236
rect 16080 4224 16086 4276
rect 16206 4224 16212 4276
rect 16264 4264 16270 4276
rect 20530 4264 20536 4276
rect 16264 4236 20536 4264
rect 16264 4224 16270 4236
rect 20530 4224 20536 4236
rect 20588 4224 20594 4276
rect 45925 4267 45983 4273
rect 45925 4264 45937 4267
rect 45296 4236 45937 4264
rect 6730 4156 6736 4208
rect 6788 4196 6794 4208
rect 6788 4168 6833 4196
rect 6788 4156 6794 4168
rect 11146 4156 11152 4208
rect 11204 4196 11210 4208
rect 12710 4196 12716 4208
rect 11204 4168 12716 4196
rect 11204 4156 11210 4168
rect 12710 4156 12716 4168
rect 12768 4156 12774 4208
rect 12805 4199 12863 4205
rect 12805 4165 12817 4199
rect 12851 4196 12863 4199
rect 15746 4196 15752 4208
rect 12851 4168 15752 4196
rect 12851 4165 12863 4168
rect 12805 4159 12863 4165
rect 15746 4156 15752 4168
rect 15804 4156 15810 4208
rect 15838 4156 15844 4208
rect 15896 4156 15902 4208
rect 16040 4168 16896 4196
rect 9674 4128 9680 4140
rect 6411 4100 6684 4128
rect 9635 4100 9680 4128
rect 6411 4097 6423 4100
rect 6365 4091 6423 4097
rect 9674 4088 9680 4100
rect 9732 4088 9738 4140
rect 11790 4088 11796 4140
rect 11848 4128 11854 4140
rect 12529 4131 12587 4137
rect 12529 4128 12541 4131
rect 11848 4100 12541 4128
rect 11848 4088 11854 4100
rect 12529 4097 12541 4100
rect 12575 4097 12587 4131
rect 12529 4091 12587 4097
rect 12728 4100 15792 4128
rect 9766 4060 9772 4072
rect 9727 4032 9772 4060
rect 9766 4020 9772 4032
rect 9824 4020 9830 4072
rect 10318 4020 10324 4072
rect 10376 4060 10382 4072
rect 10413 4063 10471 4069
rect 10413 4060 10425 4063
rect 10376 4032 10425 4060
rect 10376 4020 10382 4032
rect 10413 4029 10425 4032
rect 10459 4060 10471 4063
rect 11330 4060 11336 4072
rect 10459 4032 11336 4060
rect 10459 4029 10471 4032
rect 10413 4023 10471 4029
rect 11330 4020 11336 4032
rect 11388 4060 11394 4072
rect 11882 4060 11888 4072
rect 11388 4032 11888 4060
rect 11388 4020 11394 4032
rect 11882 4020 11888 4032
rect 11940 4020 11946 4072
rect 11974 4020 11980 4072
rect 12032 4060 12038 4072
rect 12345 4063 12403 4069
rect 12345 4060 12357 4063
rect 12032 4032 12357 4060
rect 12032 4020 12038 4032
rect 12345 4029 12357 4032
rect 12391 4029 12403 4063
rect 12345 4023 12403 4029
rect 11054 3952 11060 4004
rect 11112 3992 11118 4004
rect 12728 3992 12756 4100
rect 12894 4060 12900 4072
rect 12855 4032 12900 4060
rect 12894 4020 12900 4032
rect 12952 4020 12958 4072
rect 15764 4060 15792 4100
rect 15856 4126 15884 4156
rect 15933 4131 15991 4137
rect 15933 4126 15945 4131
rect 15856 4098 15945 4126
rect 15933 4097 15945 4098
rect 15979 4128 15991 4131
rect 16040 4128 16068 4168
rect 15979 4100 16068 4128
rect 16117 4131 16175 4137
rect 15979 4097 15991 4100
rect 15933 4091 15991 4097
rect 16117 4097 16129 4131
rect 16163 4128 16175 4131
rect 16666 4128 16672 4140
rect 16163 4100 16672 4128
rect 16163 4097 16175 4100
rect 16117 4091 16175 4097
rect 16666 4088 16672 4100
rect 16724 4088 16730 4140
rect 16868 4137 16896 4168
rect 23750 4156 23756 4208
rect 23808 4196 23814 4208
rect 24029 4199 24087 4205
rect 24029 4196 24041 4199
rect 23808 4168 24041 4196
rect 23808 4156 23814 4168
rect 24029 4165 24041 4168
rect 24075 4165 24087 4199
rect 40862 4196 40868 4208
rect 24029 4159 24087 4165
rect 40420 4168 40868 4196
rect 16853 4131 16911 4137
rect 16853 4097 16865 4131
rect 16899 4128 16911 4131
rect 16899 4100 17954 4128
rect 16899 4097 16911 4100
rect 16853 4091 16911 4097
rect 17037 4063 17095 4069
rect 17037 4060 17049 4063
rect 15764 4032 17049 4060
rect 17037 4029 17049 4032
rect 17083 4060 17095 4063
rect 17678 4060 17684 4072
rect 17083 4032 17684 4060
rect 17083 4029 17095 4032
rect 17037 4023 17095 4029
rect 17678 4020 17684 4032
rect 17736 4020 17742 4072
rect 15933 3995 15991 4001
rect 15933 3992 15945 3995
rect 11112 3964 12756 3992
rect 13280 3964 15945 3992
rect 11112 3952 11118 3964
rect 11790 3924 11796 3936
rect 11751 3896 11796 3924
rect 11790 3884 11796 3896
rect 11848 3884 11854 3936
rect 12434 3884 12440 3936
rect 12492 3924 12498 3936
rect 13280 3924 13308 3964
rect 15933 3961 15945 3964
rect 15979 3992 15991 3995
rect 16666 3992 16672 4004
rect 15979 3964 16672 3992
rect 15979 3961 15991 3964
rect 15933 3955 15991 3961
rect 16666 3952 16672 3964
rect 16724 3952 16730 4004
rect 17926 3992 17954 4100
rect 20254 4088 20260 4140
rect 20312 4128 20318 4140
rect 20533 4131 20591 4137
rect 20533 4128 20545 4131
rect 20312 4100 20545 4128
rect 20312 4088 20318 4100
rect 20533 4097 20545 4100
rect 20579 4097 20591 4131
rect 20533 4091 20591 4097
rect 20622 4088 20628 4140
rect 20680 4128 20686 4140
rect 20717 4131 20775 4137
rect 20717 4128 20729 4131
rect 20680 4100 20729 4128
rect 20680 4088 20686 4100
rect 20717 4097 20729 4100
rect 20763 4097 20775 4131
rect 20717 4091 20775 4097
rect 23845 4131 23903 4137
rect 23845 4097 23857 4131
rect 23891 4128 23903 4131
rect 24762 4128 24768 4140
rect 23891 4100 24768 4128
rect 23891 4097 23903 4100
rect 23845 4091 23903 4097
rect 24762 4088 24768 4100
rect 24820 4088 24826 4140
rect 33134 4088 33140 4140
rect 33192 4128 33198 4140
rect 33505 4131 33563 4137
rect 33505 4128 33517 4131
rect 33192 4100 33517 4128
rect 33192 4088 33198 4100
rect 33505 4097 33517 4100
rect 33551 4128 33563 4131
rect 33594 4128 33600 4140
rect 33551 4100 33600 4128
rect 33551 4097 33563 4100
rect 33505 4091 33563 4097
rect 33594 4088 33600 4100
rect 33652 4088 33658 4140
rect 33686 4088 33692 4140
rect 33744 4128 33750 4140
rect 33744 4100 33789 4128
rect 33744 4088 33750 4100
rect 35802 4088 35808 4140
rect 35860 4128 35866 4140
rect 36265 4131 36323 4137
rect 36265 4128 36277 4131
rect 35860 4100 36277 4128
rect 35860 4088 35866 4100
rect 36265 4097 36277 4100
rect 36311 4097 36323 4131
rect 36446 4128 36452 4140
rect 36407 4100 36452 4128
rect 36265 4091 36323 4097
rect 36446 4088 36452 4100
rect 36504 4088 36510 4140
rect 40420 4137 40448 4168
rect 40862 4156 40868 4168
rect 40920 4156 40926 4208
rect 42242 4156 42248 4208
rect 42300 4196 42306 4208
rect 45296 4205 45324 4236
rect 45925 4233 45937 4236
rect 45971 4233 45983 4267
rect 45925 4227 45983 4233
rect 45097 4199 45155 4205
rect 45097 4196 45109 4199
rect 42300 4168 45109 4196
rect 42300 4156 42306 4168
rect 45097 4165 45109 4168
rect 45143 4165 45155 4199
rect 45097 4159 45155 4165
rect 45281 4199 45339 4205
rect 45281 4165 45293 4199
rect 45327 4165 45339 4199
rect 46290 4196 46296 4208
rect 46251 4168 46296 4196
rect 45281 4159 45339 4165
rect 46290 4156 46296 4168
rect 46348 4156 46354 4208
rect 37645 4131 37703 4137
rect 37645 4097 37657 4131
rect 37691 4097 37703 4131
rect 37645 4091 37703 4097
rect 40404 4131 40462 4137
rect 40404 4097 40416 4131
rect 40450 4097 40462 4131
rect 40404 4091 40462 4097
rect 20901 4063 20959 4069
rect 20901 4029 20913 4063
rect 20947 4060 20959 4063
rect 21634 4060 21640 4072
rect 20947 4032 21640 4060
rect 20947 4029 20959 4032
rect 20901 4023 20959 4029
rect 21634 4020 21640 4032
rect 21692 4020 21698 4072
rect 22186 4020 22192 4072
rect 22244 4060 22250 4072
rect 22244 4032 26004 4060
rect 22244 4020 22250 4032
rect 23382 3992 23388 4004
rect 17926 3964 23388 3992
rect 23382 3952 23388 3964
rect 23440 3952 23446 4004
rect 25866 3992 25872 4004
rect 23492 3964 25872 3992
rect 12492 3896 13308 3924
rect 12492 3884 12498 3896
rect 13446 3884 13452 3936
rect 13504 3924 13510 3936
rect 14645 3927 14703 3933
rect 14645 3924 14657 3927
rect 13504 3896 14657 3924
rect 13504 3884 13510 3896
rect 14645 3893 14657 3896
rect 14691 3924 14703 3927
rect 14918 3924 14924 3936
rect 14691 3896 14924 3924
rect 14691 3893 14703 3896
rect 14645 3887 14703 3893
rect 14918 3884 14924 3896
rect 14976 3884 14982 3936
rect 16942 3884 16948 3936
rect 17000 3924 17006 3936
rect 23492 3924 23520 3964
rect 25866 3952 25872 3964
rect 25924 3952 25930 4004
rect 25976 3992 26004 4032
rect 26418 4020 26424 4072
rect 26476 4060 26482 4072
rect 36633 4063 36691 4069
rect 26476 4032 36584 4060
rect 26476 4020 26482 4032
rect 27522 3992 27528 4004
rect 25976 3964 27528 3992
rect 27522 3952 27528 3964
rect 27580 3952 27586 4004
rect 29270 3952 29276 4004
rect 29328 3992 29334 4004
rect 36556 3992 36584 4032
rect 36633 4029 36645 4063
rect 36679 4060 36691 4063
rect 37366 4060 37372 4072
rect 36679 4032 37372 4060
rect 36679 4029 36691 4032
rect 36633 4023 36691 4029
rect 37366 4020 37372 4032
rect 37424 4020 37430 4072
rect 37550 4060 37556 4072
rect 37511 4032 37556 4060
rect 37550 4020 37556 4032
rect 37608 4020 37614 4072
rect 37660 4060 37688 4091
rect 40494 4088 40500 4140
rect 40552 4128 40558 4140
rect 41322 4128 41328 4140
rect 40552 4100 40597 4128
rect 41283 4100 41328 4128
rect 40552 4088 40558 4100
rect 41322 4088 41328 4100
rect 41380 4088 41386 4140
rect 41506 4128 41512 4140
rect 41467 4100 41512 4128
rect 41506 4088 41512 4100
rect 41564 4088 41570 4140
rect 46109 4131 46167 4137
rect 46109 4097 46121 4131
rect 46155 4097 46167 4131
rect 46109 4091 46167 4097
rect 37826 4060 37832 4072
rect 37660 4032 37832 4060
rect 37826 4020 37832 4032
rect 37884 4060 37890 4072
rect 40589 4063 40647 4069
rect 40589 4060 40601 4063
rect 37884 4032 40601 4060
rect 37884 4020 37890 4032
rect 40589 4029 40601 4032
rect 40635 4029 40647 4063
rect 40589 4023 40647 4029
rect 40678 4020 40684 4072
rect 40736 4060 40742 4072
rect 40865 4063 40923 4069
rect 40736 4032 40781 4060
rect 40736 4020 40742 4032
rect 40865 4029 40877 4063
rect 40911 4060 40923 4063
rect 46124 4060 46152 4091
rect 46198 4088 46204 4140
rect 46256 4128 46262 4140
rect 46477 4131 46535 4137
rect 46256 4100 46301 4128
rect 46256 4088 46262 4100
rect 46477 4097 46489 4131
rect 46523 4097 46535 4131
rect 46477 4091 46535 4097
rect 46382 4060 46388 4072
rect 40911 4032 46388 4060
rect 40911 4029 40923 4032
rect 40865 4023 40923 4029
rect 46382 4020 46388 4032
rect 46440 4020 46446 4072
rect 42058 3992 42064 4004
rect 29328 3964 36124 3992
rect 36556 3964 42064 3992
rect 29328 3952 29334 3964
rect 17000 3896 23520 3924
rect 17000 3884 17006 3896
rect 23566 3884 23572 3936
rect 23624 3924 23630 3936
rect 23661 3927 23719 3933
rect 23661 3924 23673 3927
rect 23624 3896 23673 3924
rect 23624 3884 23630 3896
rect 23661 3893 23673 3896
rect 23707 3893 23719 3927
rect 23661 3887 23719 3893
rect 33226 3884 33232 3936
rect 33284 3924 33290 3936
rect 33505 3927 33563 3933
rect 33505 3924 33517 3927
rect 33284 3896 33517 3924
rect 33284 3884 33290 3896
rect 33505 3893 33517 3896
rect 33551 3893 33563 3927
rect 36096 3924 36124 3964
rect 42058 3952 42064 3964
rect 42116 3952 42122 4004
rect 46106 3992 46112 4004
rect 44652 3964 46112 3992
rect 36538 3924 36544 3936
rect 36096 3896 36544 3924
rect 33505 3887 33563 3893
rect 36538 3884 36544 3896
rect 36596 3884 36602 3936
rect 37369 3927 37427 3933
rect 37369 3893 37381 3927
rect 37415 3924 37427 3927
rect 37458 3924 37464 3936
rect 37415 3896 37464 3924
rect 37415 3893 37427 3896
rect 37369 3887 37427 3893
rect 37458 3884 37464 3896
rect 37516 3884 37522 3936
rect 41046 3884 41052 3936
rect 41104 3924 41110 3936
rect 41325 3927 41383 3933
rect 41325 3924 41337 3927
rect 41104 3896 41337 3924
rect 41104 3884 41110 3896
rect 41325 3893 41337 3896
rect 41371 3893 41383 3927
rect 41325 3887 41383 3893
rect 41414 3884 41420 3936
rect 41472 3924 41478 3936
rect 44652 3924 44680 3964
rect 46106 3952 46112 3964
rect 46164 3992 46170 4004
rect 46492 3992 46520 4091
rect 46164 3964 46520 3992
rect 46164 3952 46170 3964
rect 41472 3896 44680 3924
rect 44913 3927 44971 3933
rect 41472 3884 41478 3896
rect 44913 3893 44925 3927
rect 44959 3924 44971 3927
rect 45186 3924 45192 3936
rect 44959 3896 45192 3924
rect 44959 3893 44971 3896
rect 44913 3887 44971 3893
rect 45186 3884 45192 3896
rect 45244 3884 45250 3936
rect 58066 3924 58072 3936
rect 58027 3896 58072 3924
rect 58066 3884 58072 3896
rect 58124 3884 58130 3936
rect 1104 3834 58880 3856
rect 1104 3782 4214 3834
rect 4266 3782 4278 3834
rect 4330 3782 4342 3834
rect 4394 3782 4406 3834
rect 4458 3782 4470 3834
rect 4522 3782 34934 3834
rect 34986 3782 34998 3834
rect 35050 3782 35062 3834
rect 35114 3782 35126 3834
rect 35178 3782 35190 3834
rect 35242 3782 58880 3834
rect 1104 3760 58880 3782
rect 9677 3723 9735 3729
rect 9677 3689 9689 3723
rect 9723 3720 9735 3723
rect 9766 3720 9772 3732
rect 9723 3692 9772 3720
rect 9723 3689 9735 3692
rect 9677 3683 9735 3689
rect 9766 3680 9772 3692
rect 9824 3680 9830 3732
rect 10042 3680 10048 3732
rect 10100 3720 10106 3732
rect 12434 3720 12440 3732
rect 10100 3692 12440 3720
rect 10100 3680 10106 3692
rect 12434 3680 12440 3692
rect 12492 3680 12498 3732
rect 12621 3723 12679 3729
rect 12621 3689 12633 3723
rect 12667 3720 12679 3723
rect 12894 3720 12900 3732
rect 12667 3692 12900 3720
rect 12667 3689 12679 3692
rect 12621 3683 12679 3689
rect 12894 3680 12900 3692
rect 12952 3680 12958 3732
rect 14918 3680 14924 3732
rect 14976 3720 14982 3732
rect 15657 3723 15715 3729
rect 15657 3720 15669 3723
rect 14976 3692 15669 3720
rect 14976 3680 14982 3692
rect 15657 3689 15669 3692
rect 15703 3720 15715 3723
rect 26142 3720 26148 3732
rect 15703 3692 26148 3720
rect 15703 3689 15715 3692
rect 15657 3683 15715 3689
rect 26142 3680 26148 3692
rect 26200 3680 26206 3732
rect 30208 3692 36492 3720
rect 14274 3652 14280 3664
rect 2746 3624 14280 3652
rect 2038 3544 2044 3596
rect 2096 3584 2102 3596
rect 2746 3584 2774 3624
rect 14274 3612 14280 3624
rect 14332 3612 14338 3664
rect 15010 3612 15016 3664
rect 15068 3652 15074 3664
rect 15105 3655 15163 3661
rect 15105 3652 15117 3655
rect 15068 3624 15117 3652
rect 15068 3612 15074 3624
rect 15105 3621 15117 3624
rect 15151 3652 15163 3655
rect 20898 3652 20904 3664
rect 15151 3624 20904 3652
rect 15151 3621 15163 3624
rect 15105 3615 15163 3621
rect 20898 3612 20904 3624
rect 20956 3612 20962 3664
rect 2096 3556 2774 3584
rect 2096 3544 2102 3556
rect 11882 3544 11888 3596
rect 11940 3584 11946 3596
rect 14461 3587 14519 3593
rect 11940 3556 12388 3584
rect 11940 3544 11946 3556
rect 10594 3476 10600 3528
rect 10652 3516 10658 3528
rect 10652 3488 10697 3516
rect 11241 3509 11299 3515
rect 10652 3476 10658 3488
rect 11241 3475 11253 3509
rect 11287 3506 11299 3509
rect 11330 3506 11336 3528
rect 11287 3478 11336 3506
rect 11287 3475 11299 3478
rect 11330 3476 11336 3478
rect 11388 3476 11394 3528
rect 11422 3476 11428 3528
rect 11480 3516 11486 3528
rect 12360 3516 12388 3556
rect 14461 3553 14473 3587
rect 14507 3584 14519 3587
rect 18046 3584 18052 3596
rect 14507 3556 14872 3584
rect 14507 3553 14519 3556
rect 14461 3547 14519 3553
rect 12805 3519 12863 3525
rect 12805 3516 12817 3519
rect 11480 3510 11573 3516
rect 11624 3510 12112 3516
rect 11480 3488 12112 3510
rect 12360 3488 12817 3516
rect 11480 3482 11652 3488
rect 11480 3476 11486 3482
rect 11241 3469 11299 3475
rect 9861 3451 9919 3457
rect 9861 3417 9873 3451
rect 9907 3417 9919 3451
rect 10042 3448 10048 3460
rect 10003 3420 10048 3448
rect 9861 3411 9919 3417
rect 1394 3380 1400 3392
rect 1355 3352 1400 3380
rect 1394 3340 1400 3352
rect 1452 3340 1458 3392
rect 9876 3380 9904 3411
rect 10042 3408 10048 3420
rect 10100 3408 10106 3460
rect 10689 3451 10747 3457
rect 10689 3417 10701 3451
rect 10735 3448 10747 3451
rect 11974 3448 11980 3460
rect 10735 3420 11192 3448
rect 10735 3417 10747 3420
rect 10689 3411 10747 3417
rect 11054 3380 11060 3392
rect 9876 3352 11060 3380
rect 11054 3340 11060 3352
rect 11112 3340 11118 3392
rect 11164 3380 11192 3420
rect 11348 3420 11980 3448
rect 11348 3380 11376 3420
rect 11974 3408 11980 3420
rect 12032 3408 12038 3460
rect 12084 3448 12112 3488
rect 12805 3485 12817 3488
rect 12851 3485 12863 3519
rect 12805 3479 12863 3485
rect 13173 3519 13231 3525
rect 13173 3485 13185 3519
rect 13219 3516 13231 3519
rect 13446 3516 13452 3528
rect 13219 3488 13452 3516
rect 13219 3485 13231 3488
rect 13173 3479 13231 3485
rect 13446 3476 13452 3488
rect 13504 3476 13510 3528
rect 14277 3519 14335 3525
rect 14277 3516 14289 3519
rect 14108 3488 14289 3516
rect 12897 3451 12955 3457
rect 12897 3448 12909 3451
rect 12084 3420 12909 3448
rect 12897 3417 12909 3420
rect 12943 3417 12955 3451
rect 12897 3411 12955 3417
rect 12989 3451 13047 3457
rect 12989 3417 13001 3451
rect 13035 3448 13047 3451
rect 14108 3448 14136 3488
rect 14277 3485 14289 3488
rect 14323 3516 14335 3519
rect 14844 3516 14872 3556
rect 16868 3556 18052 3584
rect 14918 3516 14924 3528
rect 14323 3488 14504 3516
rect 14844 3488 14924 3516
rect 14323 3485 14335 3488
rect 14277 3479 14335 3485
rect 13035 3420 14136 3448
rect 14476 3448 14504 3488
rect 14918 3476 14924 3488
rect 14976 3476 14982 3528
rect 15102 3516 15108 3528
rect 15063 3488 15108 3516
rect 15102 3476 15108 3488
rect 15160 3476 15166 3528
rect 16666 3516 16672 3528
rect 16627 3488 16672 3516
rect 16666 3476 16672 3488
rect 16724 3476 16730 3528
rect 16868 3525 16896 3556
rect 18046 3544 18052 3556
rect 18104 3544 18110 3596
rect 19168 3556 21036 3584
rect 16853 3519 16911 3525
rect 16853 3485 16865 3519
rect 16899 3485 16911 3519
rect 17310 3516 17316 3528
rect 17271 3488 17316 3516
rect 16853 3479 16911 3485
rect 17310 3476 17316 3488
rect 17368 3476 17374 3528
rect 17402 3476 17408 3528
rect 17460 3516 17466 3528
rect 17678 3516 17684 3528
rect 17460 3488 17505 3516
rect 17639 3488 17684 3516
rect 17460 3476 17466 3488
rect 17678 3476 17684 3488
rect 17736 3476 17742 3528
rect 17819 3519 17877 3525
rect 17819 3485 17831 3519
rect 17865 3516 17877 3519
rect 19168 3516 19196 3556
rect 17865 3488 19196 3516
rect 17865 3485 17877 3488
rect 17819 3479 17877 3485
rect 19242 3476 19248 3528
rect 19300 3516 19306 3528
rect 19300 3488 19393 3516
rect 19300 3476 19306 3488
rect 15120 3448 15148 3476
rect 14476 3420 15148 3448
rect 16761 3451 16819 3457
rect 13035 3417 13047 3420
rect 12989 3411 13047 3417
rect 16761 3417 16773 3451
rect 16807 3448 16819 3451
rect 17589 3451 17647 3457
rect 17589 3448 17601 3451
rect 16807 3420 17601 3448
rect 16807 3417 16819 3420
rect 16761 3411 16819 3417
rect 17589 3417 17601 3420
rect 17635 3417 17647 3451
rect 18601 3451 18659 3457
rect 18601 3448 18613 3451
rect 17589 3411 17647 3417
rect 17696 3420 18613 3448
rect 11164 3352 11376 3380
rect 11425 3383 11483 3389
rect 11425 3349 11437 3383
rect 11471 3380 11483 3383
rect 11514 3380 11520 3392
rect 11471 3352 11520 3380
rect 11471 3349 11483 3352
rect 11425 3343 11483 3349
rect 11514 3340 11520 3352
rect 11572 3340 11578 3392
rect 14090 3380 14096 3392
rect 14051 3352 14096 3380
rect 14090 3340 14096 3352
rect 14148 3340 14154 3392
rect 14274 3340 14280 3392
rect 14332 3380 14338 3392
rect 17696 3380 17724 3420
rect 18601 3417 18613 3420
rect 18647 3417 18659 3451
rect 19352 3448 19380 3488
rect 19426 3476 19432 3528
rect 19484 3516 19490 3528
rect 20073 3519 20131 3525
rect 20073 3516 20085 3519
rect 19484 3488 20085 3516
rect 19484 3476 19490 3488
rect 20073 3485 20085 3488
rect 20119 3485 20131 3519
rect 20254 3516 20260 3528
rect 20215 3488 20260 3516
rect 20073 3479 20131 3485
rect 20254 3476 20260 3488
rect 20312 3476 20318 3528
rect 19889 3451 19947 3457
rect 19889 3448 19901 3451
rect 19352 3420 19901 3448
rect 18601 3411 18659 3417
rect 19889 3417 19901 3420
rect 19935 3417 19947 3451
rect 19889 3411 19947 3417
rect 17954 3380 17960 3392
rect 14332 3352 17724 3380
rect 17915 3352 17960 3380
rect 14332 3340 14338 3352
rect 17954 3340 17960 3352
rect 18012 3340 18018 3392
rect 18616 3380 18644 3411
rect 19334 3380 19340 3392
rect 18616 3352 19340 3380
rect 19334 3340 19340 3352
rect 19392 3340 19398 3392
rect 19429 3383 19487 3389
rect 19429 3349 19441 3383
rect 19475 3380 19487 3383
rect 20622 3380 20628 3392
rect 19475 3352 20628 3380
rect 19475 3349 19487 3352
rect 19429 3343 19487 3349
rect 20622 3340 20628 3352
rect 20680 3340 20686 3392
rect 21008 3380 21036 3556
rect 23934 3544 23940 3596
rect 23992 3584 23998 3596
rect 23992 3556 24716 3584
rect 23992 3544 23998 3556
rect 21082 3476 21088 3528
rect 21140 3516 21146 3528
rect 21269 3519 21327 3525
rect 21269 3516 21281 3519
rect 21140 3488 21281 3516
rect 21140 3476 21146 3488
rect 21269 3485 21281 3488
rect 21315 3485 21327 3519
rect 21634 3516 21640 3528
rect 21595 3488 21640 3516
rect 21269 3479 21327 3485
rect 21634 3476 21640 3488
rect 21692 3476 21698 3528
rect 23750 3476 23756 3528
rect 23808 3516 23814 3528
rect 24581 3519 24639 3525
rect 24581 3516 24593 3519
rect 23808 3488 24593 3516
rect 23808 3476 23814 3488
rect 24581 3485 24593 3488
rect 24627 3485 24639 3519
rect 24688 3516 24716 3556
rect 24762 3544 24768 3596
rect 24820 3584 24826 3596
rect 28534 3584 28540 3596
rect 24820 3556 28540 3584
rect 24820 3544 24826 3556
rect 28534 3544 28540 3556
rect 28592 3544 28598 3596
rect 28902 3584 28908 3596
rect 28863 3556 28908 3584
rect 28902 3544 28908 3556
rect 28960 3544 28966 3596
rect 26145 3519 26203 3525
rect 26145 3516 26157 3519
rect 24688 3488 26157 3516
rect 24581 3479 24639 3485
rect 26145 3485 26157 3488
rect 26191 3485 26203 3519
rect 26418 3516 26424 3528
rect 26379 3488 26424 3516
rect 26145 3479 26203 3485
rect 26418 3476 26424 3488
rect 26476 3476 26482 3528
rect 28813 3519 28871 3525
rect 28813 3485 28825 3519
rect 28859 3516 28871 3519
rect 30208 3516 30236 3692
rect 33686 3612 33692 3664
rect 33744 3612 33750 3664
rect 36464 3652 36492 3692
rect 36538 3680 36544 3732
rect 36596 3720 36602 3732
rect 57793 3723 57851 3729
rect 57793 3720 57805 3723
rect 36596 3692 57805 3720
rect 36596 3680 36602 3692
rect 57793 3689 57805 3692
rect 57839 3689 57851 3723
rect 57793 3683 57851 3689
rect 37645 3655 37703 3661
rect 36464 3624 37596 3652
rect 31941 3587 31999 3593
rect 31941 3584 31953 3587
rect 31312 3556 31953 3584
rect 31312 3525 31340 3556
rect 31941 3553 31953 3556
rect 31987 3553 31999 3587
rect 32861 3587 32919 3593
rect 32861 3584 32873 3587
rect 31941 3547 31999 3553
rect 32048 3556 32873 3584
rect 28859 3488 30236 3516
rect 31297 3519 31355 3525
rect 28859 3485 28871 3488
rect 28813 3479 28871 3485
rect 31297 3485 31309 3519
rect 31343 3485 31355 3519
rect 31297 3479 31355 3485
rect 31481 3519 31539 3525
rect 31481 3485 31493 3519
rect 31527 3516 31539 3519
rect 32048 3516 32076 3556
rect 32861 3553 32873 3556
rect 32907 3584 32919 3587
rect 33042 3584 33048 3596
rect 32907 3556 33048 3584
rect 32907 3553 32919 3556
rect 32861 3547 32919 3553
rect 33042 3544 33048 3556
rect 33100 3544 33106 3596
rect 33505 3587 33563 3593
rect 33505 3553 33517 3587
rect 33551 3584 33563 3587
rect 33704 3584 33732 3612
rect 36354 3584 36360 3596
rect 33551 3556 36360 3584
rect 33551 3553 33563 3556
rect 33505 3547 33563 3553
rect 36354 3544 36360 3556
rect 36412 3544 36418 3596
rect 31527 3488 32076 3516
rect 32125 3519 32183 3525
rect 31527 3485 31539 3488
rect 31481 3479 31539 3485
rect 32125 3485 32137 3519
rect 32171 3485 32183 3519
rect 32125 3479 32183 3485
rect 23109 3451 23167 3457
rect 23109 3417 23121 3451
rect 23155 3448 23167 3451
rect 32140 3448 32168 3479
rect 32214 3476 32220 3528
rect 32272 3516 32278 3528
rect 32769 3519 32827 3525
rect 32769 3516 32781 3519
rect 32272 3488 32781 3516
rect 32272 3476 32278 3488
rect 32769 3485 32781 3488
rect 32815 3485 32827 3519
rect 32769 3479 32827 3485
rect 32953 3519 33011 3525
rect 32953 3485 32965 3519
rect 32999 3485 33011 3519
rect 32953 3479 33011 3485
rect 32968 3448 32996 3479
rect 33594 3476 33600 3528
rect 33652 3516 33658 3528
rect 33689 3519 33747 3525
rect 33689 3516 33701 3519
rect 33652 3488 33701 3516
rect 33652 3476 33658 3488
rect 33689 3485 33701 3488
rect 33735 3485 33747 3519
rect 33870 3516 33876 3528
rect 33831 3488 33876 3516
rect 33689 3479 33747 3485
rect 33870 3476 33876 3488
rect 33928 3476 33934 3528
rect 37090 3516 37096 3528
rect 37051 3488 37096 3516
rect 37090 3476 37096 3488
rect 37148 3476 37154 3528
rect 37274 3516 37280 3528
rect 37235 3488 37280 3516
rect 37274 3476 37280 3488
rect 37332 3476 37338 3528
rect 37458 3516 37464 3528
rect 37419 3488 37464 3516
rect 37458 3476 37464 3488
rect 37516 3476 37522 3528
rect 34238 3448 34244 3460
rect 23155 3420 31754 3448
rect 32140 3420 34244 3448
rect 23155 3417 23167 3420
rect 23109 3411 23167 3417
rect 23750 3380 23756 3392
rect 21008 3352 23756 3380
rect 23750 3340 23756 3352
rect 23808 3380 23814 3392
rect 24210 3380 24216 3392
rect 23808 3352 24216 3380
rect 23808 3340 23814 3352
rect 24210 3340 24216 3352
rect 24268 3340 24274 3392
rect 24394 3380 24400 3392
rect 24355 3352 24400 3380
rect 24394 3340 24400 3352
rect 24452 3340 24458 3392
rect 25958 3380 25964 3392
rect 25919 3352 25964 3380
rect 25958 3340 25964 3352
rect 26016 3340 26022 3392
rect 26326 3380 26332 3392
rect 26287 3352 26332 3380
rect 26326 3340 26332 3352
rect 26384 3340 26390 3392
rect 26970 3380 26976 3392
rect 26931 3352 26976 3380
rect 26970 3340 26976 3352
rect 27028 3340 27034 3392
rect 27706 3380 27712 3392
rect 27667 3352 27712 3380
rect 27706 3340 27712 3352
rect 27764 3340 27770 3392
rect 28350 3340 28356 3392
rect 28408 3380 28414 3392
rect 28445 3383 28503 3389
rect 28445 3380 28457 3383
rect 28408 3352 28457 3380
rect 28408 3340 28414 3352
rect 28445 3349 28457 3352
rect 28491 3349 28503 3383
rect 28445 3343 28503 3349
rect 28534 3340 28540 3392
rect 28592 3380 28598 3392
rect 31389 3383 31447 3389
rect 31389 3380 31401 3383
rect 28592 3352 31401 3380
rect 28592 3340 28598 3352
rect 31389 3349 31401 3352
rect 31435 3349 31447 3383
rect 31726 3380 31754 3420
rect 34238 3408 34244 3420
rect 34296 3408 34302 3460
rect 37366 3408 37372 3460
rect 37424 3448 37430 3460
rect 37568 3448 37596 3624
rect 37645 3621 37657 3655
rect 37691 3621 37703 3655
rect 37645 3615 37703 3621
rect 37660 3516 37688 3615
rect 37734 3612 37740 3664
rect 37792 3652 37798 3664
rect 41598 3652 41604 3664
rect 37792 3624 41414 3652
rect 41559 3624 41604 3652
rect 37792 3612 37798 3624
rect 41386 3584 41414 3624
rect 41598 3612 41604 3624
rect 41656 3612 41662 3664
rect 42058 3652 42064 3664
rect 42019 3624 42064 3652
rect 42058 3612 42064 3624
rect 42116 3612 42122 3664
rect 46201 3587 46259 3593
rect 40144 3556 41184 3584
rect 41386 3556 45968 3584
rect 40034 3516 40040 3528
rect 37660 3488 40040 3516
rect 40034 3476 40040 3488
rect 40092 3476 40098 3528
rect 40144 3448 40172 3556
rect 40221 3519 40279 3525
rect 40221 3485 40233 3519
rect 40267 3485 40279 3519
rect 40862 3516 40868 3528
rect 40823 3488 40868 3516
rect 40221 3479 40279 3485
rect 37424 3420 37469 3448
rect 37568 3420 40172 3448
rect 40236 3448 40264 3479
rect 40862 3476 40868 3488
rect 40920 3476 40926 3528
rect 41046 3516 41052 3528
rect 41007 3488 41052 3516
rect 41046 3476 41052 3488
rect 41104 3476 41110 3528
rect 41156 3516 41184 3556
rect 43070 3516 43076 3528
rect 41156 3488 43076 3516
rect 43070 3476 43076 3488
rect 43128 3476 43134 3528
rect 43165 3519 43223 3525
rect 43165 3485 43177 3519
rect 43211 3516 43223 3519
rect 43254 3516 43260 3528
rect 43211 3488 43260 3516
rect 43211 3485 43223 3488
rect 43165 3479 43223 3485
rect 43254 3476 43260 3488
rect 43312 3516 43318 3528
rect 43809 3519 43867 3525
rect 43809 3516 43821 3519
rect 43312 3488 43821 3516
rect 43312 3476 43318 3488
rect 43809 3485 43821 3488
rect 43855 3485 43867 3519
rect 43809 3479 43867 3485
rect 40957 3451 41015 3457
rect 40957 3448 40969 3451
rect 40236 3420 40969 3448
rect 37424 3408 37430 3420
rect 40880 3392 40908 3420
rect 40957 3417 40969 3420
rect 41003 3417 41015 3451
rect 42242 3448 42248 3460
rect 42203 3420 42248 3448
rect 40957 3411 41015 3417
rect 42242 3408 42248 3420
rect 42300 3408 42306 3460
rect 42426 3448 42432 3460
rect 42387 3420 42432 3448
rect 42426 3408 42432 3420
rect 42484 3408 42490 3460
rect 42610 3408 42616 3460
rect 42668 3448 42674 3460
rect 45940 3448 45968 3556
rect 46201 3553 46213 3587
rect 46247 3584 46259 3587
rect 46290 3584 46296 3596
rect 46247 3556 46296 3584
rect 46247 3553 46259 3556
rect 46201 3547 46259 3553
rect 46290 3544 46296 3556
rect 46348 3544 46354 3596
rect 46106 3516 46112 3528
rect 46067 3488 46112 3516
rect 46106 3476 46112 3488
rect 46164 3476 46170 3528
rect 58066 3516 58072 3528
rect 58027 3488 58072 3516
rect 58066 3476 58072 3488
rect 58124 3476 58130 3528
rect 57606 3448 57612 3460
rect 42668 3420 45784 3448
rect 45940 3420 57612 3448
rect 42668 3408 42674 3420
rect 37734 3380 37740 3392
rect 31726 3352 37740 3380
rect 31389 3343 31447 3349
rect 37734 3340 37740 3352
rect 37792 3340 37798 3392
rect 40218 3380 40224 3392
rect 40179 3352 40224 3380
rect 40218 3340 40224 3352
rect 40276 3340 40282 3392
rect 40862 3340 40868 3392
rect 40920 3340 40926 3392
rect 41322 3340 41328 3392
rect 41380 3380 41386 3392
rect 43162 3380 43168 3392
rect 41380 3352 43168 3380
rect 41380 3340 41386 3352
rect 43162 3340 43168 3352
rect 43220 3340 43226 3392
rect 43346 3380 43352 3392
rect 43307 3352 43352 3380
rect 43346 3340 43352 3352
rect 43404 3340 43410 3392
rect 45756 3389 45784 3420
rect 57606 3408 57612 3420
rect 57664 3408 57670 3460
rect 45741 3383 45799 3389
rect 45741 3349 45753 3383
rect 45787 3349 45799 3383
rect 57146 3380 57152 3392
rect 57107 3352 57152 3380
rect 45741 3343 45799 3349
rect 57146 3340 57152 3352
rect 57204 3340 57210 3392
rect 1104 3290 58880 3312
rect 1104 3238 19574 3290
rect 19626 3238 19638 3290
rect 19690 3238 19702 3290
rect 19754 3238 19766 3290
rect 19818 3238 19830 3290
rect 19882 3238 50294 3290
rect 50346 3238 50358 3290
rect 50410 3238 50422 3290
rect 50474 3238 50486 3290
rect 50538 3238 50550 3290
rect 50602 3238 58880 3290
rect 1104 3216 58880 3238
rect 4617 3179 4675 3185
rect 4617 3145 4629 3179
rect 4663 3176 4675 3179
rect 4982 3176 4988 3188
rect 4663 3148 4988 3176
rect 4663 3145 4675 3148
rect 4617 3139 4675 3145
rect 4982 3136 4988 3148
rect 5040 3136 5046 3188
rect 10134 3136 10140 3188
rect 10192 3176 10198 3188
rect 11330 3176 11336 3188
rect 10192 3148 11336 3176
rect 10192 3136 10198 3148
rect 11330 3136 11336 3148
rect 11388 3136 11394 3188
rect 11514 3176 11520 3188
rect 11475 3148 11520 3176
rect 11514 3136 11520 3148
rect 11572 3136 11578 3188
rect 15102 3136 15108 3188
rect 15160 3176 15166 3188
rect 16669 3179 16727 3185
rect 16669 3176 16681 3179
rect 15160 3148 16681 3176
rect 15160 3136 15166 3148
rect 16669 3145 16681 3148
rect 16715 3145 16727 3179
rect 19242 3176 19248 3188
rect 19203 3148 19248 3176
rect 16669 3139 16727 3145
rect 19242 3136 19248 3148
rect 19300 3136 19306 3188
rect 19334 3136 19340 3188
rect 19392 3176 19398 3188
rect 19705 3179 19763 3185
rect 19705 3176 19717 3179
rect 19392 3148 19717 3176
rect 19392 3136 19398 3148
rect 19705 3145 19717 3148
rect 19751 3145 19763 3179
rect 23382 3176 23388 3188
rect 19705 3139 19763 3145
rect 20456 3148 22094 3176
rect 23343 3148 23388 3176
rect 1394 3040 1400 3052
rect 1355 3012 1400 3040
rect 1394 3000 1400 3012
rect 1452 3000 1458 3052
rect 5000 3040 5028 3136
rect 10873 3111 10931 3117
rect 10873 3108 10885 3111
rect 5460 3080 10885 3108
rect 5460 3049 5488 3080
rect 10873 3077 10885 3080
rect 10919 3077 10931 3111
rect 14090 3108 14096 3120
rect 14051 3080 14096 3108
rect 10873 3071 10931 3077
rect 5445 3043 5503 3049
rect 5445 3040 5457 3043
rect 5000 3012 5457 3040
rect 5445 3009 5457 3012
rect 5491 3009 5503 3043
rect 10134 3040 10140 3052
rect 10095 3012 10140 3040
rect 5445 3003 5503 3009
rect 10134 3000 10140 3012
rect 10192 3000 10198 3052
rect 10318 3040 10324 3052
rect 10279 3012 10324 3040
rect 10318 3000 10324 3012
rect 10376 3000 10382 3052
rect 1673 2975 1731 2981
rect 1673 2941 1685 2975
rect 1719 2972 1731 2975
rect 5537 2975 5595 2981
rect 1719 2944 5488 2972
rect 1719 2941 1731 2944
rect 1673 2935 1731 2941
rect 5074 2904 5080 2916
rect 5035 2876 5080 2904
rect 5074 2864 5080 2876
rect 5132 2864 5138 2916
rect 5460 2904 5488 2944
rect 5537 2941 5549 2975
rect 5583 2972 5595 2975
rect 9309 2975 9367 2981
rect 9309 2972 9321 2975
rect 5583 2944 9321 2972
rect 5583 2941 5595 2944
rect 5537 2935 5595 2941
rect 9309 2941 9321 2944
rect 9355 2972 9367 2975
rect 10594 2972 10600 2984
rect 9355 2944 10600 2972
rect 9355 2941 9367 2944
rect 9309 2935 9367 2941
rect 10594 2932 10600 2944
rect 10652 2932 10658 2984
rect 10888 2972 10916 3071
rect 14090 3068 14096 3080
rect 14148 3068 14154 3120
rect 14277 3111 14335 3117
rect 14277 3077 14289 3111
rect 14323 3108 14335 3111
rect 15010 3108 15016 3120
rect 14323 3080 15016 3108
rect 14323 3077 14335 3080
rect 14277 3071 14335 3077
rect 15010 3068 15016 3080
rect 15068 3068 15074 3120
rect 17773 3111 17831 3117
rect 17773 3108 17785 3111
rect 17052 3080 17785 3108
rect 11974 3040 11980 3052
rect 11935 3012 11980 3040
rect 11974 3000 11980 3012
rect 12032 3000 12038 3052
rect 17052 3049 17080 3080
rect 17773 3077 17785 3080
rect 17819 3077 17831 3111
rect 20456 3108 20484 3148
rect 21634 3108 21640 3120
rect 17773 3071 17831 3077
rect 18892 3080 20484 3108
rect 20732 3080 21640 3108
rect 13081 3043 13139 3049
rect 13081 3009 13093 3043
rect 13127 3040 13139 3043
rect 13909 3043 13967 3049
rect 13909 3040 13921 3043
rect 13127 3012 13921 3040
rect 13127 3009 13139 3012
rect 13081 3003 13139 3009
rect 13909 3009 13921 3012
rect 13955 3009 13967 3043
rect 13909 3003 13967 3009
rect 17037 3043 17095 3049
rect 17037 3009 17049 3043
rect 17083 3009 17095 3043
rect 17037 3003 17095 3009
rect 17310 3000 17316 3052
rect 17368 3040 17374 3052
rect 17681 3043 17739 3049
rect 17681 3040 17693 3043
rect 17368 3012 17693 3040
rect 17368 3000 17374 3012
rect 17681 3009 17693 3012
rect 17727 3009 17739 3043
rect 17681 3003 17739 3009
rect 17865 3043 17923 3049
rect 17865 3009 17877 3043
rect 17911 3040 17923 3043
rect 18046 3040 18052 3052
rect 17911 3012 18052 3040
rect 17911 3009 17923 3012
rect 17865 3003 17923 3009
rect 11790 2972 11796 2984
rect 10888 2944 11796 2972
rect 11790 2932 11796 2944
rect 11848 2972 11854 2984
rect 11885 2975 11943 2981
rect 11885 2972 11897 2975
rect 11848 2944 11897 2972
rect 11848 2932 11854 2944
rect 11885 2941 11897 2944
rect 11931 2941 11943 2975
rect 11885 2935 11943 2941
rect 12161 2975 12219 2981
rect 12161 2941 12173 2975
rect 12207 2972 12219 2975
rect 12989 2975 13047 2981
rect 12989 2972 13001 2975
rect 12207 2944 13001 2972
rect 12207 2941 12219 2944
rect 12161 2935 12219 2941
rect 12989 2941 13001 2944
rect 13035 2941 13047 2975
rect 16942 2972 16948 2984
rect 16903 2944 16948 2972
rect 12989 2935 13047 2941
rect 16942 2932 16948 2944
rect 17000 2932 17006 2984
rect 7374 2904 7380 2916
rect 5460 2876 7380 2904
rect 7374 2864 7380 2876
rect 7432 2864 7438 2916
rect 9674 2864 9680 2916
rect 9732 2904 9738 2916
rect 13446 2904 13452 2916
rect 9732 2876 12434 2904
rect 13407 2876 13452 2904
rect 9732 2864 9738 2876
rect 14 2796 20 2848
rect 72 2836 78 2848
rect 1486 2836 1492 2848
rect 72 2808 1492 2836
rect 72 2796 78 2808
rect 1486 2796 1492 2808
rect 1544 2836 1550 2848
rect 2317 2839 2375 2845
rect 2317 2836 2329 2839
rect 1544 2808 2329 2836
rect 1544 2796 1550 2808
rect 2317 2805 2329 2808
rect 2363 2805 2375 2839
rect 2317 2799 2375 2805
rect 2590 2796 2596 2848
rect 2648 2836 2654 2848
rect 2869 2839 2927 2845
rect 2869 2836 2881 2839
rect 2648 2808 2881 2836
rect 2648 2796 2654 2808
rect 2869 2805 2881 2808
rect 2915 2805 2927 2839
rect 8478 2836 8484 2848
rect 8439 2808 8484 2836
rect 2869 2799 2927 2805
rect 8478 2796 8484 2808
rect 8536 2796 8542 2848
rect 12406 2836 12434 2876
rect 13446 2864 13452 2876
rect 13504 2864 13510 2916
rect 17402 2836 17408 2848
rect 12406 2808 17408 2836
rect 17402 2796 17408 2808
rect 17460 2796 17466 2848
rect 17696 2836 17724 3003
rect 18046 3000 18052 3012
rect 18104 3000 18110 3052
rect 18892 3049 18920 3080
rect 18877 3043 18935 3049
rect 18877 3009 18889 3043
rect 18923 3009 18935 3043
rect 18877 3003 18935 3009
rect 20533 3043 20591 3049
rect 20533 3009 20545 3043
rect 20579 3040 20591 3043
rect 20622 3040 20628 3052
rect 20579 3012 20628 3040
rect 20579 3009 20591 3012
rect 20533 3003 20591 3009
rect 20622 3000 20628 3012
rect 20680 3000 20686 3052
rect 20732 3049 20760 3080
rect 21634 3068 21640 3080
rect 21692 3068 21698 3120
rect 22066 3108 22094 3148
rect 23382 3136 23388 3148
rect 23440 3136 23446 3188
rect 25869 3179 25927 3185
rect 25869 3176 25881 3179
rect 24044 3148 25881 3176
rect 24044 3108 24072 3148
rect 25869 3145 25881 3148
rect 25915 3145 25927 3179
rect 25869 3139 25927 3145
rect 26804 3148 27200 3176
rect 22066 3080 24072 3108
rect 24210 3068 24216 3120
rect 24268 3108 24274 3120
rect 25317 3111 25375 3117
rect 24268 3080 24440 3108
rect 24268 3068 24274 3080
rect 20717 3043 20775 3049
rect 20717 3009 20729 3043
rect 20763 3009 20775 3043
rect 20717 3003 20775 3009
rect 20809 3043 20867 3049
rect 20809 3009 20821 3043
rect 20855 3040 20867 3043
rect 20855 3012 20944 3040
rect 20855 3009 20867 3012
rect 20809 3003 20867 3009
rect 20916 2984 20944 3012
rect 21726 3000 21732 3052
rect 21784 3040 21790 3052
rect 24302 3040 24308 3052
rect 21784 3012 24308 3040
rect 21784 3000 21790 3012
rect 24302 3000 24308 3012
rect 24360 3000 24366 3052
rect 24412 3040 24440 3080
rect 25317 3077 25329 3111
rect 25363 3108 25375 3111
rect 26804 3108 26832 3148
rect 25363 3080 26832 3108
rect 25363 3077 25375 3080
rect 25317 3071 25375 3077
rect 26878 3068 26884 3120
rect 26936 3108 26942 3120
rect 26936 3080 27016 3108
rect 26936 3068 26942 3080
rect 26988 3049 27016 3080
rect 27172 3049 27200 3148
rect 31726 3148 36308 3176
rect 27338 3068 27344 3120
rect 27396 3108 27402 3120
rect 31113 3111 31171 3117
rect 27396 3080 29684 3108
rect 27396 3068 27402 3080
rect 24486 3043 24544 3049
rect 24486 3040 24498 3043
rect 24412 3012 24498 3040
rect 24486 3009 24498 3012
rect 24532 3009 24544 3043
rect 24486 3003 24544 3009
rect 25409 3043 25467 3049
rect 25409 3009 25421 3043
rect 25455 3040 25467 3043
rect 26237 3043 26295 3049
rect 26237 3040 26249 3043
rect 25455 3012 26249 3040
rect 25455 3009 25467 3012
rect 25409 3003 25467 3009
rect 26237 3009 26249 3012
rect 26283 3009 26295 3043
rect 26237 3003 26295 3009
rect 26973 3043 27031 3049
rect 26973 3009 26985 3043
rect 27019 3009 27031 3043
rect 26973 3003 27031 3009
rect 27157 3043 27215 3049
rect 27157 3009 27169 3043
rect 27203 3009 27215 3043
rect 27157 3003 27215 3009
rect 17954 2932 17960 2984
rect 18012 2972 18018 2984
rect 18785 2975 18843 2981
rect 18785 2972 18797 2975
rect 18012 2944 18797 2972
rect 18012 2932 18018 2944
rect 18785 2941 18797 2944
rect 18831 2941 18843 2975
rect 18785 2935 18843 2941
rect 20898 2932 20904 2984
rect 20956 2932 20962 2984
rect 23658 2932 23664 2984
rect 23716 2972 23722 2984
rect 23845 2975 23903 2981
rect 23845 2972 23857 2975
rect 23716 2944 23857 2972
rect 23716 2932 23722 2944
rect 23845 2941 23857 2944
rect 23891 2972 23903 2975
rect 24394 2972 24400 2984
rect 23891 2944 24400 2972
rect 23891 2941 23903 2944
rect 23845 2935 23903 2941
rect 24394 2932 24400 2944
rect 24452 2972 24458 2984
rect 24673 2975 24731 2981
rect 24673 2972 24685 2975
rect 24452 2944 24685 2972
rect 24452 2932 24458 2944
rect 24673 2941 24685 2944
rect 24719 2941 24731 2975
rect 26142 2972 26148 2984
rect 26103 2944 26148 2972
rect 24673 2935 24731 2941
rect 26142 2932 26148 2944
rect 26200 2932 26206 2984
rect 26252 2972 26280 3003
rect 27246 3000 27252 3052
rect 27304 3040 27310 3052
rect 27893 3043 27951 3049
rect 27893 3040 27905 3043
rect 27304 3012 27905 3040
rect 27304 3000 27310 3012
rect 27893 3009 27905 3012
rect 27939 3009 27951 3043
rect 28350 3040 28356 3052
rect 28311 3012 28356 3040
rect 27893 3003 27951 3009
rect 28350 3000 28356 3012
rect 28408 3000 28414 3052
rect 29656 3049 29684 3080
rect 31113 3077 31125 3111
rect 31159 3108 31171 3111
rect 31726 3108 31754 3148
rect 33870 3108 33876 3120
rect 31159 3080 31754 3108
rect 33244 3080 33548 3108
rect 33831 3080 33876 3108
rect 31159 3077 31171 3080
rect 31113 3071 31171 3077
rect 33244 3052 33272 3080
rect 28721 3043 28779 3049
rect 28721 3009 28733 3043
rect 28767 3040 28779 3043
rect 29273 3043 29331 3049
rect 29273 3040 29285 3043
rect 28767 3012 29285 3040
rect 28767 3009 28779 3012
rect 28721 3003 28779 3009
rect 29273 3009 29285 3012
rect 29319 3009 29331 3043
rect 29273 3003 29331 3009
rect 29641 3043 29699 3049
rect 29641 3009 29653 3043
rect 29687 3009 29699 3043
rect 33042 3040 33048 3052
rect 33003 3012 33048 3040
rect 29641 3003 29699 3009
rect 33042 3000 33048 3012
rect 33100 3000 33106 3052
rect 33226 3040 33232 3052
rect 33187 3012 33232 3040
rect 33226 3000 33232 3012
rect 33284 3000 33290 3052
rect 33410 3040 33416 3052
rect 33371 3012 33416 3040
rect 33410 3000 33416 3012
rect 33468 3000 33474 3052
rect 33520 3040 33548 3080
rect 33870 3068 33876 3080
rect 33928 3068 33934 3120
rect 34238 3108 34244 3120
rect 34199 3080 34244 3108
rect 34238 3068 34244 3080
rect 34296 3068 34302 3120
rect 36280 3108 36308 3148
rect 36354 3136 36360 3188
rect 36412 3176 36418 3188
rect 37277 3179 37335 3185
rect 37277 3176 37289 3179
rect 36412 3148 37289 3176
rect 36412 3136 36418 3148
rect 37277 3145 37289 3148
rect 37323 3145 37335 3179
rect 37277 3139 37335 3145
rect 40218 3136 40224 3188
rect 40276 3176 40282 3188
rect 41690 3176 41696 3188
rect 40276 3148 41696 3176
rect 40276 3136 40282 3148
rect 41690 3136 41696 3148
rect 41748 3136 41754 3188
rect 42426 3176 42432 3188
rect 42387 3148 42432 3176
rect 42426 3136 42432 3148
rect 42484 3136 42490 3188
rect 43162 3136 43168 3188
rect 43220 3176 43226 3188
rect 57146 3176 57152 3188
rect 43220 3148 57152 3176
rect 43220 3136 43226 3148
rect 57146 3136 57152 3148
rect 57204 3136 57210 3188
rect 41322 3108 41328 3120
rect 36280 3080 41328 3108
rect 41322 3068 41328 3080
rect 41380 3068 41386 3120
rect 42610 3117 42616 3120
rect 42597 3111 42616 3117
rect 42597 3077 42609 3111
rect 42597 3071 42616 3077
rect 41592 3065 41650 3071
rect 42610 3068 42616 3071
rect 42668 3068 42674 3120
rect 42797 3111 42855 3117
rect 42797 3077 42809 3111
rect 42843 3077 42855 3111
rect 42797 3071 42855 3077
rect 41592 3062 41604 3065
rect 34057 3043 34115 3049
rect 34057 3040 34069 3043
rect 33520 3012 34069 3040
rect 34057 3009 34069 3012
rect 34103 3009 34115 3043
rect 34057 3003 34115 3009
rect 35802 3000 35808 3052
rect 35860 3040 35866 3052
rect 36541 3043 36599 3049
rect 36541 3040 36553 3043
rect 35860 3012 36553 3040
rect 35860 3000 35866 3012
rect 36541 3009 36553 3012
rect 36587 3009 36599 3043
rect 36541 3003 36599 3009
rect 26326 2972 26332 2984
rect 26252 2944 26332 2972
rect 26326 2932 26332 2944
rect 26384 2972 26390 2984
rect 26384 2944 27476 2972
rect 26384 2932 26390 2944
rect 20530 2864 20536 2916
rect 20588 2904 20594 2916
rect 20625 2907 20683 2913
rect 20625 2904 20637 2907
rect 20588 2876 20637 2904
rect 20588 2864 20594 2876
rect 20625 2873 20637 2876
rect 20671 2873 20683 2907
rect 20625 2867 20683 2873
rect 20993 2907 21051 2913
rect 20993 2873 21005 2907
rect 21039 2904 21051 2907
rect 23566 2904 23572 2916
rect 21039 2876 23428 2904
rect 23527 2876 23572 2904
rect 21039 2873 21051 2876
rect 20993 2867 21051 2873
rect 21726 2836 21732 2848
rect 17696 2808 21732 2836
rect 21726 2796 21732 2808
rect 21784 2796 21790 2848
rect 21910 2836 21916 2848
rect 21871 2808 21916 2836
rect 21910 2796 21916 2808
rect 21968 2796 21974 2848
rect 23400 2836 23428 2876
rect 23566 2864 23572 2876
rect 23624 2864 23630 2916
rect 27338 2904 27344 2916
rect 26436 2876 27344 2904
rect 26436 2836 26464 2876
rect 27338 2864 27344 2876
rect 27396 2864 27402 2916
rect 27448 2904 27476 2944
rect 32582 2904 32588 2916
rect 27448 2876 32588 2904
rect 32582 2864 32588 2876
rect 32640 2904 32646 2916
rect 33045 2907 33103 2913
rect 33045 2904 33057 2907
rect 32640 2876 33057 2904
rect 32640 2864 32646 2876
rect 33045 2873 33057 2876
rect 33091 2873 33103 2907
rect 33045 2867 33103 2873
rect 23400 2808 26464 2836
rect 26510 2796 26516 2848
rect 26568 2836 26574 2848
rect 26973 2839 27031 2845
rect 26973 2836 26985 2839
rect 26568 2808 26985 2836
rect 26568 2796 26574 2808
rect 26973 2805 26985 2808
rect 27019 2805 27031 2839
rect 26973 2799 27031 2805
rect 31570 2796 31576 2848
rect 31628 2836 31634 2848
rect 32125 2839 32183 2845
rect 32125 2836 32137 2839
rect 31628 2808 32137 2836
rect 31628 2796 31634 2808
rect 32125 2805 32137 2808
rect 32171 2805 32183 2839
rect 32125 2799 32183 2805
rect 33410 2796 33416 2848
rect 33468 2836 33474 2848
rect 36265 2839 36323 2845
rect 36265 2836 36277 2839
rect 33468 2808 36277 2836
rect 33468 2796 33474 2808
rect 36265 2805 36277 2808
rect 36311 2805 36323 2839
rect 36556 2836 36584 3003
rect 37366 3000 37372 3052
rect 37424 3040 37430 3052
rect 37645 3043 37703 3049
rect 37645 3040 37657 3043
rect 37424 3012 37657 3040
rect 37424 3000 37430 3012
rect 37645 3009 37657 3012
rect 37691 3009 37703 3043
rect 37645 3003 37703 3009
rect 39761 3043 39819 3049
rect 39761 3009 39773 3043
rect 39807 3009 39819 3043
rect 39761 3003 39819 3009
rect 36633 2975 36691 2981
rect 36633 2941 36645 2975
rect 36679 2941 36691 2975
rect 36633 2935 36691 2941
rect 36648 2904 36676 2935
rect 37458 2932 37464 2984
rect 37516 2972 37522 2984
rect 37553 2975 37611 2981
rect 37553 2972 37565 2975
rect 37516 2944 37565 2972
rect 37516 2932 37522 2944
rect 37553 2941 37565 2944
rect 37599 2941 37611 2975
rect 37553 2935 37611 2941
rect 39776 2904 39804 3003
rect 40034 3000 40040 3052
rect 40092 3040 40098 3052
rect 40681 3043 40739 3049
rect 40681 3040 40693 3043
rect 40092 3012 40693 3040
rect 40092 3000 40098 3012
rect 40681 3009 40693 3012
rect 40727 3009 40739 3043
rect 40862 3040 40868 3052
rect 40823 3012 40868 3040
rect 40681 3003 40739 3009
rect 40862 3000 40868 3012
rect 40920 3000 40926 3052
rect 41432 3034 41604 3062
rect 39942 2904 39948 2916
rect 36648 2876 39948 2904
rect 39942 2864 39948 2876
rect 40000 2864 40006 2916
rect 40221 2907 40279 2913
rect 40221 2873 40233 2907
rect 40267 2904 40279 2907
rect 41432 2904 41460 3034
rect 41592 3031 41604 3034
rect 41638 3031 41650 3065
rect 41592 3025 41650 3031
rect 41877 3043 41935 3049
rect 41877 3009 41889 3043
rect 41923 3040 41935 3043
rect 42628 3040 42656 3068
rect 41923 3012 42656 3040
rect 41923 3009 41935 3012
rect 41877 3003 41935 3009
rect 41690 2932 41696 2984
rect 41748 2972 41754 2984
rect 42812 2972 42840 3071
rect 43070 3068 43076 3120
rect 43128 3108 43134 3120
rect 44545 3111 44603 3117
rect 44545 3108 44557 3111
rect 43128 3080 44557 3108
rect 43128 3068 43134 3080
rect 44545 3077 44557 3080
rect 44591 3077 44603 3111
rect 44545 3071 44603 3077
rect 45094 3068 45100 3120
rect 45152 3108 45158 3120
rect 45152 3080 51074 3108
rect 45152 3068 45158 3080
rect 43438 3000 43444 3052
rect 43496 3040 43502 3052
rect 43717 3043 43775 3049
rect 43717 3040 43729 3043
rect 43496 3012 43729 3040
rect 43496 3000 43502 3012
rect 43717 3009 43729 3012
rect 43763 3009 43775 3043
rect 44913 3043 44971 3049
rect 44913 3040 44925 3043
rect 43717 3003 43775 3009
rect 44100 3012 44925 3040
rect 43806 2972 43812 2984
rect 41748 2944 42840 2972
rect 43767 2944 43812 2972
rect 41748 2932 41754 2944
rect 43806 2932 43812 2944
rect 43864 2932 43870 2984
rect 44100 2981 44128 3012
rect 44913 3009 44925 3012
rect 44959 3009 44971 3043
rect 45186 3040 45192 3052
rect 45147 3012 45192 3040
rect 44913 3003 44971 3009
rect 45186 3000 45192 3012
rect 45244 3000 45250 3052
rect 51046 3040 51074 3080
rect 51353 3043 51411 3049
rect 51353 3040 51365 3043
rect 51046 3012 51365 3040
rect 51353 3009 51365 3012
rect 51399 3040 51411 3043
rect 51997 3043 52055 3049
rect 51997 3040 52009 3043
rect 51399 3012 52009 3040
rect 51399 3009 51411 3012
rect 51353 3003 51411 3009
rect 51997 3009 52009 3012
rect 52043 3009 52055 3043
rect 57164 3040 57192 3136
rect 57885 3043 57943 3049
rect 57885 3040 57897 3043
rect 57164 3012 57897 3040
rect 51997 3003 52055 3009
rect 57885 3009 57897 3012
rect 57931 3009 57943 3043
rect 57885 3003 57943 3009
rect 44085 2975 44143 2981
rect 44085 2941 44097 2975
rect 44131 2941 44143 2975
rect 44085 2935 44143 2941
rect 51537 2907 51595 2913
rect 40267 2876 42656 2904
rect 40267 2873 40279 2876
rect 40221 2867 40279 2873
rect 39853 2839 39911 2845
rect 39853 2836 39865 2839
rect 36556 2808 39865 2836
rect 36265 2799 36323 2805
rect 39853 2805 39865 2808
rect 39899 2805 39911 2839
rect 39853 2799 39911 2805
rect 40126 2796 40132 2848
rect 40184 2836 40190 2848
rect 41049 2839 41107 2845
rect 41049 2836 41061 2839
rect 40184 2808 41061 2836
rect 40184 2796 40190 2808
rect 41049 2805 41061 2808
rect 41095 2805 41107 2839
rect 41049 2799 41107 2805
rect 41877 2839 41935 2845
rect 41877 2805 41889 2839
rect 41923 2836 41935 2839
rect 42242 2836 42248 2848
rect 41923 2808 42248 2836
rect 41923 2805 41935 2808
rect 41877 2799 41935 2805
rect 42242 2796 42248 2808
rect 42300 2796 42306 2848
rect 42628 2845 42656 2876
rect 51537 2873 51549 2907
rect 51583 2904 51595 2907
rect 52730 2904 52736 2916
rect 51583 2876 52736 2904
rect 51583 2873 51595 2876
rect 51537 2867 51595 2873
rect 52730 2864 52736 2876
rect 52788 2864 52794 2916
rect 42613 2839 42671 2845
rect 42613 2805 42625 2839
rect 42659 2805 42671 2839
rect 42613 2799 42671 2805
rect 56042 2796 56048 2848
rect 56100 2836 56106 2848
rect 56597 2839 56655 2845
rect 56597 2836 56609 2839
rect 56100 2808 56609 2836
rect 56100 2796 56106 2808
rect 56597 2805 56609 2808
rect 56643 2805 56655 2839
rect 57238 2836 57244 2848
rect 57199 2808 57244 2836
rect 56597 2799 56655 2805
rect 57238 2796 57244 2808
rect 57296 2796 57302 2848
rect 58069 2839 58127 2845
rect 58069 2805 58081 2839
rect 58115 2836 58127 2839
rect 59906 2836 59912 2848
rect 58115 2808 59912 2836
rect 58115 2805 58127 2808
rect 58069 2799 58127 2805
rect 59906 2796 59912 2808
rect 59964 2796 59970 2848
rect 1104 2746 58880 2768
rect 1104 2694 4214 2746
rect 4266 2694 4278 2746
rect 4330 2694 4342 2746
rect 4394 2694 4406 2746
rect 4458 2694 4470 2746
rect 4522 2694 34934 2746
rect 34986 2694 34998 2746
rect 35050 2694 35062 2746
rect 35114 2694 35126 2746
rect 35178 2694 35190 2746
rect 35242 2694 58880 2746
rect 1104 2672 58880 2694
rect 2777 2635 2835 2641
rect 2777 2601 2789 2635
rect 2823 2632 2835 2635
rect 4890 2632 4896 2644
rect 2823 2604 4896 2632
rect 2823 2601 2835 2604
rect 2777 2595 2835 2601
rect 4890 2592 4896 2604
rect 4948 2592 4954 2644
rect 21266 2632 21272 2644
rect 6886 2604 21272 2632
rect 2041 2499 2099 2505
rect 2041 2465 2053 2499
rect 2087 2496 2099 2499
rect 5718 2496 5724 2508
rect 2087 2468 5724 2496
rect 2087 2465 2099 2468
rect 2041 2459 2099 2465
rect 5718 2456 5724 2468
rect 5776 2496 5782 2508
rect 6886 2496 6914 2604
rect 21266 2592 21272 2604
rect 21324 2592 21330 2644
rect 22189 2635 22247 2641
rect 22189 2601 22201 2635
rect 22235 2632 22247 2635
rect 22554 2632 22560 2644
rect 22235 2604 22560 2632
rect 22235 2601 22247 2604
rect 22189 2595 22247 2601
rect 22554 2592 22560 2604
rect 22612 2592 22618 2644
rect 23753 2635 23811 2641
rect 23753 2601 23765 2635
rect 23799 2632 23811 2635
rect 23842 2632 23848 2644
rect 23799 2604 23848 2632
rect 23799 2601 23811 2604
rect 23753 2595 23811 2601
rect 23842 2592 23848 2604
rect 23900 2592 23906 2644
rect 24210 2592 24216 2644
rect 24268 2632 24274 2644
rect 26878 2632 26884 2644
rect 24268 2604 26884 2632
rect 24268 2592 24274 2604
rect 26878 2592 26884 2604
rect 26936 2592 26942 2644
rect 27062 2592 27068 2644
rect 27120 2632 27126 2644
rect 27157 2635 27215 2641
rect 27157 2632 27169 2635
rect 27120 2604 27169 2632
rect 27120 2592 27126 2604
rect 27157 2601 27169 2604
rect 27203 2601 27215 2635
rect 27157 2595 27215 2601
rect 28074 2592 28080 2644
rect 28132 2632 28138 2644
rect 31389 2635 31447 2641
rect 31389 2632 31401 2635
rect 28132 2604 31401 2632
rect 28132 2592 28138 2604
rect 31389 2601 31401 2604
rect 31435 2601 31447 2635
rect 31389 2595 31447 2601
rect 31726 2604 32628 2632
rect 8754 2524 8760 2576
rect 8812 2564 8818 2576
rect 31726 2564 31754 2604
rect 8812 2536 31754 2564
rect 8812 2524 8818 2536
rect 8110 2496 8116 2508
rect 5776 2468 6914 2496
rect 8071 2468 8116 2496
rect 5776 2456 5782 2468
rect 8110 2456 8116 2468
rect 8168 2456 8174 2508
rect 10045 2499 10103 2505
rect 10045 2465 10057 2499
rect 10091 2496 10103 2499
rect 10134 2496 10140 2508
rect 10091 2468 10140 2496
rect 10091 2465 10103 2468
rect 10045 2459 10103 2465
rect 10134 2456 10140 2468
rect 10192 2456 10198 2508
rect 10502 2456 10508 2508
rect 10560 2496 10566 2508
rect 15565 2499 15623 2505
rect 15565 2496 15577 2499
rect 10560 2468 15577 2496
rect 10560 2456 10566 2468
rect 15565 2465 15577 2468
rect 15611 2465 15623 2499
rect 15565 2459 15623 2465
rect 20622 2456 20628 2508
rect 20680 2496 20686 2508
rect 21082 2496 21088 2508
rect 20680 2468 20944 2496
rect 21043 2468 21088 2496
rect 20680 2456 20686 2468
rect 1486 2428 1492 2440
rect 1447 2400 1492 2428
rect 1486 2388 1492 2400
rect 1544 2388 1550 2440
rect 1946 2388 1952 2440
rect 2004 2428 2010 2440
rect 2590 2428 2596 2440
rect 2004 2400 2596 2428
rect 2004 2388 2010 2400
rect 2590 2388 2596 2400
rect 2648 2388 2654 2440
rect 4249 2431 4307 2437
rect 4249 2397 4261 2431
rect 4295 2428 4307 2431
rect 5074 2428 5080 2440
rect 4295 2400 5080 2428
rect 4295 2397 4307 2400
rect 4249 2391 4307 2397
rect 5074 2388 5080 2400
rect 5132 2388 5138 2440
rect 7742 2388 7748 2440
rect 7800 2428 7806 2440
rect 8389 2431 8447 2437
rect 8389 2428 8401 2431
rect 7800 2400 8401 2428
rect 7800 2388 7806 2400
rect 8389 2397 8401 2400
rect 8435 2428 8447 2431
rect 8478 2428 8484 2440
rect 8435 2400 8484 2428
rect 8435 2397 8447 2400
rect 8389 2391 8447 2397
rect 8478 2388 8484 2400
rect 8536 2388 8542 2440
rect 9309 2431 9367 2437
rect 9309 2397 9321 2431
rect 9355 2428 9367 2431
rect 9674 2428 9680 2440
rect 9355 2400 9680 2428
rect 9355 2397 9367 2400
rect 9309 2391 9367 2397
rect 9674 2388 9680 2400
rect 9732 2428 9738 2440
rect 9769 2431 9827 2437
rect 9769 2428 9781 2431
rect 9732 2400 9781 2428
rect 9732 2388 9738 2400
rect 9769 2397 9781 2400
rect 9815 2397 9827 2431
rect 9769 2391 9827 2397
rect 11977 2431 12035 2437
rect 11977 2397 11989 2431
rect 12023 2428 12035 2431
rect 12023 2400 12572 2428
rect 12023 2397 12035 2400
rect 11977 2391 12035 2397
rect 12544 2304 12572 2400
rect 13446 2388 13452 2440
rect 13504 2428 13510 2440
rect 14093 2431 14151 2437
rect 14093 2428 14105 2431
rect 13504 2400 14105 2428
rect 13504 2388 13510 2400
rect 14093 2397 14105 2400
rect 14139 2397 14151 2431
rect 14093 2391 14151 2397
rect 15289 2431 15347 2437
rect 15289 2397 15301 2431
rect 15335 2428 15347 2431
rect 15470 2428 15476 2440
rect 15335 2400 15476 2428
rect 15335 2397 15347 2400
rect 15289 2391 15347 2397
rect 15470 2388 15476 2400
rect 15528 2388 15534 2440
rect 17681 2431 17739 2437
rect 17681 2397 17693 2431
rect 17727 2428 17739 2431
rect 18414 2428 18420 2440
rect 17727 2400 18420 2428
rect 17727 2397 17739 2400
rect 17681 2391 17739 2397
rect 18414 2388 18420 2400
rect 18472 2388 18478 2440
rect 19150 2388 19156 2440
rect 19208 2428 19214 2440
rect 20806 2428 20812 2440
rect 19208 2400 20208 2428
rect 20767 2400 20812 2428
rect 19208 2388 19214 2400
rect 15488 2360 15516 2388
rect 16669 2363 16727 2369
rect 16669 2360 16681 2363
rect 15488 2332 16681 2360
rect 16669 2329 16681 2332
rect 16715 2329 16727 2363
rect 16669 2323 16727 2329
rect 19521 2363 19579 2369
rect 19521 2329 19533 2363
rect 19567 2360 19579 2363
rect 19978 2360 19984 2372
rect 19567 2332 19984 2360
rect 19567 2329 19579 2332
rect 19521 2323 19579 2329
rect 19978 2320 19984 2332
rect 20036 2360 20042 2372
rect 20073 2363 20131 2369
rect 20073 2360 20085 2363
rect 20036 2332 20085 2360
rect 20036 2320 20042 2332
rect 20073 2329 20085 2332
rect 20119 2329 20131 2363
rect 20180 2360 20208 2400
rect 20806 2388 20812 2400
rect 20864 2388 20870 2440
rect 20916 2437 20944 2468
rect 21082 2456 21088 2468
rect 21140 2456 21146 2508
rect 23658 2496 23664 2508
rect 21192 2468 23060 2496
rect 20901 2431 20959 2437
rect 20901 2397 20913 2431
rect 20947 2397 20959 2431
rect 20901 2391 20959 2397
rect 21192 2360 21220 2468
rect 21910 2388 21916 2440
rect 21968 2428 21974 2440
rect 22005 2431 22063 2437
rect 22005 2428 22017 2431
rect 21968 2400 22017 2428
rect 21968 2388 21974 2400
rect 22005 2397 22017 2400
rect 22051 2397 22063 2431
rect 22005 2391 22063 2397
rect 20180 2332 21220 2360
rect 20073 2323 20131 2329
rect 3878 2252 3884 2304
rect 3936 2292 3942 2304
rect 4065 2295 4123 2301
rect 4065 2292 4077 2295
rect 3936 2264 4077 2292
rect 3936 2252 3942 2264
rect 4065 2261 4077 2264
rect 4111 2261 4123 2295
rect 4065 2255 4123 2261
rect 11606 2252 11612 2304
rect 11664 2292 11670 2304
rect 11793 2295 11851 2301
rect 11793 2292 11805 2295
rect 11664 2264 11805 2292
rect 11664 2252 11670 2264
rect 11793 2261 11805 2264
rect 11839 2261 11851 2295
rect 12526 2292 12532 2304
rect 12487 2264 12532 2292
rect 11793 2255 11851 2261
rect 12526 2252 12532 2264
rect 12584 2252 12590 2304
rect 13538 2252 13544 2304
rect 13596 2292 13602 2304
rect 14277 2295 14335 2301
rect 14277 2292 14289 2295
rect 13596 2264 14289 2292
rect 13596 2252 13602 2264
rect 14277 2261 14289 2264
rect 14323 2261 14335 2295
rect 14277 2255 14335 2261
rect 18046 2252 18052 2304
rect 18104 2292 18110 2304
rect 18233 2295 18291 2301
rect 18233 2292 18245 2295
rect 18104 2264 18245 2292
rect 18104 2252 18110 2264
rect 18233 2261 18245 2264
rect 18279 2261 18291 2295
rect 20162 2292 20168 2304
rect 20123 2264 20168 2292
rect 18233 2255 18291 2261
rect 20162 2252 20168 2264
rect 20220 2252 20226 2304
rect 23032 2292 23060 2468
rect 23584 2468 23664 2496
rect 23584 2437 23612 2468
rect 23658 2456 23664 2468
rect 23716 2456 23722 2508
rect 25133 2499 25191 2505
rect 25133 2465 25145 2499
rect 25179 2496 25191 2499
rect 25774 2496 25780 2508
rect 25179 2468 25780 2496
rect 25179 2465 25191 2468
rect 25133 2459 25191 2465
rect 25774 2456 25780 2468
rect 25832 2456 25838 2508
rect 25958 2496 25964 2508
rect 25919 2468 25964 2496
rect 25958 2456 25964 2468
rect 26016 2456 26022 2508
rect 26326 2496 26332 2508
rect 26160 2468 26332 2496
rect 23569 2431 23627 2437
rect 23569 2397 23581 2431
rect 23615 2397 23627 2431
rect 23750 2428 23756 2440
rect 23711 2400 23756 2428
rect 23569 2391 23627 2397
rect 23750 2388 23756 2400
rect 23808 2388 23814 2440
rect 25866 2428 25872 2440
rect 25827 2400 25872 2428
rect 25866 2388 25872 2400
rect 25924 2388 25930 2440
rect 26160 2437 26188 2468
rect 26326 2456 26332 2468
rect 26384 2456 26390 2508
rect 26421 2499 26479 2505
rect 26421 2465 26433 2499
rect 26467 2496 26479 2499
rect 26694 2496 26700 2508
rect 26467 2468 26700 2496
rect 26467 2465 26479 2468
rect 26421 2459 26479 2465
rect 26694 2456 26700 2468
rect 26752 2456 26758 2508
rect 26878 2456 26884 2508
rect 26936 2496 26942 2508
rect 32217 2499 32275 2505
rect 32217 2496 32229 2499
rect 26936 2468 32229 2496
rect 26936 2456 26942 2468
rect 32217 2465 32229 2468
rect 32263 2465 32275 2499
rect 32600 2496 32628 2604
rect 33042 2592 33048 2644
rect 33100 2632 33106 2644
rect 33229 2635 33287 2641
rect 33229 2632 33241 2635
rect 33100 2604 33241 2632
rect 33100 2592 33106 2604
rect 33229 2601 33241 2604
rect 33275 2601 33287 2635
rect 39942 2632 39948 2644
rect 39903 2604 39948 2632
rect 33229 2595 33287 2601
rect 39942 2592 39948 2604
rect 40000 2592 40006 2644
rect 46106 2592 46112 2644
rect 46164 2632 46170 2644
rect 46661 2635 46719 2641
rect 46661 2632 46673 2635
rect 46164 2604 46673 2632
rect 46164 2592 46170 2604
rect 46661 2601 46673 2604
rect 46707 2632 46719 2635
rect 50982 2632 50988 2644
rect 46707 2604 50988 2632
rect 46707 2601 46719 2604
rect 46661 2595 46719 2601
rect 50982 2592 50988 2604
rect 51040 2592 51046 2644
rect 51166 2632 51172 2644
rect 51079 2604 51172 2632
rect 51166 2592 51172 2604
rect 51224 2632 51230 2644
rect 52362 2632 52368 2644
rect 51224 2604 52368 2632
rect 51224 2592 51230 2604
rect 52362 2592 52368 2604
rect 52420 2592 52426 2644
rect 55858 2592 55864 2644
rect 55916 2632 55922 2644
rect 56965 2635 57023 2641
rect 56965 2632 56977 2635
rect 55916 2604 56977 2632
rect 55916 2592 55922 2604
rect 56965 2601 56977 2604
rect 57011 2601 57023 2635
rect 56965 2595 57023 2601
rect 32674 2524 32680 2576
rect 32732 2564 32738 2576
rect 36357 2567 36415 2573
rect 32732 2536 35894 2564
rect 32732 2524 32738 2536
rect 34885 2499 34943 2505
rect 34885 2496 34897 2499
rect 32600 2468 34897 2496
rect 32217 2459 32275 2465
rect 34885 2465 34897 2468
rect 34931 2465 34943 2499
rect 35866 2496 35894 2536
rect 36357 2533 36369 2567
rect 36403 2564 36415 2567
rect 48498 2564 48504 2576
rect 36403 2536 48504 2564
rect 36403 2533 36415 2536
rect 36357 2527 36415 2533
rect 48498 2524 48504 2536
rect 48556 2524 48562 2576
rect 48593 2567 48651 2573
rect 48593 2533 48605 2567
rect 48639 2564 48651 2567
rect 52546 2564 52552 2576
rect 48639 2536 52552 2564
rect 48639 2533 48651 2536
rect 48593 2527 48651 2533
rect 35866 2468 45554 2496
rect 34885 2459 34943 2465
rect 26145 2431 26203 2437
rect 26145 2397 26157 2431
rect 26191 2397 26203 2431
rect 26145 2391 26203 2397
rect 26237 2431 26295 2437
rect 26237 2397 26249 2431
rect 26283 2428 26295 2431
rect 26510 2428 26516 2440
rect 26283 2400 26516 2428
rect 26283 2397 26295 2400
rect 26237 2391 26295 2397
rect 26510 2388 26516 2400
rect 26568 2388 26574 2440
rect 26970 2428 26976 2440
rect 26931 2400 26976 2428
rect 26970 2388 26976 2400
rect 27028 2388 27034 2440
rect 27706 2388 27712 2440
rect 27764 2428 27770 2440
rect 27801 2431 27859 2437
rect 27801 2428 27813 2431
rect 27764 2400 27813 2428
rect 27764 2388 27770 2400
rect 27801 2397 27813 2400
rect 27847 2397 27859 2431
rect 27801 2391 27859 2397
rect 28442 2388 28448 2440
rect 28500 2428 28506 2440
rect 31570 2428 31576 2440
rect 28500 2400 30328 2428
rect 31531 2400 31576 2428
rect 28500 2388 28506 2400
rect 23109 2363 23167 2369
rect 23109 2329 23121 2363
rect 23155 2360 23167 2363
rect 23842 2360 23848 2372
rect 23155 2332 23848 2360
rect 23155 2329 23167 2332
rect 23109 2323 23167 2329
rect 23842 2320 23848 2332
rect 23900 2360 23906 2372
rect 24857 2363 24915 2369
rect 24857 2360 24869 2363
rect 23900 2332 24869 2360
rect 23900 2320 23906 2332
rect 24857 2329 24869 2332
rect 24903 2329 24915 2363
rect 24857 2323 24915 2329
rect 26694 2320 26700 2372
rect 26752 2360 26758 2372
rect 27246 2360 27252 2372
rect 26752 2332 27252 2360
rect 26752 2320 26758 2332
rect 27246 2320 27252 2332
rect 27304 2320 27310 2372
rect 28077 2363 28135 2369
rect 28077 2329 28089 2363
rect 28123 2329 28135 2363
rect 28077 2323 28135 2329
rect 28997 2363 29055 2369
rect 28997 2329 29009 2363
rect 29043 2360 29055 2363
rect 29638 2360 29644 2372
rect 29043 2332 29644 2360
rect 29043 2329 29055 2332
rect 28997 2323 29055 2329
rect 28092 2292 28120 2323
rect 29638 2320 29644 2332
rect 29696 2360 29702 2372
rect 30009 2363 30067 2369
rect 30009 2360 30021 2363
rect 29696 2332 30021 2360
rect 29696 2320 29702 2332
rect 30009 2329 30021 2332
rect 30055 2329 30067 2363
rect 30300 2360 30328 2400
rect 31570 2388 31576 2400
rect 31628 2388 31634 2440
rect 32401 2431 32459 2437
rect 32401 2397 32413 2431
rect 32447 2397 32459 2431
rect 32582 2428 32588 2440
rect 32543 2400 32588 2428
rect 32401 2391 32459 2397
rect 32416 2360 32444 2391
rect 32582 2388 32588 2400
rect 32640 2388 32646 2440
rect 33226 2428 33232 2440
rect 33187 2400 33232 2428
rect 33226 2388 33232 2400
rect 33284 2388 33290 2440
rect 33410 2388 33416 2440
rect 33468 2428 33474 2440
rect 34701 2431 34759 2437
rect 34701 2428 34713 2431
rect 33468 2400 33513 2428
rect 34164 2400 34713 2428
rect 33468 2388 33474 2400
rect 30300 2332 31754 2360
rect 32416 2332 33088 2360
rect 30009 2323 30067 2329
rect 30098 2292 30104 2304
rect 23032 2264 28120 2292
rect 30059 2264 30104 2292
rect 30098 2252 30104 2264
rect 30156 2252 30162 2304
rect 31726 2292 31754 2332
rect 32674 2292 32680 2304
rect 31726 2264 32680 2292
rect 32674 2252 32680 2264
rect 32732 2252 32738 2304
rect 33060 2301 33088 2332
rect 34164 2304 34192 2400
rect 34701 2397 34713 2400
rect 34747 2397 34759 2431
rect 34701 2391 34759 2397
rect 35713 2431 35771 2437
rect 35713 2397 35725 2431
rect 35759 2428 35771 2431
rect 36078 2428 36084 2440
rect 35759 2400 36084 2428
rect 35759 2397 35771 2400
rect 35713 2391 35771 2397
rect 36078 2388 36084 2400
rect 36136 2428 36142 2440
rect 36173 2431 36231 2437
rect 36173 2428 36185 2431
rect 36136 2400 36185 2428
rect 36136 2388 36142 2400
rect 36173 2397 36185 2400
rect 36219 2397 36231 2431
rect 38105 2431 38163 2437
rect 38105 2428 38117 2431
rect 36173 2391 36231 2397
rect 37568 2400 38117 2428
rect 37568 2304 37596 2400
rect 38105 2397 38117 2400
rect 38151 2397 38163 2431
rect 40126 2428 40132 2440
rect 40087 2400 40132 2428
rect 38105 2391 38163 2397
rect 40126 2388 40132 2400
rect 40184 2388 40190 2440
rect 40218 2388 40224 2440
rect 40276 2428 40282 2440
rect 41049 2431 41107 2437
rect 40276 2400 40321 2428
rect 40276 2388 40282 2400
rect 41049 2397 41061 2431
rect 41095 2428 41107 2431
rect 41598 2428 41604 2440
rect 41095 2400 41604 2428
rect 41095 2397 41107 2400
rect 41049 2391 41107 2397
rect 41598 2388 41604 2400
rect 41656 2388 41662 2440
rect 42429 2431 42487 2437
rect 42429 2428 42441 2431
rect 41892 2400 42441 2428
rect 41892 2304 41920 2400
rect 42429 2397 42441 2400
rect 42475 2397 42487 2431
rect 42429 2391 42487 2397
rect 43346 2388 43352 2440
rect 43404 2428 43410 2440
rect 43901 2431 43959 2437
rect 43901 2428 43913 2431
rect 43404 2400 43913 2428
rect 43404 2388 43410 2400
rect 43901 2397 43913 2400
rect 43947 2397 43959 2431
rect 43901 2391 43959 2397
rect 42702 2360 42708 2372
rect 42663 2332 42708 2360
rect 42702 2320 42708 2332
rect 42760 2320 42766 2372
rect 45526 2360 45554 2468
rect 46106 2428 46112 2440
rect 46067 2400 46112 2428
rect 46106 2388 46112 2400
rect 46164 2388 46170 2440
rect 48041 2431 48099 2437
rect 48041 2397 48053 2431
rect 48087 2428 48099 2431
rect 48608 2428 48636 2527
rect 52546 2524 52552 2536
rect 52604 2524 52610 2576
rect 56137 2499 56195 2505
rect 56137 2496 56149 2499
rect 48087 2400 48636 2428
rect 48700 2468 56149 2496
rect 48087 2397 48099 2400
rect 48041 2391 48099 2397
rect 48700 2360 48728 2468
rect 56137 2465 56149 2468
rect 56183 2465 56195 2499
rect 56137 2459 56195 2465
rect 50617 2431 50675 2437
rect 50617 2397 50629 2431
rect 50663 2428 50675 2431
rect 51166 2428 51172 2440
rect 50663 2400 51172 2428
rect 50663 2397 50675 2400
rect 50617 2391 50675 2397
rect 51166 2388 51172 2400
rect 51224 2388 51230 2440
rect 52730 2428 52736 2440
rect 52691 2400 52736 2428
rect 52730 2388 52736 2400
rect 52788 2388 52794 2440
rect 54202 2388 54208 2440
rect 54260 2428 54266 2440
rect 54665 2431 54723 2437
rect 54665 2428 54677 2431
rect 54260 2400 54677 2428
rect 54260 2388 54266 2400
rect 54665 2397 54677 2400
rect 54711 2428 54723 2431
rect 55309 2431 55367 2437
rect 55309 2428 55321 2431
rect 54711 2400 55321 2428
rect 54711 2397 54723 2400
rect 54665 2391 54723 2397
rect 55309 2397 55321 2400
rect 55355 2397 55367 2431
rect 55309 2391 55367 2397
rect 56042 2388 56048 2440
rect 56100 2428 56106 2440
rect 56413 2431 56471 2437
rect 56413 2428 56425 2431
rect 56100 2400 56425 2428
rect 56100 2388 56106 2400
rect 56413 2397 56425 2400
rect 56459 2397 56471 2431
rect 57882 2428 57888 2440
rect 57843 2400 57888 2428
rect 56413 2391 56471 2397
rect 57882 2388 57888 2400
rect 57940 2388 57946 2440
rect 45526 2332 48728 2360
rect 49786 2320 49792 2372
rect 49844 2360 49850 2372
rect 54113 2363 54171 2369
rect 54113 2360 54125 2363
rect 49844 2332 54125 2360
rect 49844 2320 49850 2332
rect 54113 2329 54125 2332
rect 54159 2329 54171 2363
rect 57238 2360 57244 2372
rect 57199 2332 57244 2360
rect 54113 2323 54171 2329
rect 57238 2320 57244 2332
rect 57296 2320 57302 2372
rect 33045 2295 33103 2301
rect 33045 2261 33057 2295
rect 33091 2261 33103 2295
rect 34146 2292 34152 2304
rect 34107 2264 34152 2292
rect 33045 2255 33103 2261
rect 34146 2252 34152 2264
rect 34204 2252 34210 2304
rect 37550 2292 37556 2304
rect 37511 2264 37556 2292
rect 37550 2252 37556 2264
rect 37608 2252 37614 2304
rect 38010 2252 38016 2304
rect 38068 2292 38074 2304
rect 38289 2295 38347 2301
rect 38289 2292 38301 2295
rect 38068 2264 38301 2292
rect 38068 2252 38074 2264
rect 38289 2261 38301 2264
rect 38335 2261 38347 2295
rect 38289 2255 38347 2261
rect 40034 2252 40040 2304
rect 40092 2292 40098 2304
rect 40865 2295 40923 2301
rect 40865 2292 40877 2295
rect 40092 2264 40877 2292
rect 40092 2252 40098 2264
rect 40865 2261 40877 2264
rect 40911 2261 40923 2295
rect 41874 2292 41880 2304
rect 41835 2264 41880 2292
rect 40865 2255 40923 2261
rect 41874 2252 41880 2264
rect 41932 2252 41938 2304
rect 43346 2292 43352 2304
rect 43307 2264 43352 2292
rect 43346 2252 43352 2264
rect 43404 2252 43410 2304
rect 43806 2252 43812 2304
rect 43864 2292 43870 2304
rect 44085 2295 44143 2301
rect 44085 2292 44097 2295
rect 43864 2264 44097 2292
rect 43864 2252 43870 2264
rect 44085 2261 44097 2264
rect 44131 2261 44143 2295
rect 44085 2255 44143 2261
rect 45738 2252 45744 2304
rect 45796 2292 45802 2304
rect 45925 2295 45983 2301
rect 45925 2292 45937 2295
rect 45796 2264 45937 2292
rect 45796 2252 45802 2264
rect 45925 2261 45937 2264
rect 45971 2261 45983 2295
rect 45925 2255 45983 2261
rect 47670 2252 47676 2304
rect 47728 2292 47734 2304
rect 47857 2295 47915 2301
rect 47857 2292 47869 2295
rect 47728 2264 47869 2292
rect 47728 2252 47734 2264
rect 47857 2261 47869 2264
rect 47903 2261 47915 2295
rect 47857 2255 47915 2261
rect 50154 2252 50160 2304
rect 50212 2292 50218 2304
rect 50433 2295 50491 2301
rect 50433 2292 50445 2295
rect 50212 2264 50445 2292
rect 50212 2252 50218 2264
rect 50433 2261 50445 2264
rect 50479 2261 50491 2295
rect 50433 2255 50491 2261
rect 52178 2252 52184 2304
rect 52236 2292 52242 2304
rect 52917 2295 52975 2301
rect 52917 2292 52929 2295
rect 52236 2264 52929 2292
rect 52236 2252 52242 2264
rect 52917 2261 52929 2264
rect 52963 2261 52975 2295
rect 52917 2255 52975 2261
rect 57974 2252 57980 2304
rect 58032 2292 58038 2304
rect 58069 2295 58127 2301
rect 58069 2292 58081 2295
rect 58032 2264 58081 2292
rect 58032 2252 58038 2264
rect 58069 2261 58081 2264
rect 58115 2261 58127 2295
rect 58069 2255 58127 2261
rect 1104 2202 58880 2224
rect 1104 2150 19574 2202
rect 19626 2150 19638 2202
rect 19690 2150 19702 2202
rect 19754 2150 19766 2202
rect 19818 2150 19830 2202
rect 19882 2150 50294 2202
rect 50346 2150 50358 2202
rect 50410 2150 50422 2202
rect 50474 2150 50486 2202
rect 50538 2150 50550 2202
rect 50602 2150 58880 2202
rect 1104 2128 58880 2150
rect 5166 2048 5172 2100
rect 5224 2088 5230 2100
rect 37550 2088 37556 2100
rect 5224 2060 37556 2088
rect 5224 2048 5230 2060
rect 37550 2048 37556 2060
rect 37608 2048 37614 2100
rect 48498 2048 48504 2100
rect 48556 2088 48562 2100
rect 54570 2088 54576 2100
rect 48556 2060 54576 2088
rect 48556 2048 48562 2060
rect 54570 2048 54576 2060
rect 54628 2048 54634 2100
rect 12526 1980 12532 2032
rect 12584 2020 12590 2032
rect 46474 2020 46480 2032
rect 12584 1992 46480 2020
rect 12584 1980 12590 1992
rect 46474 1980 46480 1992
rect 46532 1980 46538 2032
rect 18414 1912 18420 1964
rect 18472 1952 18478 1964
rect 26602 1952 26608 1964
rect 18472 1924 26608 1952
rect 18472 1912 18478 1924
rect 26602 1912 26608 1924
rect 26660 1912 26666 1964
rect 42702 1912 42708 1964
rect 42760 1952 42766 1964
rect 48774 1952 48780 1964
rect 42760 1924 48780 1952
rect 42760 1912 42766 1924
rect 48774 1912 48780 1924
rect 48832 1912 48838 1964
rect 14182 1844 14188 1896
rect 14240 1884 14246 1896
rect 30098 1884 30104 1896
rect 14240 1856 30104 1884
rect 14240 1844 14246 1856
rect 30098 1844 30104 1856
rect 30156 1844 30162 1896
rect 20162 1776 20168 1828
rect 20220 1816 20226 1828
rect 43346 1816 43352 1828
rect 20220 1788 43352 1816
rect 20220 1776 20226 1788
rect 43346 1776 43352 1788
rect 43404 1776 43410 1828
rect 26234 1708 26240 1760
rect 26292 1748 26298 1760
rect 26970 1748 26976 1760
rect 26292 1720 26976 1748
rect 26292 1708 26298 1720
rect 26970 1708 26976 1720
rect 27028 1708 27034 1760
rect 27522 1708 27528 1760
rect 27580 1748 27586 1760
rect 49786 1748 49792 1760
rect 27580 1720 49792 1748
rect 27580 1708 27586 1720
rect 49786 1708 49792 1720
rect 49844 1708 49850 1760
<< via1 >>
rect 37556 37612 37608 37664
rect 39120 37612 39172 37664
rect 4214 37510 4266 37562
rect 4278 37510 4330 37562
rect 4342 37510 4394 37562
rect 4406 37510 4458 37562
rect 4470 37510 4522 37562
rect 34934 37510 34986 37562
rect 34998 37510 35050 37562
rect 35062 37510 35114 37562
rect 35126 37510 35178 37562
rect 35190 37510 35242 37562
rect 37556 37408 37608 37460
rect 37648 37408 37700 37460
rect 48596 37408 48648 37460
rect 5724 37340 5776 37392
rect 23848 37383 23900 37392
rect 23848 37349 23857 37383
rect 23857 37349 23891 37383
rect 23891 37349 23900 37383
rect 23848 37340 23900 37349
rect 4620 37272 4672 37324
rect 12256 37272 12308 37324
rect 2412 37247 2464 37256
rect 2412 37213 2421 37247
rect 2421 37213 2455 37247
rect 2455 37213 2464 37247
rect 2412 37204 2464 37213
rect 3884 37204 3936 37256
rect 5816 37204 5868 37256
rect 7748 37204 7800 37256
rect 9680 37204 9732 37256
rect 14188 37272 14240 37324
rect 16672 37247 16724 37256
rect 7104 37136 7156 37188
rect 16672 37213 16681 37247
rect 16681 37213 16715 37247
rect 16715 37213 16724 37247
rect 16672 37204 16724 37213
rect 20 37068 72 37120
rect 1952 37068 2004 37120
rect 5908 37068 5960 37120
rect 8024 37111 8076 37120
rect 8024 37077 8033 37111
rect 8033 37077 8067 37111
rect 8067 37077 8076 37111
rect 8024 37068 8076 37077
rect 11520 37068 11572 37120
rect 16580 37068 16632 37120
rect 18052 37068 18104 37120
rect 19984 37204 20036 37256
rect 28908 37272 28960 37324
rect 30288 37272 30340 37324
rect 20260 37136 20312 37188
rect 22192 37136 22244 37188
rect 25780 37204 25832 37256
rect 28356 37204 28408 37256
rect 46756 37340 46808 37392
rect 47032 37272 47084 37324
rect 32588 37247 32640 37256
rect 32588 37213 32597 37247
rect 32597 37213 32631 37247
rect 32631 37213 32640 37247
rect 32588 37204 32640 37213
rect 34152 37204 34204 37256
rect 35808 37204 35860 37256
rect 36176 37204 36228 37256
rect 37188 37204 37240 37256
rect 39028 37247 39080 37256
rect 39028 37213 39037 37247
rect 39037 37213 39071 37247
rect 39071 37213 39080 37247
rect 39028 37204 39080 37213
rect 39120 37247 39172 37256
rect 39120 37213 39129 37247
rect 39129 37213 39163 37247
rect 39163 37213 39172 37247
rect 40132 37247 40184 37256
rect 39120 37204 39172 37213
rect 40132 37213 40141 37247
rect 40141 37213 40175 37247
rect 40175 37213 40184 37247
rect 40132 37204 40184 37213
rect 41052 37204 41104 37256
rect 41880 37204 41932 37256
rect 42524 37204 42576 37256
rect 28632 37136 28684 37188
rect 34796 37179 34848 37188
rect 34796 37145 34805 37179
rect 34805 37145 34839 37179
rect 34839 37145 34848 37179
rect 34796 37136 34848 37145
rect 35624 37179 35676 37188
rect 22284 37111 22336 37120
rect 22284 37077 22293 37111
rect 22293 37077 22327 37111
rect 22327 37077 22336 37111
rect 22284 37068 22336 37077
rect 24584 37111 24636 37120
rect 24584 37077 24593 37111
rect 24593 37077 24627 37111
rect 24627 37077 24636 37111
rect 24584 37068 24636 37077
rect 26148 37068 26200 37120
rect 32220 37068 32272 37120
rect 34704 37068 34756 37120
rect 35624 37145 35633 37179
rect 35633 37145 35667 37179
rect 35667 37145 35676 37179
rect 35624 37136 35676 37145
rect 35532 37068 35584 37120
rect 38016 37136 38068 37188
rect 47584 37204 47636 37256
rect 48412 37204 48464 37256
rect 48964 37247 49016 37256
rect 48964 37213 48973 37247
rect 48973 37213 49007 37247
rect 49007 37213 49016 37247
rect 48964 37204 49016 37213
rect 50252 37204 50304 37256
rect 52552 37204 52604 37256
rect 54208 37247 54260 37256
rect 54208 37213 54217 37247
rect 54217 37213 54251 37247
rect 54251 37213 54260 37247
rect 54208 37204 54260 37213
rect 56048 37204 56100 37256
rect 57980 37204 58032 37256
rect 38292 37068 38344 37120
rect 39212 37068 39264 37120
rect 40040 37068 40092 37120
rect 43720 37136 43772 37188
rect 46112 37136 46164 37188
rect 42616 37068 42668 37120
rect 46572 37068 46624 37120
rect 46940 37136 46992 37188
rect 48228 37136 48280 37188
rect 56692 37179 56744 37188
rect 56692 37145 56701 37179
rect 56701 37145 56735 37179
rect 56735 37145 56744 37179
rect 56692 37136 56744 37145
rect 50068 37068 50120 37120
rect 50712 37111 50764 37120
rect 50712 37077 50721 37111
rect 50721 37077 50755 37111
rect 50755 37077 50764 37111
rect 50712 37068 50764 37077
rect 52184 37068 52236 37120
rect 54116 37068 54168 37120
rect 56600 37068 56652 37120
rect 58164 37068 58216 37120
rect 59912 37068 59964 37120
rect 19574 36966 19626 37018
rect 19638 36966 19690 37018
rect 19702 36966 19754 37018
rect 19766 36966 19818 37018
rect 19830 36966 19882 37018
rect 50294 36966 50346 37018
rect 50358 36966 50410 37018
rect 50422 36966 50474 37018
rect 50486 36966 50538 37018
rect 50550 36966 50602 37018
rect 1492 36907 1544 36916
rect 1492 36873 1501 36907
rect 1501 36873 1535 36907
rect 1535 36873 1544 36907
rect 1492 36864 1544 36873
rect 3884 36864 3936 36916
rect 4068 36864 4120 36916
rect 24584 36864 24636 36916
rect 32404 36864 32456 36916
rect 37188 36864 37240 36916
rect 39028 36864 39080 36916
rect 14188 36839 14240 36848
rect 14188 36805 14197 36839
rect 14197 36805 14231 36839
rect 14231 36805 14240 36839
rect 14188 36796 14240 36805
rect 26516 36796 26568 36848
rect 28080 36839 28132 36848
rect 2044 36728 2096 36780
rect 6736 36728 6788 36780
rect 7472 36771 7524 36780
rect 7472 36737 7481 36771
rect 7481 36737 7515 36771
rect 7515 36737 7524 36771
rect 7472 36728 7524 36737
rect 8300 36771 8352 36780
rect 8300 36737 8309 36771
rect 8309 36737 8343 36771
rect 8343 36737 8352 36771
rect 8300 36728 8352 36737
rect 8576 36771 8628 36780
rect 8576 36737 8585 36771
rect 8585 36737 8619 36771
rect 8619 36737 8628 36771
rect 8576 36728 8628 36737
rect 21272 36728 21324 36780
rect 23480 36728 23532 36780
rect 23848 36728 23900 36780
rect 5816 36703 5868 36712
rect 5816 36669 5825 36703
rect 5825 36669 5859 36703
rect 5859 36669 5868 36703
rect 5816 36660 5868 36669
rect 7104 36703 7156 36712
rect 7104 36669 7113 36703
rect 7113 36669 7147 36703
rect 7147 36669 7156 36703
rect 7104 36660 7156 36669
rect 19432 36660 19484 36712
rect 21732 36660 21784 36712
rect 24400 36660 24452 36712
rect 25688 36703 25740 36712
rect 25688 36669 25697 36703
rect 25697 36669 25731 36703
rect 25731 36669 25740 36703
rect 25688 36660 25740 36669
rect 26424 36660 26476 36712
rect 28080 36805 28089 36839
rect 28089 36805 28123 36839
rect 28123 36805 28132 36839
rect 28080 36796 28132 36805
rect 27896 36728 27948 36780
rect 31300 36728 31352 36780
rect 34704 36771 34756 36780
rect 34704 36737 34713 36771
rect 34713 36737 34747 36771
rect 34747 36737 34756 36771
rect 34704 36728 34756 36737
rect 34796 36728 34848 36780
rect 35532 36771 35584 36780
rect 35532 36737 35541 36771
rect 35541 36737 35575 36771
rect 35575 36737 35584 36771
rect 35532 36728 35584 36737
rect 38292 36771 38344 36780
rect 38292 36737 38301 36771
rect 38301 36737 38335 36771
rect 38335 36737 38344 36771
rect 38292 36728 38344 36737
rect 31576 36660 31628 36712
rect 33416 36660 33468 36712
rect 23480 36592 23532 36644
rect 30840 36592 30892 36644
rect 33600 36592 33652 36644
rect 40132 36864 40184 36916
rect 47400 36864 47452 36916
rect 47584 36907 47636 36916
rect 47584 36873 47593 36907
rect 47593 36873 47627 36907
rect 47627 36873 47636 36907
rect 47584 36864 47636 36873
rect 48228 36864 48280 36916
rect 48964 36907 49016 36916
rect 48964 36873 48973 36907
rect 48973 36873 49007 36907
rect 49007 36873 49016 36907
rect 48964 36864 49016 36873
rect 50160 36864 50212 36916
rect 57980 36864 58032 36916
rect 41880 36771 41932 36780
rect 39212 36660 39264 36712
rect 40132 36660 40184 36712
rect 41880 36737 41889 36771
rect 41889 36737 41923 36771
rect 41923 36737 41932 36771
rect 41880 36728 41932 36737
rect 46388 36796 46440 36848
rect 57888 36796 57940 36848
rect 42708 36728 42760 36780
rect 43720 36771 43772 36780
rect 43720 36737 43729 36771
rect 43729 36737 43763 36771
rect 43763 36737 43772 36771
rect 43720 36728 43772 36737
rect 46112 36771 46164 36780
rect 46112 36737 46121 36771
rect 46121 36737 46155 36771
rect 46155 36737 46164 36771
rect 46112 36728 46164 36737
rect 46572 36771 46624 36780
rect 46572 36737 46581 36771
rect 46581 36737 46615 36771
rect 46615 36737 46624 36771
rect 46572 36728 46624 36737
rect 47124 36728 47176 36780
rect 42616 36660 42668 36712
rect 47676 36660 47728 36712
rect 56600 36660 56652 36712
rect 6644 36524 6696 36576
rect 29092 36567 29144 36576
rect 29092 36533 29101 36567
rect 29101 36533 29135 36567
rect 29135 36533 29144 36567
rect 29092 36524 29144 36533
rect 30196 36567 30248 36576
rect 30196 36533 30205 36567
rect 30205 36533 30239 36567
rect 30239 36533 30248 36567
rect 30196 36524 30248 36533
rect 32496 36524 32548 36576
rect 35808 36567 35860 36576
rect 35808 36533 35817 36567
rect 35817 36533 35851 36567
rect 35851 36533 35860 36567
rect 35808 36524 35860 36533
rect 36452 36524 36504 36576
rect 39304 36524 39356 36576
rect 39396 36567 39448 36576
rect 39396 36533 39405 36567
rect 39405 36533 39439 36567
rect 39439 36533 39448 36567
rect 39396 36524 39448 36533
rect 40316 36524 40368 36576
rect 41420 36567 41472 36576
rect 41420 36533 41429 36567
rect 41429 36533 41463 36567
rect 41463 36533 41472 36567
rect 41420 36524 41472 36533
rect 42616 36567 42668 36576
rect 42616 36533 42625 36567
rect 42625 36533 42659 36567
rect 42659 36533 42668 36567
rect 42616 36524 42668 36533
rect 42984 36567 43036 36576
rect 42984 36533 42993 36567
rect 42993 36533 43027 36567
rect 43027 36533 43036 36567
rect 42984 36524 43036 36533
rect 56600 36524 56652 36576
rect 4214 36422 4266 36474
rect 4278 36422 4330 36474
rect 4342 36422 4394 36474
rect 4406 36422 4458 36474
rect 4470 36422 4522 36474
rect 34934 36422 34986 36474
rect 34998 36422 35050 36474
rect 35062 36422 35114 36474
rect 35126 36422 35178 36474
rect 35190 36422 35242 36474
rect 8300 36320 8352 36372
rect 8944 36363 8996 36372
rect 8944 36329 8953 36363
rect 8953 36329 8987 36363
rect 8987 36329 8996 36363
rect 8944 36320 8996 36329
rect 19432 36363 19484 36372
rect 19432 36329 19441 36363
rect 19441 36329 19475 36363
rect 19475 36329 19484 36363
rect 19432 36320 19484 36329
rect 21732 36363 21784 36372
rect 21732 36329 21741 36363
rect 21741 36329 21775 36363
rect 21775 36329 21784 36363
rect 21732 36320 21784 36329
rect 23848 36363 23900 36372
rect 23848 36329 23857 36363
rect 23857 36329 23891 36363
rect 23891 36329 23900 36363
rect 23848 36320 23900 36329
rect 6644 36252 6696 36304
rect 8576 36252 8628 36304
rect 21272 36252 21324 36304
rect 1676 36159 1728 36168
rect 1676 36125 1685 36159
rect 1685 36125 1719 36159
rect 1719 36125 1728 36159
rect 1676 36116 1728 36125
rect 8024 36116 8076 36168
rect 20076 36184 20128 36236
rect 8852 36116 8904 36168
rect 19248 36159 19300 36168
rect 19248 36125 19257 36159
rect 19257 36125 19291 36159
rect 19291 36125 19300 36159
rect 19248 36116 19300 36125
rect 19340 36116 19392 36168
rect 21272 36159 21324 36168
rect 21272 36125 21281 36159
rect 21281 36125 21315 36159
rect 21315 36125 21324 36159
rect 21272 36116 21324 36125
rect 22100 36116 22152 36168
rect 25688 36320 25740 36372
rect 26424 36363 26476 36372
rect 26424 36329 26433 36363
rect 26433 36329 26467 36363
rect 26467 36329 26476 36363
rect 26424 36320 26476 36329
rect 28632 36363 28684 36372
rect 28632 36329 28641 36363
rect 28641 36329 28675 36363
rect 28675 36329 28684 36363
rect 28632 36320 28684 36329
rect 31576 36363 31628 36372
rect 31576 36329 31585 36363
rect 31585 36329 31619 36363
rect 31619 36329 31628 36363
rect 31576 36320 31628 36329
rect 23664 36159 23716 36168
rect 23664 36125 23673 36159
rect 23673 36125 23707 36159
rect 23707 36125 23716 36159
rect 23664 36116 23716 36125
rect 23848 36159 23900 36168
rect 23848 36125 23857 36159
rect 23857 36125 23891 36159
rect 23891 36125 23900 36159
rect 24400 36159 24452 36168
rect 23848 36116 23900 36125
rect 24400 36125 24409 36159
rect 24409 36125 24443 36159
rect 24443 36125 24452 36159
rect 24400 36116 24452 36125
rect 24492 36159 24544 36168
rect 24492 36125 24501 36159
rect 24501 36125 24535 36159
rect 24535 36125 24544 36159
rect 24492 36116 24544 36125
rect 27896 36252 27948 36304
rect 39028 36320 39080 36372
rect 34796 36252 34848 36304
rect 35624 36252 35676 36304
rect 26516 36116 26568 36168
rect 28448 36159 28500 36168
rect 28448 36125 28457 36159
rect 28457 36125 28491 36159
rect 28491 36125 28500 36159
rect 28448 36116 28500 36125
rect 28632 36159 28684 36168
rect 28632 36125 28641 36159
rect 28641 36125 28675 36159
rect 28675 36125 28684 36159
rect 28632 36116 28684 36125
rect 29092 36116 29144 36168
rect 32496 36227 32548 36236
rect 32496 36193 32505 36227
rect 32505 36193 32539 36227
rect 32539 36193 32548 36227
rect 32496 36184 32548 36193
rect 30840 36159 30892 36168
rect 30840 36125 30849 36159
rect 30849 36125 30883 36159
rect 30883 36125 30892 36159
rect 30840 36116 30892 36125
rect 31300 36159 31352 36168
rect 31300 36125 31309 36159
rect 31309 36125 31343 36159
rect 31343 36125 31352 36159
rect 31300 36116 31352 36125
rect 32404 36159 32456 36168
rect 32404 36125 32413 36159
rect 32413 36125 32447 36159
rect 32447 36125 32456 36159
rect 32404 36116 32456 36125
rect 33416 36116 33468 36168
rect 34704 36116 34756 36168
rect 1492 36023 1544 36032
rect 1492 35989 1501 36023
rect 1501 35989 1535 36023
rect 1535 35989 1544 36023
rect 1492 35980 1544 35989
rect 8760 35980 8812 36032
rect 23664 35980 23716 36032
rect 24492 35980 24544 36032
rect 29644 36023 29696 36032
rect 29644 35989 29653 36023
rect 29653 35989 29687 36023
rect 29687 35989 29696 36023
rect 29644 35980 29696 35989
rect 31760 36023 31812 36032
rect 31760 35989 31769 36023
rect 31769 35989 31803 36023
rect 31803 35989 31812 36023
rect 33232 36023 33284 36032
rect 31760 35980 31812 35989
rect 33232 35989 33241 36023
rect 33241 35989 33275 36023
rect 33275 35989 33284 36023
rect 33232 35980 33284 35989
rect 33600 36091 33652 36100
rect 33600 36057 33609 36091
rect 33609 36057 33643 36091
rect 33643 36057 33652 36091
rect 35532 36091 35584 36100
rect 33600 36048 33652 36057
rect 35532 36057 35541 36091
rect 35541 36057 35575 36091
rect 35575 36057 35584 36091
rect 35532 36048 35584 36057
rect 36452 36159 36504 36168
rect 36452 36125 36461 36159
rect 36461 36125 36495 36159
rect 36495 36125 36504 36159
rect 36452 36116 36504 36125
rect 38108 36227 38160 36236
rect 38108 36193 38117 36227
rect 38117 36193 38151 36227
rect 38151 36193 38160 36227
rect 38108 36184 38160 36193
rect 41420 36320 41472 36372
rect 47400 36320 47452 36372
rect 39304 36252 39356 36304
rect 46112 36252 46164 36304
rect 41420 36227 41472 36236
rect 41420 36193 41429 36227
rect 41429 36193 41463 36227
rect 41463 36193 41472 36227
rect 41420 36184 41472 36193
rect 49056 36227 49108 36236
rect 49056 36193 49065 36227
rect 49065 36193 49099 36227
rect 49099 36193 49108 36227
rect 49056 36184 49108 36193
rect 38200 36159 38252 36168
rect 38200 36125 38209 36159
rect 38209 36125 38243 36159
rect 38243 36125 38252 36159
rect 38200 36116 38252 36125
rect 38292 36116 38344 36168
rect 40316 36159 40368 36168
rect 40316 36125 40325 36159
rect 40325 36125 40359 36159
rect 40359 36125 40368 36159
rect 40316 36116 40368 36125
rect 42984 36159 43036 36168
rect 41880 36048 41932 36100
rect 42984 36125 42993 36159
rect 42993 36125 43027 36159
rect 43027 36125 43036 36159
rect 42984 36116 43036 36125
rect 47124 36159 47176 36168
rect 47124 36125 47133 36159
rect 47133 36125 47167 36159
rect 47167 36125 47176 36159
rect 47124 36116 47176 36125
rect 47676 36159 47728 36168
rect 47676 36125 47685 36159
rect 47685 36125 47719 36159
rect 47719 36125 47728 36159
rect 47676 36116 47728 36125
rect 48964 36159 49016 36168
rect 48964 36125 48973 36159
rect 48973 36125 49007 36159
rect 49007 36125 49016 36159
rect 48964 36116 49016 36125
rect 58164 36159 58216 36168
rect 58164 36125 58173 36159
rect 58173 36125 58207 36159
rect 58207 36125 58216 36159
rect 58164 36116 58216 36125
rect 44640 36048 44692 36100
rect 46572 36048 46624 36100
rect 57796 36048 57848 36100
rect 39120 36023 39172 36032
rect 39120 35989 39129 36023
rect 39129 35989 39163 36023
rect 39163 35989 39172 36023
rect 39120 35980 39172 35989
rect 40132 35980 40184 36032
rect 19574 35878 19626 35930
rect 19638 35878 19690 35930
rect 19702 35878 19754 35930
rect 19766 35878 19818 35930
rect 19830 35878 19882 35930
rect 50294 35878 50346 35930
rect 50358 35878 50410 35930
rect 50422 35878 50474 35930
rect 50486 35878 50538 35930
rect 50550 35878 50602 35930
rect 6644 35819 6696 35828
rect 6644 35785 6653 35819
rect 6653 35785 6687 35819
rect 6687 35785 6696 35819
rect 6644 35776 6696 35785
rect 6736 35819 6788 35828
rect 6736 35785 6745 35819
rect 6745 35785 6779 35819
rect 6779 35785 6788 35819
rect 6736 35776 6788 35785
rect 16580 35776 16632 35828
rect 17776 35776 17828 35828
rect 7012 35708 7064 35760
rect 7472 35708 7524 35760
rect 8024 35751 8076 35760
rect 8024 35717 8033 35751
rect 8033 35717 8067 35751
rect 8067 35717 8076 35751
rect 8024 35708 8076 35717
rect 18144 35708 18196 35760
rect 19248 35708 19300 35760
rect 7748 35640 7800 35692
rect 8116 35683 8168 35692
rect 8116 35649 8125 35683
rect 8125 35649 8159 35683
rect 8159 35649 8168 35683
rect 8116 35640 8168 35649
rect 8300 35683 8352 35692
rect 8300 35649 8309 35683
rect 8309 35649 8343 35683
rect 8343 35649 8352 35683
rect 8300 35640 8352 35649
rect 8760 35683 8812 35692
rect 8760 35649 8769 35683
rect 8769 35649 8803 35683
rect 8803 35649 8812 35683
rect 8760 35640 8812 35649
rect 8944 35683 8996 35692
rect 8944 35649 8953 35683
rect 8953 35649 8987 35683
rect 8987 35649 8996 35683
rect 8944 35640 8996 35649
rect 11704 35683 11756 35692
rect 11704 35649 11713 35683
rect 11713 35649 11747 35683
rect 11747 35649 11756 35683
rect 11704 35640 11756 35649
rect 11888 35683 11940 35692
rect 11888 35649 11897 35683
rect 11897 35649 11931 35683
rect 11931 35649 11940 35683
rect 11888 35640 11940 35649
rect 22100 35708 22152 35760
rect 23848 35708 23900 35760
rect 8852 35572 8904 35624
rect 5540 35504 5592 35556
rect 12348 35504 12400 35556
rect 19340 35572 19392 35624
rect 21088 35640 21140 35692
rect 28724 35776 28776 35828
rect 38200 35776 38252 35828
rect 40132 35819 40184 35828
rect 40132 35785 40141 35819
rect 40141 35785 40175 35819
rect 40175 35785 40184 35819
rect 40132 35776 40184 35785
rect 47124 35776 47176 35828
rect 49056 35776 49108 35828
rect 58164 35819 58216 35828
rect 58164 35785 58173 35819
rect 58173 35785 58207 35819
rect 58207 35785 58216 35819
rect 58164 35776 58216 35785
rect 27988 35708 28040 35760
rect 50712 35708 50764 35760
rect 29644 35640 29696 35692
rect 30196 35640 30248 35692
rect 31760 35640 31812 35692
rect 32404 35640 32456 35692
rect 33232 35640 33284 35692
rect 45100 35640 45152 35692
rect 49424 35683 49476 35692
rect 24952 35572 25004 35624
rect 29092 35572 29144 35624
rect 43628 35572 43680 35624
rect 49424 35649 49433 35683
rect 49433 35649 49467 35683
rect 49467 35649 49476 35683
rect 49424 35640 49476 35649
rect 49976 35572 50028 35624
rect 23664 35504 23716 35556
rect 28632 35547 28684 35556
rect 28632 35513 28641 35547
rect 28641 35513 28675 35547
rect 28675 35513 28684 35547
rect 28632 35504 28684 35513
rect 7932 35436 7984 35488
rect 8852 35436 8904 35488
rect 12440 35436 12492 35488
rect 18696 35436 18748 35488
rect 20076 35436 20128 35488
rect 28356 35436 28408 35488
rect 30196 35479 30248 35488
rect 30196 35445 30205 35479
rect 30205 35445 30239 35479
rect 30239 35445 30248 35479
rect 30196 35436 30248 35445
rect 41052 35479 41104 35488
rect 41052 35445 41061 35479
rect 41061 35445 41095 35479
rect 41095 35445 41104 35479
rect 41052 35436 41104 35445
rect 4214 35334 4266 35386
rect 4278 35334 4330 35386
rect 4342 35334 4394 35386
rect 4406 35334 4458 35386
rect 4470 35334 4522 35386
rect 34934 35334 34986 35386
rect 34998 35334 35050 35386
rect 35062 35334 35114 35386
rect 35126 35334 35178 35386
rect 35190 35334 35242 35386
rect 7012 35232 7064 35284
rect 7748 35275 7800 35284
rect 7748 35241 7757 35275
rect 7757 35241 7791 35275
rect 7791 35241 7800 35275
rect 7748 35232 7800 35241
rect 9588 35275 9640 35284
rect 7012 35139 7064 35148
rect 7012 35105 7021 35139
rect 7021 35105 7055 35139
rect 7055 35105 7064 35139
rect 7012 35096 7064 35105
rect 8300 35096 8352 35148
rect 9588 35241 9597 35275
rect 9597 35241 9631 35275
rect 9631 35241 9640 35275
rect 9588 35232 9640 35241
rect 11888 35232 11940 35284
rect 16580 35275 16632 35284
rect 16580 35241 16589 35275
rect 16589 35241 16623 35275
rect 16623 35241 16632 35275
rect 16580 35232 16632 35241
rect 18328 35232 18380 35284
rect 18696 35275 18748 35284
rect 18696 35241 18705 35275
rect 18705 35241 18739 35275
rect 18739 35241 18748 35275
rect 18696 35232 18748 35241
rect 22100 35232 22152 35284
rect 12440 35096 12492 35148
rect 7932 35071 7984 35080
rect 7932 35037 7941 35071
rect 7941 35037 7975 35071
rect 7975 35037 7984 35071
rect 7932 35028 7984 35037
rect 8024 35028 8076 35080
rect 11520 35071 11572 35080
rect 11520 35037 11529 35071
rect 11529 35037 11563 35071
rect 11563 35037 11572 35071
rect 11520 35028 11572 35037
rect 12164 35071 12216 35080
rect 12164 35037 12173 35071
rect 12173 35037 12207 35071
rect 12207 35037 12216 35071
rect 12164 35028 12216 35037
rect 12716 35071 12768 35080
rect 12716 35037 12725 35071
rect 12725 35037 12759 35071
rect 12759 35037 12768 35071
rect 12716 35028 12768 35037
rect 12900 34960 12952 35012
rect 16580 34960 16632 35012
rect 17868 34960 17920 35012
rect 12532 34935 12584 34944
rect 12532 34901 12541 34935
rect 12541 34901 12575 34935
rect 12575 34901 12584 34935
rect 12532 34892 12584 34901
rect 18420 34892 18472 34944
rect 20812 35028 20864 35080
rect 23480 35071 23532 35080
rect 21272 34960 21324 35012
rect 23480 35037 23489 35071
rect 23489 35037 23523 35071
rect 23523 35037 23532 35071
rect 23480 35028 23532 35037
rect 27896 35232 27948 35284
rect 28448 35232 28500 35284
rect 32588 35232 32640 35284
rect 24492 35164 24544 35216
rect 34704 35207 34756 35216
rect 25136 35071 25188 35080
rect 25136 35037 25145 35071
rect 25145 35037 25179 35071
rect 25179 35037 25188 35071
rect 25136 35028 25188 35037
rect 34704 35173 34713 35207
rect 34713 35173 34747 35207
rect 34747 35173 34756 35207
rect 34704 35164 34756 35173
rect 35992 35232 36044 35284
rect 37372 35232 37424 35284
rect 43628 35275 43680 35284
rect 43628 35241 43637 35275
rect 43637 35241 43671 35275
rect 43671 35241 43680 35275
rect 43628 35232 43680 35241
rect 22652 34960 22704 35012
rect 28356 35071 28408 35080
rect 22192 34892 22244 34944
rect 24952 34892 25004 34944
rect 28356 35037 28365 35071
rect 28365 35037 28399 35071
rect 28399 35037 28408 35071
rect 28356 35028 28408 35037
rect 27988 34892 28040 34944
rect 35900 35096 35952 35148
rect 37188 35096 37240 35148
rect 43260 35139 43312 35148
rect 43260 35105 43269 35139
rect 43269 35105 43303 35139
rect 43303 35105 43312 35139
rect 43260 35096 43312 35105
rect 54208 35164 54260 35216
rect 28724 35028 28776 35080
rect 35348 35028 35400 35080
rect 37464 35071 37516 35080
rect 37464 35037 37473 35071
rect 37473 35037 37507 35071
rect 37507 35037 37516 35071
rect 37464 35028 37516 35037
rect 43352 35071 43404 35080
rect 43352 35037 43361 35071
rect 43361 35037 43395 35071
rect 43395 35037 43404 35071
rect 43352 35028 43404 35037
rect 48504 35028 48556 35080
rect 49516 35096 49568 35148
rect 52184 35096 52236 35148
rect 57888 35139 57940 35148
rect 57888 35105 57897 35139
rect 57897 35105 57931 35139
rect 57931 35105 57940 35139
rect 57888 35096 57940 35105
rect 28908 34960 28960 35012
rect 40316 34960 40368 35012
rect 35992 34892 36044 34944
rect 38936 34892 38988 34944
rect 48412 34892 48464 34944
rect 49056 35028 49108 35080
rect 48688 34960 48740 35012
rect 53564 35028 53616 35080
rect 58164 35071 58216 35080
rect 58164 35037 58173 35071
rect 58173 35037 58207 35071
rect 58207 35037 58216 35071
rect 58164 35028 58216 35037
rect 49976 34892 50028 34944
rect 19574 34790 19626 34842
rect 19638 34790 19690 34842
rect 19702 34790 19754 34842
rect 19766 34790 19818 34842
rect 19830 34790 19882 34842
rect 50294 34790 50346 34842
rect 50358 34790 50410 34842
rect 50422 34790 50474 34842
rect 50486 34790 50538 34842
rect 50550 34790 50602 34842
rect 8300 34688 8352 34740
rect 18144 34688 18196 34740
rect 19340 34688 19392 34740
rect 20812 34688 20864 34740
rect 21088 34731 21140 34740
rect 21088 34697 21097 34731
rect 21097 34697 21131 34731
rect 21131 34697 21140 34731
rect 21088 34688 21140 34697
rect 22192 34688 22244 34740
rect 48596 34688 48648 34740
rect 48964 34688 49016 34740
rect 52184 34731 52236 34740
rect 52184 34697 52193 34731
rect 52193 34697 52227 34731
rect 52227 34697 52236 34731
rect 52184 34688 52236 34697
rect 53564 34731 53616 34740
rect 53564 34697 53573 34731
rect 53573 34697 53607 34731
rect 53607 34697 53616 34731
rect 53564 34688 53616 34697
rect 58164 34731 58216 34740
rect 58164 34697 58173 34731
rect 58173 34697 58207 34731
rect 58207 34697 58216 34731
rect 58164 34688 58216 34697
rect 12440 34620 12492 34672
rect 15292 34620 15344 34672
rect 16488 34620 16540 34672
rect 7840 34595 7892 34604
rect 7840 34561 7849 34595
rect 7849 34561 7883 34595
rect 7883 34561 7892 34595
rect 7840 34552 7892 34561
rect 9496 34552 9548 34604
rect 11520 34552 11572 34604
rect 12348 34595 12400 34604
rect 12348 34561 12357 34595
rect 12357 34561 12391 34595
rect 12391 34561 12400 34595
rect 12348 34552 12400 34561
rect 12532 34552 12584 34604
rect 15844 34552 15896 34604
rect 17408 34552 17460 34604
rect 17868 34552 17920 34604
rect 18328 34595 18380 34604
rect 18328 34561 18337 34595
rect 18337 34561 18371 34595
rect 18371 34561 18380 34595
rect 18328 34552 18380 34561
rect 18420 34595 18472 34604
rect 18420 34561 18429 34595
rect 18429 34561 18463 34595
rect 18463 34561 18472 34595
rect 18420 34552 18472 34561
rect 7012 34484 7064 34536
rect 7932 34484 7984 34536
rect 11612 34484 11664 34536
rect 15200 34527 15252 34536
rect 15200 34493 15209 34527
rect 15209 34493 15243 34527
rect 15243 34493 15252 34527
rect 15200 34484 15252 34493
rect 16120 34527 16172 34536
rect 16120 34493 16129 34527
rect 16129 34493 16163 34527
rect 16163 34493 16172 34527
rect 16120 34484 16172 34493
rect 11152 34416 11204 34468
rect 18328 34416 18380 34468
rect 20168 34552 20220 34604
rect 22652 34620 22704 34672
rect 24492 34620 24544 34672
rect 27896 34663 27948 34672
rect 27896 34629 27905 34663
rect 27905 34629 27939 34663
rect 27939 34629 27948 34663
rect 27896 34620 27948 34629
rect 34796 34620 34848 34672
rect 24952 34595 25004 34604
rect 24952 34561 24961 34595
rect 24961 34561 24995 34595
rect 24995 34561 25004 34595
rect 24952 34552 25004 34561
rect 25136 34552 25188 34604
rect 27804 34552 27856 34604
rect 28448 34552 28500 34604
rect 32404 34595 32456 34604
rect 32404 34561 32413 34595
rect 32413 34561 32447 34595
rect 32447 34561 32456 34595
rect 32404 34552 32456 34561
rect 32772 34595 32824 34604
rect 32772 34561 32781 34595
rect 32781 34561 32815 34595
rect 32815 34561 32824 34595
rect 32772 34552 32824 34561
rect 35992 34595 36044 34604
rect 35992 34561 36001 34595
rect 36001 34561 36035 34595
rect 36035 34561 36044 34595
rect 35992 34552 36044 34561
rect 37832 34595 37884 34604
rect 37832 34561 37841 34595
rect 37841 34561 37875 34595
rect 37875 34561 37884 34595
rect 37832 34552 37884 34561
rect 38200 34552 38252 34604
rect 38936 34595 38988 34604
rect 38936 34561 38945 34595
rect 38945 34561 38979 34595
rect 38979 34561 38988 34595
rect 38936 34552 38988 34561
rect 40040 34595 40092 34604
rect 35348 34484 35400 34536
rect 37464 34484 37516 34536
rect 38292 34484 38344 34536
rect 40040 34561 40049 34595
rect 40049 34561 40083 34595
rect 40083 34561 40092 34595
rect 40040 34552 40092 34561
rect 40132 34527 40184 34536
rect 27988 34459 28040 34468
rect 7656 34391 7708 34400
rect 7656 34357 7665 34391
rect 7665 34357 7699 34391
rect 7699 34357 7708 34391
rect 7656 34348 7708 34357
rect 14096 34348 14148 34400
rect 27988 34425 27997 34459
rect 27997 34425 28031 34459
rect 28031 34425 28040 34459
rect 27988 34416 28040 34425
rect 33600 34459 33652 34468
rect 33600 34425 33609 34459
rect 33609 34425 33643 34459
rect 33643 34425 33652 34459
rect 33600 34416 33652 34425
rect 35900 34459 35952 34468
rect 35900 34425 35909 34459
rect 35909 34425 35943 34459
rect 35943 34425 35952 34459
rect 35900 34416 35952 34425
rect 38384 34416 38436 34468
rect 40132 34493 40141 34527
rect 40141 34493 40175 34527
rect 40175 34493 40184 34527
rect 40132 34484 40184 34493
rect 40316 34620 40368 34672
rect 48688 34620 48740 34672
rect 42892 34552 42944 34604
rect 43168 34595 43220 34604
rect 43168 34561 43177 34595
rect 43177 34561 43211 34595
rect 43211 34561 43220 34595
rect 43168 34552 43220 34561
rect 48412 34552 48464 34604
rect 45100 34484 45152 34536
rect 48872 34484 48924 34536
rect 40316 34416 40368 34468
rect 43260 34416 43312 34468
rect 48504 34416 48556 34468
rect 49976 34595 50028 34604
rect 49976 34561 49985 34595
rect 49985 34561 50019 34595
rect 50019 34561 50028 34595
rect 49976 34552 50028 34561
rect 52460 34620 52512 34672
rect 49516 34484 49568 34536
rect 52184 34416 52236 34468
rect 28448 34391 28500 34400
rect 28448 34357 28457 34391
rect 28457 34357 28491 34391
rect 28491 34357 28500 34391
rect 28448 34348 28500 34357
rect 38108 34391 38160 34400
rect 38108 34357 38117 34391
rect 38117 34357 38151 34391
rect 38151 34357 38160 34391
rect 38108 34348 38160 34357
rect 49424 34348 49476 34400
rect 52644 34552 52696 34604
rect 52828 34595 52880 34604
rect 52828 34561 52837 34595
rect 52837 34561 52871 34595
rect 52871 34561 52880 34595
rect 53472 34595 53524 34604
rect 52828 34552 52880 34561
rect 53472 34561 53481 34595
rect 53481 34561 53515 34595
rect 53515 34561 53524 34595
rect 53472 34552 53524 34561
rect 52920 34348 52972 34400
rect 4214 34246 4266 34298
rect 4278 34246 4330 34298
rect 4342 34246 4394 34298
rect 4406 34246 4458 34298
rect 4470 34246 4522 34298
rect 34934 34246 34986 34298
rect 34998 34246 35050 34298
rect 35062 34246 35114 34298
rect 35126 34246 35178 34298
rect 35190 34246 35242 34298
rect 11704 34144 11756 34196
rect 15200 34187 15252 34196
rect 15200 34153 15209 34187
rect 15209 34153 15243 34187
rect 15243 34153 15252 34187
rect 15200 34144 15252 34153
rect 17408 34144 17460 34196
rect 18420 34144 18472 34196
rect 25136 34187 25188 34196
rect 25136 34153 25145 34187
rect 25145 34153 25179 34187
rect 25179 34153 25188 34187
rect 25136 34144 25188 34153
rect 27620 34144 27672 34196
rect 27896 34187 27948 34196
rect 27896 34153 27905 34187
rect 27905 34153 27939 34187
rect 27939 34153 27948 34187
rect 27896 34144 27948 34153
rect 28540 34187 28592 34196
rect 28540 34153 28549 34187
rect 28549 34153 28583 34187
rect 28583 34153 28592 34187
rect 28540 34144 28592 34153
rect 32772 34187 32824 34196
rect 11796 34076 11848 34128
rect 12164 34076 12216 34128
rect 16120 34076 16172 34128
rect 24952 34119 25004 34128
rect 24952 34085 24961 34119
rect 24961 34085 24995 34119
rect 24995 34085 25004 34119
rect 24952 34076 25004 34085
rect 28356 34076 28408 34128
rect 11888 34008 11940 34060
rect 12072 34008 12124 34060
rect 22284 34008 22336 34060
rect 22652 34051 22704 34060
rect 22652 34017 22661 34051
rect 22661 34017 22695 34051
rect 22695 34017 22704 34051
rect 22652 34008 22704 34017
rect 23388 34051 23440 34060
rect 23388 34017 23397 34051
rect 23397 34017 23431 34051
rect 23431 34017 23440 34051
rect 23388 34008 23440 34017
rect 32772 34153 32781 34187
rect 32781 34153 32815 34187
rect 32815 34153 32824 34187
rect 32772 34144 32824 34153
rect 34796 34144 34848 34196
rect 38384 34187 38436 34196
rect 38384 34153 38393 34187
rect 38393 34153 38427 34187
rect 38427 34153 38436 34187
rect 38384 34144 38436 34153
rect 40132 34144 40184 34196
rect 43168 34144 43220 34196
rect 48688 34187 48740 34196
rect 48688 34153 48697 34187
rect 48697 34153 48731 34187
rect 48731 34153 48740 34187
rect 48688 34144 48740 34153
rect 49424 34144 49476 34196
rect 38292 34119 38344 34128
rect 38292 34085 38301 34119
rect 38301 34085 38335 34119
rect 38335 34085 38344 34119
rect 38292 34076 38344 34085
rect 40224 34076 40276 34128
rect 35900 34051 35952 34060
rect 35900 34017 35909 34051
rect 35909 34017 35943 34051
rect 35943 34017 35952 34051
rect 35900 34008 35952 34017
rect 37832 34008 37884 34060
rect 7840 33940 7892 33992
rect 8208 33940 8260 33992
rect 9128 33940 9180 33992
rect 9772 33940 9824 33992
rect 11152 33940 11204 33992
rect 11612 33940 11664 33992
rect 12900 33983 12952 33992
rect 8300 33872 8352 33924
rect 9496 33915 9548 33924
rect 9496 33881 9505 33915
rect 9505 33881 9539 33915
rect 9539 33881 9548 33915
rect 9496 33872 9548 33881
rect 12900 33949 12909 33983
rect 12909 33949 12943 33983
rect 12943 33949 12952 33983
rect 12900 33940 12952 33949
rect 14188 33940 14240 33992
rect 7288 33804 7340 33856
rect 12716 33872 12768 33924
rect 13728 33872 13780 33924
rect 15292 33940 15344 33992
rect 15844 33983 15896 33992
rect 15844 33949 15853 33983
rect 15853 33949 15887 33983
rect 15887 33949 15896 33983
rect 15844 33940 15896 33949
rect 18420 33983 18472 33992
rect 18420 33949 18429 33983
rect 18429 33949 18463 33983
rect 18463 33949 18472 33983
rect 18420 33940 18472 33949
rect 18512 33915 18564 33924
rect 18512 33881 18521 33915
rect 18521 33881 18555 33915
rect 18555 33881 18564 33915
rect 18512 33872 18564 33881
rect 18328 33804 18380 33856
rect 19248 33940 19300 33992
rect 18788 33872 18840 33924
rect 23204 33983 23256 33992
rect 23204 33949 23213 33983
rect 23213 33949 23247 33983
rect 23247 33949 23256 33983
rect 23204 33940 23256 33949
rect 28264 33940 28316 33992
rect 24676 33915 24728 33924
rect 24676 33881 24685 33915
rect 24685 33881 24719 33915
rect 24719 33881 24728 33915
rect 24676 33872 24728 33881
rect 27712 33915 27764 33924
rect 27712 33881 27721 33915
rect 27721 33881 27755 33915
rect 27755 33881 27764 33915
rect 27712 33872 27764 33881
rect 27804 33872 27856 33924
rect 31116 33940 31168 33992
rect 31392 33983 31444 33992
rect 31392 33949 31401 33983
rect 31401 33949 31435 33983
rect 31435 33949 31444 33983
rect 31392 33940 31444 33949
rect 32404 33940 32456 33992
rect 35440 33940 35492 33992
rect 37188 33983 37240 33992
rect 37188 33949 37197 33983
rect 37197 33949 37231 33983
rect 37231 33949 37240 33983
rect 37188 33940 37240 33949
rect 37372 33983 37424 33992
rect 37372 33949 37381 33983
rect 37381 33949 37415 33983
rect 37415 33949 37424 33983
rect 37372 33940 37424 33949
rect 39948 33983 40000 33992
rect 39948 33949 39957 33983
rect 39957 33949 39991 33983
rect 39991 33949 40000 33983
rect 39948 33940 40000 33949
rect 40316 33940 40368 33992
rect 41788 34051 41840 34060
rect 41788 34017 41797 34051
rect 41797 34017 41831 34051
rect 41831 34017 41840 34051
rect 41788 34008 41840 34017
rect 42892 34076 42944 34128
rect 42892 33983 42944 33992
rect 35348 33915 35400 33924
rect 35348 33881 35357 33915
rect 35357 33881 35391 33915
rect 35391 33881 35400 33915
rect 35348 33872 35400 33881
rect 20168 33804 20220 33856
rect 28080 33847 28132 33856
rect 28080 33813 28089 33847
rect 28089 33813 28123 33847
rect 28123 33813 28132 33847
rect 28080 33804 28132 33813
rect 42892 33949 42901 33983
rect 42901 33949 42935 33983
rect 42935 33949 42944 33983
rect 42892 33940 42944 33949
rect 42616 33872 42668 33924
rect 43352 33940 43404 33992
rect 46940 34076 46992 34128
rect 45008 33983 45060 33992
rect 45008 33949 45017 33983
rect 45017 33949 45051 33983
rect 45051 33949 45060 33983
rect 45008 33940 45060 33949
rect 45100 33983 45152 33992
rect 45100 33949 45109 33983
rect 45109 33949 45143 33983
rect 45143 33949 45152 33983
rect 45100 33940 45152 33949
rect 48688 33940 48740 33992
rect 51264 33983 51316 33992
rect 51264 33949 51273 33983
rect 51273 33949 51307 33983
rect 51307 33949 51316 33983
rect 51264 33940 51316 33949
rect 52460 34008 52512 34060
rect 53472 34051 53524 34060
rect 53472 34017 53481 34051
rect 53481 34017 53515 34051
rect 53515 34017 53524 34051
rect 53472 34008 53524 34017
rect 52184 33983 52236 33992
rect 52184 33949 52193 33983
rect 52193 33949 52227 33983
rect 52227 33949 52236 33983
rect 52184 33940 52236 33949
rect 52920 33983 52972 33992
rect 49056 33872 49108 33924
rect 52920 33949 52929 33983
rect 52929 33949 52963 33983
rect 52963 33949 52972 33983
rect 52920 33940 52972 33949
rect 55588 33872 55640 33924
rect 43168 33804 43220 33856
rect 43352 33847 43404 33856
rect 43352 33813 43361 33847
rect 43361 33813 43395 33847
rect 43395 33813 43404 33847
rect 43352 33804 43404 33813
rect 45836 33804 45888 33856
rect 52184 33804 52236 33856
rect 19574 33702 19626 33754
rect 19638 33702 19690 33754
rect 19702 33702 19754 33754
rect 19766 33702 19818 33754
rect 19830 33702 19882 33754
rect 50294 33702 50346 33754
rect 50358 33702 50410 33754
rect 50422 33702 50474 33754
rect 50486 33702 50538 33754
rect 50550 33702 50602 33754
rect 11796 33643 11848 33652
rect 11796 33609 11805 33643
rect 11805 33609 11839 33643
rect 11839 33609 11848 33643
rect 11796 33600 11848 33609
rect 17776 33600 17828 33652
rect 27620 33643 27672 33652
rect 27620 33609 27629 33643
rect 27629 33609 27663 33643
rect 27663 33609 27672 33643
rect 27620 33600 27672 33609
rect 27804 33600 27856 33652
rect 31392 33600 31444 33652
rect 35716 33600 35768 33652
rect 1584 33464 1636 33516
rect 9128 33575 9180 33584
rect 9128 33541 9137 33575
rect 9137 33541 9171 33575
rect 9171 33541 9180 33575
rect 9128 33532 9180 33541
rect 12072 33532 12124 33584
rect 17132 33575 17184 33584
rect 17132 33541 17141 33575
rect 17141 33541 17175 33575
rect 17175 33541 17184 33575
rect 17132 33532 17184 33541
rect 23388 33532 23440 33584
rect 25320 33532 25372 33584
rect 7104 33328 7156 33380
rect 8208 33464 8260 33516
rect 8300 33464 8352 33516
rect 9772 33464 9824 33516
rect 11612 33464 11664 33516
rect 22468 33464 22520 33516
rect 23204 33507 23256 33516
rect 23204 33473 23213 33507
rect 23213 33473 23247 33507
rect 23247 33473 23256 33507
rect 23204 33464 23256 33473
rect 24676 33464 24728 33516
rect 27712 33464 27764 33516
rect 28448 33532 28500 33584
rect 28908 33532 28960 33584
rect 28632 33507 28684 33516
rect 28632 33473 28641 33507
rect 28641 33473 28675 33507
rect 28675 33473 28684 33507
rect 28632 33464 28684 33473
rect 31208 33507 31260 33516
rect 8944 33396 8996 33448
rect 12164 33439 12216 33448
rect 12164 33405 12173 33439
rect 12173 33405 12207 33439
rect 12207 33405 12216 33439
rect 12164 33396 12216 33405
rect 24952 33439 25004 33448
rect 24952 33405 24961 33439
rect 24961 33405 24995 33439
rect 24995 33405 25004 33439
rect 24952 33396 25004 33405
rect 28356 33396 28408 33448
rect 31208 33473 31217 33507
rect 31217 33473 31251 33507
rect 31251 33473 31260 33507
rect 31208 33464 31260 33473
rect 35440 33464 35492 33516
rect 31116 33396 31168 33448
rect 39948 33396 40000 33448
rect 48504 33532 48556 33584
rect 52460 33532 52512 33584
rect 41788 33464 41840 33516
rect 42616 33507 42668 33516
rect 42616 33473 42625 33507
rect 42625 33473 42659 33507
rect 42659 33473 42668 33507
rect 42616 33464 42668 33473
rect 43352 33464 43404 33516
rect 44732 33464 44784 33516
rect 44916 33507 44968 33516
rect 44916 33473 44925 33507
rect 44925 33473 44959 33507
rect 44959 33473 44968 33507
rect 44916 33464 44968 33473
rect 45100 33507 45152 33516
rect 45100 33473 45109 33507
rect 45109 33473 45143 33507
rect 45143 33473 45152 33507
rect 45100 33464 45152 33473
rect 45192 33464 45244 33516
rect 48964 33507 49016 33516
rect 48964 33473 48973 33507
rect 48973 33473 49007 33507
rect 49007 33473 49016 33507
rect 48964 33464 49016 33473
rect 49332 33507 49384 33516
rect 45008 33396 45060 33448
rect 49332 33473 49341 33507
rect 49341 33473 49375 33507
rect 49375 33473 49384 33507
rect 49332 33464 49384 33473
rect 51264 33464 51316 33516
rect 52644 33464 52696 33516
rect 58164 33507 58216 33516
rect 58164 33473 58173 33507
rect 58173 33473 58207 33507
rect 58207 33473 58216 33507
rect 58164 33464 58216 33473
rect 7656 33328 7708 33380
rect 8116 33328 8168 33380
rect 26332 33328 26384 33380
rect 1768 33260 1820 33312
rect 32404 33328 32456 33380
rect 45560 33328 45612 33380
rect 53472 33328 53524 33380
rect 27988 33260 28040 33312
rect 28540 33260 28592 33312
rect 30196 33260 30248 33312
rect 35716 33260 35768 33312
rect 35900 33303 35952 33312
rect 35900 33269 35909 33303
rect 35909 33269 35943 33303
rect 35943 33269 35952 33303
rect 35900 33260 35952 33269
rect 52184 33260 52236 33312
rect 52828 33260 52880 33312
rect 4214 33158 4266 33210
rect 4278 33158 4330 33210
rect 4342 33158 4394 33210
rect 4406 33158 4458 33210
rect 4470 33158 4522 33210
rect 34934 33158 34986 33210
rect 34998 33158 35050 33210
rect 35062 33158 35114 33210
rect 35126 33158 35178 33210
rect 35190 33158 35242 33210
rect 1584 33099 1636 33108
rect 1584 33065 1593 33099
rect 1593 33065 1627 33099
rect 1627 33065 1636 33099
rect 1584 33056 1636 33065
rect 8944 33099 8996 33108
rect 8944 33065 8953 33099
rect 8953 33065 8987 33099
rect 8987 33065 8996 33099
rect 8944 33056 8996 33065
rect 18420 33056 18472 33108
rect 27988 33056 28040 33108
rect 28632 33056 28684 33108
rect 48872 33099 48924 33108
rect 48872 33065 48881 33099
rect 48881 33065 48915 33099
rect 48915 33065 48924 33099
rect 48872 33056 48924 33065
rect 58164 33099 58216 33108
rect 58164 33065 58173 33099
rect 58173 33065 58207 33099
rect 58207 33065 58216 33099
rect 58164 33056 58216 33065
rect 17132 32988 17184 33040
rect 19248 33031 19300 33040
rect 19248 32997 19257 33031
rect 19257 32997 19291 33031
rect 19291 32997 19300 33031
rect 19248 32988 19300 32997
rect 7656 32963 7708 32972
rect 7656 32929 7665 32963
rect 7665 32929 7699 32963
rect 7699 32929 7708 32963
rect 7656 32920 7708 32929
rect 18788 32920 18840 32972
rect 23204 32920 23256 32972
rect 26332 32963 26384 32972
rect 26332 32929 26341 32963
rect 26341 32929 26375 32963
rect 26375 32929 26384 32963
rect 38660 32988 38712 33040
rect 28264 32963 28316 32972
rect 26332 32920 26384 32929
rect 7104 32895 7156 32904
rect 7104 32861 7113 32895
rect 7113 32861 7147 32895
rect 7147 32861 7156 32895
rect 7104 32852 7156 32861
rect 7288 32895 7340 32904
rect 7288 32861 7297 32895
rect 7297 32861 7331 32895
rect 7331 32861 7340 32895
rect 7288 32852 7340 32861
rect 8116 32895 8168 32904
rect 8116 32861 8125 32895
rect 8125 32861 8159 32895
rect 8159 32861 8168 32895
rect 8116 32852 8168 32861
rect 11152 32852 11204 32904
rect 11612 32895 11664 32904
rect 11612 32861 11621 32895
rect 11621 32861 11655 32895
rect 11655 32861 11664 32895
rect 11612 32852 11664 32861
rect 11980 32895 12032 32904
rect 11980 32861 11989 32895
rect 11989 32861 12023 32895
rect 12023 32861 12032 32895
rect 11980 32852 12032 32861
rect 12164 32852 12216 32904
rect 16580 32852 16632 32904
rect 10876 32784 10928 32836
rect 17224 32784 17276 32836
rect 7380 32716 7432 32768
rect 8116 32716 8168 32768
rect 13268 32716 13320 32768
rect 13728 32716 13780 32768
rect 18328 32852 18380 32904
rect 18512 32895 18564 32904
rect 18512 32861 18521 32895
rect 18521 32861 18555 32895
rect 18555 32861 18564 32895
rect 18512 32852 18564 32861
rect 19340 32852 19392 32904
rect 22008 32895 22060 32904
rect 18236 32827 18288 32836
rect 18236 32793 18245 32827
rect 18245 32793 18279 32827
rect 18279 32793 18288 32827
rect 18236 32784 18288 32793
rect 17592 32716 17644 32768
rect 22008 32861 22017 32895
rect 22017 32861 22051 32895
rect 22051 32861 22060 32895
rect 22008 32852 22060 32861
rect 22284 32895 22336 32904
rect 22284 32861 22293 32895
rect 22293 32861 22327 32895
rect 22327 32861 22336 32895
rect 22284 32852 22336 32861
rect 28264 32929 28273 32963
rect 28273 32929 28307 32963
rect 28307 32929 28316 32963
rect 28264 32920 28316 32929
rect 30472 32963 30524 32972
rect 30472 32929 30481 32963
rect 30481 32929 30515 32963
rect 30515 32929 30524 32963
rect 30472 32920 30524 32929
rect 31392 32920 31444 32972
rect 35900 32920 35952 32972
rect 49332 32920 49384 32972
rect 27988 32895 28040 32904
rect 27988 32861 27997 32895
rect 27997 32861 28031 32895
rect 28031 32861 28040 32895
rect 27988 32852 28040 32861
rect 30656 32852 30708 32904
rect 34520 32852 34572 32904
rect 35716 32852 35768 32904
rect 37280 32852 37332 32904
rect 27528 32827 27580 32836
rect 24768 32716 24820 32768
rect 26976 32716 27028 32768
rect 27528 32793 27537 32827
rect 27537 32793 27571 32827
rect 27571 32793 27580 32827
rect 27528 32784 27580 32793
rect 38292 32784 38344 32836
rect 44916 32852 44968 32904
rect 45192 32895 45244 32904
rect 45192 32861 45201 32895
rect 45201 32861 45235 32895
rect 45235 32861 45244 32895
rect 45192 32852 45244 32861
rect 45836 32895 45888 32904
rect 45836 32861 45845 32895
rect 45845 32861 45879 32895
rect 45879 32861 45888 32895
rect 45836 32852 45888 32861
rect 46204 32895 46256 32904
rect 46204 32861 46213 32895
rect 46213 32861 46247 32895
rect 46247 32861 46256 32895
rect 46204 32852 46256 32861
rect 48780 32895 48832 32904
rect 48780 32861 48789 32895
rect 48789 32861 48823 32895
rect 48823 32861 48832 32895
rect 48780 32852 48832 32861
rect 48964 32895 49016 32904
rect 48964 32861 48973 32895
rect 48973 32861 49007 32895
rect 49007 32861 49016 32895
rect 48964 32852 49016 32861
rect 47032 32784 47084 32836
rect 52920 32784 52972 32836
rect 27896 32716 27948 32768
rect 33600 32716 33652 32768
rect 35532 32716 35584 32768
rect 39028 32716 39080 32768
rect 45652 32716 45704 32768
rect 19574 32614 19626 32666
rect 19638 32614 19690 32666
rect 19702 32614 19754 32666
rect 19766 32614 19818 32666
rect 19830 32614 19882 32666
rect 50294 32614 50346 32666
rect 50358 32614 50410 32666
rect 50422 32614 50474 32666
rect 50486 32614 50538 32666
rect 50550 32614 50602 32666
rect 2228 32512 2280 32564
rect 33600 32512 33652 32564
rect 8944 32444 8996 32496
rect 9312 32444 9364 32496
rect 15844 32444 15896 32496
rect 7380 32419 7432 32428
rect 7380 32385 7389 32419
rect 7389 32385 7423 32419
rect 7423 32385 7432 32419
rect 7380 32376 7432 32385
rect 8116 32419 8168 32428
rect 8116 32385 8125 32419
rect 8125 32385 8159 32419
rect 8159 32385 8168 32419
rect 8116 32376 8168 32385
rect 10416 32419 10468 32428
rect 10416 32385 10425 32419
rect 10425 32385 10459 32419
rect 10459 32385 10468 32419
rect 10416 32376 10468 32385
rect 13268 32419 13320 32428
rect 13268 32385 13277 32419
rect 13277 32385 13311 32419
rect 13311 32385 13320 32419
rect 13268 32376 13320 32385
rect 13728 32376 13780 32428
rect 15200 32419 15252 32428
rect 15200 32385 15209 32419
rect 15209 32385 15243 32419
rect 15243 32385 15252 32419
rect 15200 32376 15252 32385
rect 10232 32308 10284 32360
rect 10692 32351 10744 32360
rect 10692 32317 10701 32351
rect 10701 32317 10735 32351
rect 10735 32317 10744 32351
rect 10692 32308 10744 32317
rect 15108 32308 15160 32360
rect 15660 32376 15712 32428
rect 18604 32444 18656 32496
rect 24400 32487 24452 32496
rect 24400 32453 24409 32487
rect 24409 32453 24443 32487
rect 24443 32453 24452 32487
rect 24400 32444 24452 32453
rect 24676 32444 24728 32496
rect 24768 32444 24820 32496
rect 18236 32419 18288 32428
rect 18236 32385 18245 32419
rect 18245 32385 18279 32419
rect 18279 32385 18288 32419
rect 18236 32376 18288 32385
rect 18328 32419 18380 32428
rect 18328 32385 18337 32419
rect 18337 32385 18371 32419
rect 18371 32385 18380 32419
rect 18328 32376 18380 32385
rect 18512 32419 18564 32428
rect 18512 32385 18521 32419
rect 18521 32385 18555 32419
rect 18555 32385 18564 32419
rect 24216 32419 24268 32428
rect 18512 32376 18564 32385
rect 24216 32385 24225 32419
rect 24225 32385 24259 32419
rect 24259 32385 24268 32419
rect 24216 32376 24268 32385
rect 22008 32351 22060 32360
rect 22008 32317 22017 32351
rect 22017 32317 22051 32351
rect 22051 32317 22060 32351
rect 22008 32308 22060 32317
rect 22468 32351 22520 32360
rect 22468 32317 22477 32351
rect 22477 32317 22511 32351
rect 22511 32317 22520 32351
rect 22468 32308 22520 32317
rect 8392 32240 8444 32292
rect 15292 32240 15344 32292
rect 16212 32240 16264 32292
rect 22100 32240 22152 32292
rect 22284 32283 22336 32292
rect 22284 32249 22293 32283
rect 22293 32249 22327 32283
rect 22327 32249 22336 32283
rect 22284 32240 22336 32249
rect 31208 32444 31260 32496
rect 37464 32512 37516 32564
rect 38292 32555 38344 32564
rect 38292 32521 38301 32555
rect 38301 32521 38335 32555
rect 38335 32521 38344 32555
rect 38292 32512 38344 32521
rect 40040 32555 40092 32564
rect 40040 32521 40049 32555
rect 40049 32521 40083 32555
rect 40083 32521 40092 32555
rect 40040 32512 40092 32521
rect 46204 32512 46256 32564
rect 48964 32512 49016 32564
rect 30472 32419 30524 32428
rect 30472 32385 30481 32419
rect 30481 32385 30515 32419
rect 30515 32385 30524 32419
rect 30472 32376 30524 32385
rect 30656 32419 30708 32428
rect 30656 32385 30665 32419
rect 30665 32385 30699 32419
rect 30699 32385 30708 32419
rect 30656 32376 30708 32385
rect 35716 32444 35768 32496
rect 33784 32419 33836 32428
rect 33784 32385 33793 32419
rect 33793 32385 33827 32419
rect 33827 32385 33836 32419
rect 33784 32376 33836 32385
rect 33968 32419 34020 32428
rect 33968 32385 33977 32419
rect 33977 32385 34011 32419
rect 34011 32385 34020 32419
rect 33968 32376 34020 32385
rect 34520 32419 34572 32428
rect 34520 32385 34529 32419
rect 34529 32385 34563 32419
rect 34563 32385 34572 32419
rect 34520 32376 34572 32385
rect 34152 32308 34204 32360
rect 56692 32444 56744 32496
rect 37280 32419 37332 32428
rect 37280 32385 37289 32419
rect 37289 32385 37323 32419
rect 37323 32385 37332 32419
rect 37280 32376 37332 32385
rect 38200 32419 38252 32428
rect 38200 32385 38209 32419
rect 38209 32385 38243 32419
rect 38243 32385 38252 32419
rect 38200 32376 38252 32385
rect 39028 32419 39080 32428
rect 37464 32351 37516 32360
rect 37464 32317 37473 32351
rect 37473 32317 37507 32351
rect 37507 32317 37516 32351
rect 37464 32308 37516 32317
rect 10508 32215 10560 32224
rect 10508 32181 10517 32215
rect 10517 32181 10551 32215
rect 10551 32181 10560 32215
rect 10508 32172 10560 32181
rect 14280 32172 14332 32224
rect 14464 32172 14516 32224
rect 16488 32172 16540 32224
rect 17132 32172 17184 32224
rect 21180 32172 21232 32224
rect 27896 32172 27948 32224
rect 38016 32240 38068 32292
rect 39028 32385 39037 32419
rect 39037 32385 39071 32419
rect 39071 32385 39080 32419
rect 39028 32376 39080 32385
rect 39212 32419 39264 32428
rect 39212 32385 39221 32419
rect 39221 32385 39255 32419
rect 39255 32385 39264 32419
rect 39212 32376 39264 32385
rect 41328 32419 41380 32428
rect 41328 32385 41337 32419
rect 41337 32385 41371 32419
rect 41371 32385 41380 32419
rect 41328 32376 41380 32385
rect 43352 32419 43404 32428
rect 43352 32385 43361 32419
rect 43361 32385 43395 32419
rect 43395 32385 43404 32419
rect 43352 32376 43404 32385
rect 44916 32376 44968 32428
rect 45652 32419 45704 32428
rect 45652 32385 45661 32419
rect 45661 32385 45695 32419
rect 45695 32385 45704 32419
rect 45652 32376 45704 32385
rect 47952 32376 48004 32428
rect 49792 32376 49844 32428
rect 52920 32419 52972 32428
rect 52920 32385 52929 32419
rect 52929 32385 52963 32419
rect 52963 32385 52972 32419
rect 52920 32376 52972 32385
rect 41236 32351 41288 32360
rect 41236 32317 41245 32351
rect 41245 32317 41279 32351
rect 41279 32317 41288 32351
rect 41236 32308 41288 32317
rect 41788 32308 41840 32360
rect 45100 32351 45152 32360
rect 45100 32317 45109 32351
rect 45109 32317 45143 32351
rect 45143 32317 45152 32351
rect 45100 32308 45152 32317
rect 53288 32308 53340 32360
rect 45192 32172 45244 32224
rect 52736 32215 52788 32224
rect 52736 32181 52745 32215
rect 52745 32181 52779 32215
rect 52779 32181 52788 32215
rect 52736 32172 52788 32181
rect 4214 32070 4266 32122
rect 4278 32070 4330 32122
rect 4342 32070 4394 32122
rect 4406 32070 4458 32122
rect 4470 32070 4522 32122
rect 34934 32070 34986 32122
rect 34998 32070 35050 32122
rect 35062 32070 35114 32122
rect 35126 32070 35178 32122
rect 35190 32070 35242 32122
rect 1676 31968 1728 32020
rect 8392 32011 8444 32020
rect 8392 31977 8401 32011
rect 8401 31977 8435 32011
rect 8435 31977 8444 32011
rect 8392 31968 8444 31977
rect 8760 31968 8812 32020
rect 9312 32011 9364 32020
rect 9312 31977 9321 32011
rect 9321 31977 9355 32011
rect 9355 31977 9364 32011
rect 9312 31968 9364 31977
rect 10048 31968 10100 32020
rect 10416 31968 10468 32020
rect 15200 31968 15252 32020
rect 15660 32011 15712 32020
rect 15660 31977 15669 32011
rect 15669 31977 15703 32011
rect 15703 31977 15712 32011
rect 15660 31968 15712 31977
rect 16488 32011 16540 32020
rect 9772 31832 9824 31884
rect 9956 31832 10008 31884
rect 10692 31875 10744 31884
rect 10692 31841 10701 31875
rect 10701 31841 10735 31875
rect 10735 31841 10744 31875
rect 10692 31832 10744 31841
rect 14188 31900 14240 31952
rect 14280 31900 14332 31952
rect 16488 31977 16497 32011
rect 16497 31977 16531 32011
rect 16531 31977 16540 32011
rect 16488 31968 16540 31977
rect 16580 31968 16632 32020
rect 17040 32011 17092 32020
rect 17040 31977 17049 32011
rect 17049 31977 17083 32011
rect 17083 31977 17092 32011
rect 17040 31968 17092 31977
rect 18236 31968 18288 32020
rect 1952 31764 2004 31816
rect 3240 31764 3292 31816
rect 1584 31696 1636 31748
rect 7196 31764 7248 31816
rect 8208 31764 8260 31816
rect 10048 31807 10100 31816
rect 10048 31773 10057 31807
rect 10057 31773 10091 31807
rect 10091 31773 10100 31807
rect 10048 31764 10100 31773
rect 10140 31807 10192 31816
rect 10140 31773 10149 31807
rect 10149 31773 10183 31807
rect 10183 31773 10192 31807
rect 10140 31764 10192 31773
rect 10508 31764 10560 31816
rect 13544 31807 13596 31816
rect 13544 31773 13553 31807
rect 13553 31773 13587 31807
rect 13587 31773 13596 31807
rect 13544 31764 13596 31773
rect 7288 31696 7340 31748
rect 13360 31696 13412 31748
rect 17224 31900 17276 31952
rect 27068 31968 27120 32020
rect 27528 31968 27580 32020
rect 33968 31968 34020 32020
rect 34152 32011 34204 32020
rect 34152 31977 34161 32011
rect 34161 31977 34195 32011
rect 34195 31977 34204 32011
rect 34152 31968 34204 31977
rect 43352 31968 43404 32020
rect 45008 31968 45060 32020
rect 47952 32011 48004 32020
rect 47952 31977 47961 32011
rect 47961 31977 47995 32011
rect 47995 31977 48004 32011
rect 47952 31968 48004 31977
rect 49056 32011 49108 32020
rect 49056 31977 49065 32011
rect 49065 31977 49099 32011
rect 49099 31977 49108 32011
rect 49056 31968 49108 31977
rect 53288 31968 53340 32020
rect 16212 31764 16264 31816
rect 17960 31807 18012 31816
rect 17960 31773 17969 31807
rect 17969 31773 18003 31807
rect 18003 31773 18012 31807
rect 17960 31764 18012 31773
rect 18052 31764 18104 31816
rect 30472 31900 30524 31952
rect 32128 31900 32180 31952
rect 20996 31832 21048 31884
rect 22008 31832 22060 31884
rect 24216 31832 24268 31884
rect 26884 31832 26936 31884
rect 28632 31832 28684 31884
rect 30656 31875 30708 31884
rect 30656 31841 30665 31875
rect 30665 31841 30699 31875
rect 30699 31841 30708 31875
rect 30656 31832 30708 31841
rect 35716 31875 35768 31884
rect 24400 31764 24452 31816
rect 26976 31807 27028 31816
rect 26976 31773 26985 31807
rect 26985 31773 27019 31807
rect 27019 31773 27028 31807
rect 26976 31764 27028 31773
rect 27804 31764 27856 31816
rect 28356 31696 28408 31748
rect 29736 31764 29788 31816
rect 33968 31807 34020 31816
rect 33968 31773 33977 31807
rect 33977 31773 34011 31807
rect 34011 31773 34020 31807
rect 33968 31764 34020 31773
rect 34152 31807 34204 31816
rect 34152 31773 34161 31807
rect 34161 31773 34195 31807
rect 34195 31773 34204 31807
rect 34152 31764 34204 31773
rect 32220 31696 32272 31748
rect 35716 31841 35725 31875
rect 35725 31841 35759 31875
rect 35759 31841 35768 31875
rect 35716 31832 35768 31841
rect 38660 31875 38712 31884
rect 38660 31841 38669 31875
rect 38669 31841 38703 31875
rect 38703 31841 38712 31875
rect 38660 31832 38712 31841
rect 38016 31807 38068 31816
rect 38016 31773 38025 31807
rect 38025 31773 38059 31807
rect 38059 31773 38068 31807
rect 38016 31764 38068 31773
rect 38200 31807 38252 31816
rect 38200 31773 38209 31807
rect 38209 31773 38243 31807
rect 38243 31773 38252 31807
rect 38200 31764 38252 31773
rect 39028 31900 39080 31952
rect 41052 31900 41104 31952
rect 41236 31832 41288 31884
rect 41328 31832 41380 31884
rect 39212 31764 39264 31816
rect 45652 31832 45704 31884
rect 45100 31807 45152 31816
rect 45100 31773 45109 31807
rect 45109 31773 45143 31807
rect 45143 31773 45152 31807
rect 45100 31764 45152 31773
rect 45560 31807 45612 31816
rect 45560 31773 45569 31807
rect 45569 31773 45603 31807
rect 45603 31773 45612 31807
rect 48228 31832 48280 31884
rect 48412 31832 48464 31884
rect 45560 31764 45612 31773
rect 48688 31807 48740 31816
rect 45376 31739 45428 31748
rect 45376 31705 45385 31739
rect 45385 31705 45419 31739
rect 45419 31705 45428 31739
rect 48688 31773 48697 31807
rect 48697 31773 48731 31807
rect 48731 31773 48740 31807
rect 48688 31764 48740 31773
rect 52920 31807 52972 31816
rect 52920 31773 52929 31807
rect 52929 31773 52963 31807
rect 52963 31773 52972 31807
rect 52920 31764 52972 31773
rect 53288 31807 53340 31816
rect 53288 31773 53297 31807
rect 53297 31773 53331 31807
rect 53331 31773 53340 31807
rect 53288 31764 53340 31773
rect 45376 31696 45428 31705
rect 48596 31696 48648 31748
rect 52276 31696 52328 31748
rect 55496 31764 55548 31816
rect 56324 31807 56376 31816
rect 56324 31773 56333 31807
rect 56333 31773 56367 31807
rect 56367 31773 56376 31807
rect 56324 31764 56376 31773
rect 57888 31764 57940 31816
rect 8944 31671 8996 31680
rect 8944 31637 8953 31671
rect 8953 31637 8987 31671
rect 8987 31637 8996 31671
rect 8944 31628 8996 31637
rect 13176 31628 13228 31680
rect 18236 31628 18288 31680
rect 29092 31628 29144 31680
rect 19574 31526 19626 31578
rect 19638 31526 19690 31578
rect 19702 31526 19754 31578
rect 19766 31526 19818 31578
rect 19830 31526 19882 31578
rect 50294 31526 50346 31578
rect 50358 31526 50410 31578
rect 50422 31526 50474 31578
rect 50486 31526 50538 31578
rect 50550 31526 50602 31578
rect 10048 31467 10100 31476
rect 10048 31433 10057 31467
rect 10057 31433 10091 31467
rect 10091 31433 10100 31467
rect 10048 31424 10100 31433
rect 15108 31424 15160 31476
rect 1584 31399 1636 31408
rect 1584 31365 1593 31399
rect 1593 31365 1627 31399
rect 1627 31365 1636 31399
rect 1584 31356 1636 31365
rect 7104 31356 7156 31408
rect 8944 31356 8996 31408
rect 13360 31399 13412 31408
rect 13360 31365 13369 31399
rect 13369 31365 13403 31399
rect 13403 31365 13412 31399
rect 13360 31356 13412 31365
rect 13544 31399 13596 31408
rect 13544 31365 13569 31399
rect 13569 31365 13596 31399
rect 13544 31356 13596 31365
rect 17960 31356 18012 31408
rect 19524 31356 19576 31408
rect 22836 31399 22888 31408
rect 7196 31331 7248 31340
rect 7196 31297 7205 31331
rect 7205 31297 7239 31331
rect 7239 31297 7248 31331
rect 7196 31288 7248 31297
rect 8116 31288 8168 31340
rect 10048 31288 10100 31340
rect 18052 31331 18104 31340
rect 18052 31297 18061 31331
rect 18061 31297 18095 31331
rect 18095 31297 18104 31331
rect 18052 31288 18104 31297
rect 18236 31331 18288 31340
rect 18236 31297 18245 31331
rect 18245 31297 18279 31331
rect 18279 31297 18288 31331
rect 18236 31288 18288 31297
rect 18512 31331 18564 31340
rect 18512 31297 18521 31331
rect 18521 31297 18555 31331
rect 18555 31297 18564 31331
rect 18512 31288 18564 31297
rect 9496 31220 9548 31272
rect 10600 31220 10652 31272
rect 18328 31220 18380 31272
rect 22836 31365 22845 31399
rect 22845 31365 22879 31399
rect 22879 31365 22888 31399
rect 22836 31356 22888 31365
rect 27068 31399 27120 31408
rect 27068 31365 27077 31399
rect 27077 31365 27111 31399
rect 27111 31365 27120 31399
rect 27068 31356 27120 31365
rect 27804 31356 27856 31408
rect 7564 31152 7616 31204
rect 22284 31152 22336 31204
rect 9864 31127 9916 31136
rect 9864 31093 9873 31127
rect 9873 31093 9907 31127
rect 9907 31093 9916 31127
rect 9864 31084 9916 31093
rect 10324 31084 10376 31136
rect 13176 31084 13228 31136
rect 18328 31084 18380 31136
rect 26700 31220 26752 31272
rect 28632 31331 28684 31340
rect 28632 31297 28641 31331
rect 28641 31297 28675 31331
rect 28675 31297 28684 31331
rect 28632 31288 28684 31297
rect 33784 31424 33836 31476
rect 38200 31424 38252 31476
rect 48596 31424 48648 31476
rect 48688 31424 48740 31476
rect 49792 31467 49844 31476
rect 49792 31433 49801 31467
rect 49801 31433 49835 31467
rect 49835 31433 49844 31467
rect 49792 31424 49844 31433
rect 32128 31399 32180 31408
rect 32128 31365 32137 31399
rect 32137 31365 32171 31399
rect 32171 31365 32180 31399
rect 32128 31356 32180 31365
rect 29736 31288 29788 31340
rect 33968 31288 34020 31340
rect 37556 31288 37608 31340
rect 40500 31288 40552 31340
rect 45376 31288 45428 31340
rect 45652 31288 45704 31340
rect 48320 31288 48372 31340
rect 52736 31356 52788 31408
rect 54944 31399 54996 31408
rect 54944 31365 54953 31399
rect 54953 31365 54987 31399
rect 54987 31365 54996 31399
rect 54944 31356 54996 31365
rect 37372 31263 37424 31272
rect 37372 31229 37381 31263
rect 37381 31229 37415 31263
rect 37415 31229 37424 31263
rect 37372 31220 37424 31229
rect 40684 31263 40736 31272
rect 40684 31229 40693 31263
rect 40693 31229 40727 31263
rect 40727 31229 40736 31263
rect 40684 31220 40736 31229
rect 41328 31220 41380 31272
rect 45100 31220 45152 31272
rect 45284 31220 45336 31272
rect 48228 31220 48280 31272
rect 48780 31220 48832 31272
rect 52368 31288 52420 31340
rect 55404 31331 55456 31340
rect 55404 31297 55413 31331
rect 55413 31297 55447 31331
rect 55447 31297 55456 31331
rect 55404 31288 55456 31297
rect 52276 31220 52328 31272
rect 55312 31220 55364 31272
rect 32220 31152 32272 31204
rect 44824 31195 44876 31204
rect 44824 31161 44833 31195
rect 44833 31161 44867 31195
rect 44867 31161 44876 31195
rect 44824 31152 44876 31161
rect 45652 31195 45704 31204
rect 45652 31161 45661 31195
rect 45661 31161 45695 31195
rect 45695 31161 45704 31195
rect 45652 31152 45704 31161
rect 49976 31152 50028 31204
rect 50068 31152 50120 31204
rect 52368 31152 52420 31204
rect 28356 31127 28408 31136
rect 28356 31093 28365 31127
rect 28365 31093 28399 31127
rect 28399 31093 28408 31127
rect 28356 31084 28408 31093
rect 29092 31127 29144 31136
rect 29092 31093 29101 31127
rect 29101 31093 29135 31127
rect 29135 31093 29144 31127
rect 29092 31084 29144 31093
rect 48320 31084 48372 31136
rect 52000 31084 52052 31136
rect 4214 30982 4266 31034
rect 4278 30982 4330 31034
rect 4342 30982 4394 31034
rect 4406 30982 4458 31034
rect 4470 30982 4522 31034
rect 34934 30982 34986 31034
rect 34998 30982 35050 31034
rect 35062 30982 35114 31034
rect 35126 30982 35178 31034
rect 35190 30982 35242 31034
rect 10140 30880 10192 30932
rect 12900 30880 12952 30932
rect 19340 30923 19392 30932
rect 19340 30889 19349 30923
rect 19349 30889 19383 30923
rect 19383 30889 19392 30923
rect 19340 30880 19392 30889
rect 22100 30880 22152 30932
rect 27804 30923 27856 30932
rect 27804 30889 27813 30923
rect 27813 30889 27847 30923
rect 27847 30889 27856 30923
rect 27804 30880 27856 30889
rect 37372 30923 37424 30932
rect 37372 30889 37381 30923
rect 37381 30889 37415 30923
rect 37415 30889 37424 30923
rect 37372 30880 37424 30889
rect 45192 30880 45244 30932
rect 45284 30880 45336 30932
rect 55496 30923 55548 30932
rect 55496 30889 55505 30923
rect 55505 30889 55539 30923
rect 55539 30889 55548 30923
rect 55496 30880 55548 30889
rect 10324 30855 10376 30864
rect 10324 30821 10333 30855
rect 10333 30821 10367 30855
rect 10367 30821 10376 30855
rect 10324 30812 10376 30821
rect 13360 30812 13412 30864
rect 7288 30719 7340 30728
rect 7288 30685 7297 30719
rect 7297 30685 7331 30719
rect 7331 30685 7340 30719
rect 7288 30676 7340 30685
rect 9864 30676 9916 30728
rect 10600 30744 10652 30796
rect 12716 30744 12768 30796
rect 13268 30744 13320 30796
rect 12992 30719 13044 30728
rect 10048 30540 10100 30592
rect 12992 30685 13001 30719
rect 13001 30685 13035 30719
rect 13035 30685 13044 30719
rect 12992 30676 13044 30685
rect 13084 30719 13136 30728
rect 13084 30685 13093 30719
rect 13093 30685 13127 30719
rect 13127 30685 13136 30719
rect 16948 30812 17000 30864
rect 18052 30855 18104 30864
rect 18052 30821 18061 30855
rect 18061 30821 18095 30855
rect 18095 30821 18104 30855
rect 18052 30812 18104 30821
rect 22836 30812 22888 30864
rect 18328 30787 18380 30796
rect 18328 30753 18337 30787
rect 18337 30753 18371 30787
rect 18371 30753 18380 30787
rect 18328 30744 18380 30753
rect 26884 30787 26936 30796
rect 26884 30753 26893 30787
rect 26893 30753 26927 30787
rect 26927 30753 26936 30787
rect 30472 30787 30524 30796
rect 26884 30744 26936 30753
rect 14372 30719 14424 30728
rect 13084 30676 13136 30685
rect 14372 30685 14381 30719
rect 14381 30685 14415 30719
rect 14415 30685 14424 30719
rect 14372 30676 14424 30685
rect 14556 30719 14608 30728
rect 14556 30685 14565 30719
rect 14565 30685 14599 30719
rect 14599 30685 14608 30719
rect 14556 30676 14608 30685
rect 15844 30676 15896 30728
rect 11244 30608 11296 30660
rect 19340 30676 19392 30728
rect 19432 30676 19484 30728
rect 22836 30719 22888 30728
rect 19524 30608 19576 30660
rect 22836 30685 22845 30719
rect 22845 30685 22879 30719
rect 22879 30685 22888 30719
rect 22836 30676 22888 30685
rect 23112 30719 23164 30728
rect 23112 30685 23121 30719
rect 23121 30685 23155 30719
rect 23155 30685 23164 30719
rect 23112 30676 23164 30685
rect 26976 30719 27028 30728
rect 26976 30685 26985 30719
rect 26985 30685 27019 30719
rect 27019 30685 27028 30719
rect 26976 30676 27028 30685
rect 30472 30753 30481 30787
rect 30481 30753 30515 30787
rect 30515 30753 30524 30787
rect 30472 30744 30524 30753
rect 32128 30812 32180 30864
rect 51356 30812 51408 30864
rect 28724 30676 28776 30728
rect 45008 30787 45060 30796
rect 45008 30753 45017 30787
rect 45017 30753 45051 30787
rect 45051 30753 45060 30787
rect 45008 30744 45060 30753
rect 55312 30787 55364 30796
rect 55312 30753 55321 30787
rect 55321 30753 55355 30787
rect 55355 30753 55364 30787
rect 55312 30744 55364 30753
rect 34520 30676 34572 30728
rect 37188 30719 37240 30728
rect 37188 30685 37197 30719
rect 37197 30685 37231 30719
rect 37231 30685 37240 30719
rect 37188 30676 37240 30685
rect 37464 30676 37516 30728
rect 44364 30676 44416 30728
rect 45376 30676 45428 30728
rect 48320 30719 48372 30728
rect 48320 30685 48329 30719
rect 48329 30685 48363 30719
rect 48363 30685 48372 30719
rect 48320 30676 48372 30685
rect 48412 30719 48464 30728
rect 48412 30685 48421 30719
rect 48421 30685 48455 30719
rect 48455 30685 48464 30719
rect 48412 30676 48464 30685
rect 48596 30719 48648 30728
rect 48596 30685 48605 30719
rect 48605 30685 48639 30719
rect 48639 30685 48648 30719
rect 48780 30719 48832 30728
rect 48596 30676 48648 30685
rect 48780 30685 48789 30719
rect 48789 30685 48823 30719
rect 48823 30685 48832 30719
rect 48780 30676 48832 30685
rect 49976 30676 50028 30728
rect 50896 30719 50948 30728
rect 50896 30685 50905 30719
rect 50905 30685 50939 30719
rect 50939 30685 50948 30719
rect 50896 30676 50948 30685
rect 52276 30719 52328 30728
rect 52276 30685 52285 30719
rect 52285 30685 52319 30719
rect 52319 30685 52328 30719
rect 52276 30676 52328 30685
rect 52368 30676 52420 30728
rect 55772 30719 55824 30728
rect 55772 30685 55781 30719
rect 55781 30685 55815 30719
rect 55815 30685 55824 30719
rect 55772 30676 55824 30685
rect 29092 30608 29144 30660
rect 44824 30608 44876 30660
rect 48228 30608 48280 30660
rect 51080 30651 51132 30660
rect 51080 30617 51089 30651
rect 51089 30617 51123 30651
rect 51123 30617 51132 30651
rect 51080 30608 51132 30617
rect 52184 30608 52236 30660
rect 12716 30540 12768 30592
rect 13084 30540 13136 30592
rect 13544 30540 13596 30592
rect 17500 30540 17552 30592
rect 19432 30540 19484 30592
rect 19984 30540 20036 30592
rect 22192 30583 22244 30592
rect 22192 30549 22201 30583
rect 22201 30549 22235 30583
rect 22235 30549 22244 30583
rect 23020 30583 23072 30592
rect 22192 30540 22244 30549
rect 23020 30549 23029 30583
rect 23029 30549 23063 30583
rect 23063 30549 23072 30583
rect 23020 30540 23072 30549
rect 24768 30540 24820 30592
rect 27712 30540 27764 30592
rect 28724 30583 28776 30592
rect 28724 30549 28733 30583
rect 28733 30549 28767 30583
rect 28767 30549 28776 30583
rect 28724 30540 28776 30549
rect 45468 30583 45520 30592
rect 45468 30549 45477 30583
rect 45477 30549 45511 30583
rect 45511 30549 45520 30583
rect 45468 30540 45520 30549
rect 51632 30540 51684 30592
rect 56048 30540 56100 30592
rect 19574 30438 19626 30490
rect 19638 30438 19690 30490
rect 19702 30438 19754 30490
rect 19766 30438 19818 30490
rect 19830 30438 19882 30490
rect 50294 30438 50346 30490
rect 50358 30438 50410 30490
rect 50422 30438 50474 30490
rect 50486 30438 50538 30490
rect 50550 30438 50602 30490
rect 10324 30336 10376 30388
rect 10784 30336 10836 30388
rect 10968 30336 11020 30388
rect 9496 30268 9548 30320
rect 10048 30268 10100 30320
rect 13176 30311 13228 30320
rect 13176 30277 13185 30311
rect 13185 30277 13219 30311
rect 13219 30277 13228 30311
rect 13176 30268 13228 30277
rect 16028 30268 16080 30320
rect 5448 30200 5500 30252
rect 6920 30200 6972 30252
rect 7656 30243 7708 30252
rect 7656 30209 7665 30243
rect 7665 30209 7699 30243
rect 7699 30209 7708 30243
rect 7656 30200 7708 30209
rect 10692 30200 10744 30252
rect 12900 30243 12952 30252
rect 12900 30209 12909 30243
rect 12909 30209 12943 30243
rect 12943 30209 12952 30243
rect 12900 30200 12952 30209
rect 12992 30243 13044 30252
rect 12992 30209 13001 30243
rect 13001 30209 13035 30243
rect 13035 30209 13044 30243
rect 12992 30200 13044 30209
rect 9128 30132 9180 30184
rect 12440 30132 12492 30184
rect 13268 30132 13320 30184
rect 14556 30132 14608 30184
rect 13820 30064 13872 30116
rect 15568 30243 15620 30252
rect 15568 30209 15577 30243
rect 15577 30209 15611 30243
rect 15611 30209 15620 30243
rect 15844 30243 15896 30252
rect 15568 30200 15620 30209
rect 15844 30209 15853 30243
rect 15853 30209 15887 30243
rect 15887 30209 15896 30243
rect 15844 30200 15896 30209
rect 15936 30200 15988 30252
rect 16948 30243 17000 30252
rect 16948 30209 16957 30243
rect 16957 30209 16991 30243
rect 16991 30209 17000 30243
rect 16948 30200 17000 30209
rect 17868 30200 17920 30252
rect 19984 30268 20036 30320
rect 22836 30336 22888 30388
rect 24400 30336 24452 30388
rect 26976 30336 27028 30388
rect 28724 30336 28776 30388
rect 40408 30336 40460 30388
rect 40684 30336 40736 30388
rect 44364 30379 44416 30388
rect 44364 30345 44373 30379
rect 44373 30345 44407 30379
rect 44407 30345 44416 30379
rect 44364 30336 44416 30345
rect 44824 30336 44876 30388
rect 48780 30336 48832 30388
rect 55312 30336 55364 30388
rect 55404 30336 55456 30388
rect 19800 30175 19852 30184
rect 18236 30064 18288 30116
rect 19800 30141 19809 30175
rect 19809 30141 19843 30175
rect 19843 30141 19852 30175
rect 19800 30132 19852 30141
rect 22928 30200 22980 30252
rect 23112 30200 23164 30252
rect 30380 30268 30432 30320
rect 34152 30268 34204 30320
rect 37188 30268 37240 30320
rect 24860 30200 24912 30252
rect 32680 30200 32732 30252
rect 34428 30200 34480 30252
rect 24308 30132 24360 30184
rect 32772 30175 32824 30184
rect 32772 30141 32781 30175
rect 32781 30141 32815 30175
rect 32815 30141 32824 30175
rect 32772 30132 32824 30141
rect 32956 30132 33008 30184
rect 37464 30200 37516 30252
rect 40500 30268 40552 30320
rect 43076 30268 43128 30320
rect 42432 30243 42484 30252
rect 39672 30175 39724 30184
rect 39672 30141 39681 30175
rect 39681 30141 39715 30175
rect 39715 30141 39724 30175
rect 39672 30132 39724 30141
rect 20996 30064 21048 30116
rect 27068 30064 27120 30116
rect 30932 30064 30984 30116
rect 37556 30064 37608 30116
rect 42432 30209 42441 30243
rect 42441 30209 42475 30243
rect 42475 30209 42484 30243
rect 42432 30200 42484 30209
rect 44272 30243 44324 30252
rect 39856 30132 39908 30184
rect 42524 30132 42576 30184
rect 44272 30209 44281 30243
rect 44281 30209 44315 30243
rect 44315 30209 44324 30243
rect 44272 30200 44324 30209
rect 45008 30200 45060 30252
rect 45100 30200 45152 30252
rect 48044 30200 48096 30252
rect 51632 30243 51684 30252
rect 49516 30064 49568 30116
rect 51632 30209 51641 30243
rect 51641 30209 51675 30243
rect 51675 30209 51684 30243
rect 51632 30200 51684 30209
rect 55312 30243 55364 30252
rect 55312 30209 55321 30243
rect 55321 30209 55355 30243
rect 55355 30209 55364 30243
rect 55312 30200 55364 30209
rect 55680 30200 55732 30252
rect 52092 30175 52144 30184
rect 52092 30141 52101 30175
rect 52101 30141 52135 30175
rect 52135 30141 52144 30175
rect 52092 30132 52144 30141
rect 51724 30064 51776 30116
rect 10508 29996 10560 30048
rect 11060 29996 11112 30048
rect 15384 29996 15436 30048
rect 18420 29996 18472 30048
rect 22192 29996 22244 30048
rect 22928 29996 22980 30048
rect 24768 29996 24820 30048
rect 34428 29996 34480 30048
rect 40592 30039 40644 30048
rect 40592 30005 40601 30039
rect 40601 30005 40635 30039
rect 40635 30005 40644 30039
rect 40592 29996 40644 30005
rect 45192 29996 45244 30048
rect 45376 29996 45428 30048
rect 48504 29996 48556 30048
rect 53012 29996 53064 30048
rect 56048 29996 56100 30048
rect 4214 29894 4266 29946
rect 4278 29894 4330 29946
rect 4342 29894 4394 29946
rect 4406 29894 4458 29946
rect 4470 29894 4522 29946
rect 34934 29894 34986 29946
rect 34998 29894 35050 29946
rect 35062 29894 35114 29946
rect 35126 29894 35178 29946
rect 35190 29894 35242 29946
rect 2228 29835 2280 29844
rect 2228 29801 2237 29835
rect 2237 29801 2271 29835
rect 2271 29801 2280 29835
rect 2228 29792 2280 29801
rect 7380 29792 7432 29844
rect 9680 29835 9732 29844
rect 9680 29801 9689 29835
rect 9689 29801 9723 29835
rect 9723 29801 9732 29835
rect 9680 29792 9732 29801
rect 9864 29835 9916 29844
rect 9864 29801 9873 29835
rect 9873 29801 9907 29835
rect 9907 29801 9916 29835
rect 9864 29792 9916 29801
rect 10692 29835 10744 29844
rect 10692 29801 10701 29835
rect 10701 29801 10735 29835
rect 10735 29801 10744 29835
rect 10692 29792 10744 29801
rect 10784 29792 10836 29844
rect 12992 29835 13044 29844
rect 12992 29801 13001 29835
rect 13001 29801 13035 29835
rect 13035 29801 13044 29835
rect 12992 29792 13044 29801
rect 14464 29835 14516 29844
rect 14464 29801 14473 29835
rect 14473 29801 14507 29835
rect 14507 29801 14516 29835
rect 14464 29792 14516 29801
rect 15108 29792 15160 29844
rect 15384 29835 15436 29844
rect 15384 29801 15393 29835
rect 15393 29801 15427 29835
rect 15427 29801 15436 29835
rect 15384 29792 15436 29801
rect 15844 29835 15896 29844
rect 15844 29801 15853 29835
rect 15853 29801 15887 29835
rect 15887 29801 15896 29835
rect 15844 29792 15896 29801
rect 19984 29792 20036 29844
rect 22928 29835 22980 29844
rect 22928 29801 22937 29835
rect 22937 29801 22971 29835
rect 22971 29801 22980 29835
rect 22928 29792 22980 29801
rect 23020 29792 23072 29844
rect 11060 29724 11112 29776
rect 19064 29724 19116 29776
rect 19156 29724 19208 29776
rect 3332 29656 3384 29708
rect 5724 29699 5776 29708
rect 5724 29665 5733 29699
rect 5733 29665 5767 29699
rect 5767 29665 5776 29699
rect 5724 29656 5776 29665
rect 7656 29699 7708 29708
rect 7656 29665 7665 29699
rect 7665 29665 7699 29699
rect 7699 29665 7708 29699
rect 7656 29656 7708 29665
rect 19432 29656 19484 29708
rect 2228 29588 2280 29640
rect 5448 29588 5500 29640
rect 7380 29631 7432 29640
rect 7380 29597 7389 29631
rect 7389 29597 7423 29631
rect 7423 29597 7432 29631
rect 7380 29588 7432 29597
rect 9680 29588 9732 29640
rect 12440 29631 12492 29640
rect 12440 29597 12449 29631
rect 12449 29597 12483 29631
rect 12483 29597 12492 29631
rect 12440 29588 12492 29597
rect 13636 29588 13688 29640
rect 15016 29631 15068 29640
rect 15016 29597 15025 29631
rect 15025 29597 15059 29631
rect 15059 29597 15068 29631
rect 15016 29588 15068 29597
rect 15108 29588 15160 29640
rect 16028 29631 16080 29640
rect 16028 29597 16037 29631
rect 16037 29597 16071 29631
rect 16071 29597 16080 29631
rect 16028 29588 16080 29597
rect 16212 29631 16264 29640
rect 16212 29597 16221 29631
rect 16221 29597 16255 29631
rect 16255 29597 16264 29631
rect 16212 29588 16264 29597
rect 17868 29588 17920 29640
rect 7472 29520 7524 29572
rect 12624 29563 12676 29572
rect 12624 29529 12633 29563
rect 12633 29529 12667 29563
rect 12667 29529 12676 29563
rect 12624 29520 12676 29529
rect 1492 29495 1544 29504
rect 1492 29461 1501 29495
rect 1501 29461 1535 29495
rect 1535 29461 1544 29495
rect 1492 29452 1544 29461
rect 4344 29495 4396 29504
rect 4344 29461 4353 29495
rect 4353 29461 4387 29495
rect 4387 29461 4396 29495
rect 4344 29452 4396 29461
rect 4896 29495 4948 29504
rect 4896 29461 4905 29495
rect 4905 29461 4939 29495
rect 4939 29461 4948 29495
rect 4896 29452 4948 29461
rect 9864 29452 9916 29504
rect 12256 29452 12308 29504
rect 12348 29452 12400 29504
rect 14188 29520 14240 29572
rect 19800 29520 19852 29572
rect 23112 29656 23164 29708
rect 24860 29724 24912 29776
rect 25412 29724 25464 29776
rect 27804 29792 27856 29844
rect 28356 29792 28408 29844
rect 30380 29792 30432 29844
rect 32956 29835 33008 29844
rect 32956 29801 32965 29835
rect 32965 29801 32999 29835
rect 32999 29801 33008 29835
rect 32956 29792 33008 29801
rect 37188 29792 37240 29844
rect 37464 29835 37516 29844
rect 37464 29801 37473 29835
rect 37473 29801 37507 29835
rect 37507 29801 37516 29835
rect 37464 29792 37516 29801
rect 42524 29792 42576 29844
rect 45468 29792 45520 29844
rect 48320 29835 48372 29844
rect 48320 29801 48329 29835
rect 48329 29801 48363 29835
rect 48363 29801 48372 29835
rect 48320 29792 48372 29801
rect 30840 29724 30892 29776
rect 30932 29699 30984 29708
rect 22928 29588 22980 29640
rect 23848 29631 23900 29640
rect 23848 29597 23857 29631
rect 23857 29597 23891 29631
rect 23891 29597 23900 29631
rect 23848 29588 23900 29597
rect 24400 29631 24452 29640
rect 24400 29597 24409 29631
rect 24409 29597 24443 29631
rect 24443 29597 24452 29631
rect 24400 29588 24452 29597
rect 30932 29665 30941 29699
rect 30941 29665 30975 29699
rect 30975 29665 30984 29699
rect 30932 29656 30984 29665
rect 32680 29699 32732 29708
rect 32680 29665 32689 29699
rect 32689 29665 32723 29699
rect 32723 29665 32732 29699
rect 32680 29656 32732 29665
rect 32772 29699 32824 29708
rect 32772 29665 32781 29699
rect 32781 29665 32815 29699
rect 32815 29665 32824 29699
rect 32772 29656 32824 29665
rect 24768 29631 24820 29640
rect 24768 29597 24777 29631
rect 24777 29597 24811 29631
rect 24811 29597 24820 29631
rect 27712 29631 27764 29640
rect 24768 29588 24820 29597
rect 27712 29597 27721 29631
rect 27721 29597 27755 29631
rect 27755 29597 27764 29631
rect 27712 29588 27764 29597
rect 27896 29588 27948 29640
rect 28080 29588 28132 29640
rect 30380 29588 30432 29640
rect 30656 29588 30708 29640
rect 36452 29631 36504 29640
rect 36452 29597 36461 29631
rect 36461 29597 36495 29631
rect 36495 29597 36504 29631
rect 36452 29588 36504 29597
rect 36636 29631 36688 29640
rect 36636 29597 36645 29631
rect 36645 29597 36679 29631
rect 36679 29597 36688 29631
rect 36636 29588 36688 29597
rect 44272 29656 44324 29708
rect 40408 29631 40460 29640
rect 13728 29452 13780 29504
rect 14096 29452 14148 29504
rect 15476 29452 15528 29504
rect 17592 29452 17644 29504
rect 22376 29452 22428 29504
rect 24124 29452 24176 29504
rect 27160 29452 27212 29504
rect 40408 29597 40417 29631
rect 40417 29597 40451 29631
rect 40451 29597 40460 29631
rect 40408 29588 40460 29597
rect 40592 29588 40644 29640
rect 45008 29631 45060 29640
rect 45008 29597 45017 29631
rect 45017 29597 45051 29631
rect 45051 29597 45060 29631
rect 45008 29588 45060 29597
rect 55220 29656 55272 29708
rect 47676 29631 47728 29640
rect 47676 29597 47685 29631
rect 47685 29597 47719 29631
rect 47719 29597 47728 29631
rect 47676 29588 47728 29597
rect 48044 29588 48096 29640
rect 48504 29631 48556 29640
rect 48504 29597 48513 29631
rect 48513 29597 48547 29631
rect 48547 29597 48556 29631
rect 48504 29588 48556 29597
rect 48780 29631 48832 29640
rect 48780 29597 48789 29631
rect 48789 29597 48823 29631
rect 48823 29597 48832 29631
rect 48780 29588 48832 29597
rect 52092 29631 52144 29640
rect 52092 29597 52101 29631
rect 52101 29597 52135 29631
rect 52135 29597 52144 29631
rect 52092 29588 52144 29597
rect 53012 29631 53064 29640
rect 53012 29597 53021 29631
rect 53021 29597 53055 29631
rect 53055 29597 53064 29631
rect 53012 29588 53064 29597
rect 55312 29631 55364 29640
rect 55312 29597 55321 29631
rect 55321 29597 55355 29631
rect 55355 29597 55364 29631
rect 55312 29588 55364 29597
rect 55680 29631 55732 29640
rect 55680 29597 55689 29631
rect 55689 29597 55723 29631
rect 55723 29597 55732 29631
rect 55680 29588 55732 29597
rect 56324 29631 56376 29640
rect 56324 29597 56333 29631
rect 56333 29597 56367 29631
rect 56367 29597 56376 29631
rect 56324 29588 56376 29597
rect 56968 29588 57020 29640
rect 43076 29520 43128 29572
rect 51540 29563 51592 29572
rect 51540 29529 51549 29563
rect 51549 29529 51583 29563
rect 51583 29529 51592 29563
rect 51540 29520 51592 29529
rect 56048 29520 56100 29572
rect 57704 29588 57756 29640
rect 57888 29588 57940 29640
rect 28172 29452 28224 29504
rect 32312 29495 32364 29504
rect 32312 29461 32321 29495
rect 32321 29461 32355 29495
rect 32355 29461 32364 29495
rect 32312 29452 32364 29461
rect 40500 29495 40552 29504
rect 40500 29461 40509 29495
rect 40509 29461 40543 29495
rect 40543 29461 40552 29495
rect 40500 29452 40552 29461
rect 42432 29452 42484 29504
rect 19574 29350 19626 29402
rect 19638 29350 19690 29402
rect 19702 29350 19754 29402
rect 19766 29350 19818 29402
rect 19830 29350 19882 29402
rect 50294 29350 50346 29402
rect 50358 29350 50410 29402
rect 50422 29350 50474 29402
rect 50486 29350 50538 29402
rect 50550 29350 50602 29402
rect 4344 29180 4396 29232
rect 6920 29223 6972 29232
rect 6920 29189 6929 29223
rect 6929 29189 6963 29223
rect 6963 29189 6972 29223
rect 6920 29180 6972 29189
rect 7472 29248 7524 29300
rect 9128 29180 9180 29232
rect 3332 29112 3384 29164
rect 8944 29112 8996 29164
rect 10508 29180 10560 29232
rect 10600 29155 10652 29164
rect 10600 29121 10609 29155
rect 10609 29121 10643 29155
rect 10643 29121 10652 29155
rect 10600 29112 10652 29121
rect 5724 29044 5776 29096
rect 9772 29044 9824 29096
rect 9864 28976 9916 29028
rect 10416 28976 10468 29028
rect 11152 29112 11204 29164
rect 12624 29248 12676 29300
rect 13084 29248 13136 29300
rect 13452 29248 13504 29300
rect 14096 29248 14148 29300
rect 15568 29248 15620 29300
rect 21180 29291 21232 29300
rect 21180 29257 21189 29291
rect 21189 29257 21223 29291
rect 21223 29257 21232 29291
rect 21180 29248 21232 29257
rect 23112 29248 23164 29300
rect 24860 29248 24912 29300
rect 17040 29180 17092 29232
rect 13912 29112 13964 29164
rect 14648 29155 14700 29164
rect 14648 29121 14657 29155
rect 14657 29121 14691 29155
rect 14691 29121 14700 29155
rect 14648 29112 14700 29121
rect 14740 29155 14792 29164
rect 14740 29121 14749 29155
rect 14749 29121 14783 29155
rect 14783 29121 14792 29155
rect 14740 29112 14792 29121
rect 14924 29112 14976 29164
rect 15476 29155 15528 29164
rect 15476 29121 15485 29155
rect 15485 29121 15519 29155
rect 15519 29121 15528 29155
rect 15476 29112 15528 29121
rect 17960 29180 18012 29232
rect 19156 29223 19208 29232
rect 19156 29189 19165 29223
rect 19165 29189 19199 29223
rect 19199 29189 19208 29223
rect 19156 29180 19208 29189
rect 19432 29180 19484 29232
rect 17592 29112 17644 29164
rect 19248 29112 19300 29164
rect 27068 29180 27120 29232
rect 22744 29112 22796 29164
rect 13636 28976 13688 29028
rect 13728 28976 13780 29028
rect 7380 28908 7432 28960
rect 11980 28908 12032 28960
rect 14188 28976 14240 29028
rect 18604 29044 18656 29096
rect 24124 29087 24176 29096
rect 17224 28976 17276 29028
rect 18052 29019 18104 29028
rect 18052 28985 18061 29019
rect 18061 28985 18095 29019
rect 18095 28985 18104 29019
rect 18052 28976 18104 28985
rect 18512 28976 18564 29028
rect 19340 29019 19392 29028
rect 19340 28985 19349 29019
rect 19349 28985 19383 29019
rect 19383 28985 19392 29019
rect 19340 28976 19392 28985
rect 24124 29053 24133 29087
rect 24133 29053 24167 29087
rect 24167 29053 24176 29087
rect 24124 29044 24176 29053
rect 27160 29155 27212 29164
rect 24584 29044 24636 29096
rect 27160 29121 27169 29155
rect 27169 29121 27203 29155
rect 27203 29121 27212 29155
rect 27160 29112 27212 29121
rect 28080 29112 28132 29164
rect 28172 29155 28224 29164
rect 28172 29121 28181 29155
rect 28181 29121 28215 29155
rect 28215 29121 28224 29155
rect 28172 29112 28224 29121
rect 24308 28976 24360 29028
rect 27712 28976 27764 29028
rect 28264 29044 28316 29096
rect 32220 29248 32272 29300
rect 32680 29248 32732 29300
rect 36452 29248 36504 29300
rect 48780 29248 48832 29300
rect 49608 29291 49660 29300
rect 49608 29257 49617 29291
rect 49617 29257 49651 29291
rect 49651 29257 49660 29291
rect 49608 29248 49660 29257
rect 51724 29291 51776 29300
rect 51724 29257 51733 29291
rect 51733 29257 51767 29291
rect 51767 29257 51776 29291
rect 51724 29248 51776 29257
rect 55312 29248 55364 29300
rect 56324 29248 56376 29300
rect 30932 29112 30984 29164
rect 32220 29155 32272 29164
rect 32220 29121 32229 29155
rect 32229 29121 32263 29155
rect 32263 29121 32272 29155
rect 32220 29112 32272 29121
rect 34520 29112 34572 29164
rect 43076 29155 43128 29164
rect 43076 29121 43085 29155
rect 43085 29121 43119 29155
rect 43119 29121 43128 29155
rect 43076 29112 43128 29121
rect 33140 29044 33192 29096
rect 42892 29087 42944 29096
rect 42892 29053 42901 29087
rect 42901 29053 42935 29087
rect 42935 29053 42944 29087
rect 42892 29044 42944 29053
rect 45008 29180 45060 29232
rect 47676 29180 47728 29232
rect 45468 29112 45520 29164
rect 49148 29112 49200 29164
rect 29276 28976 29328 29028
rect 45192 29044 45244 29096
rect 48504 29087 48556 29096
rect 48504 29053 48513 29087
rect 48513 29053 48547 29087
rect 48547 29053 48556 29087
rect 48504 29044 48556 29053
rect 51080 29180 51132 29232
rect 48412 28976 48464 29028
rect 50896 29112 50948 29164
rect 57612 29180 57664 29232
rect 56048 29112 56100 29164
rect 57888 29112 57940 29164
rect 58164 29155 58216 29164
rect 58164 29121 58173 29155
rect 58173 29121 58207 29155
rect 58207 29121 58216 29155
rect 58164 29112 58216 29121
rect 55772 29044 55824 29096
rect 57704 29044 57756 29096
rect 22468 28908 22520 28960
rect 27620 28951 27672 28960
rect 27620 28917 27629 28951
rect 27629 28917 27663 28951
rect 27663 28917 27672 28951
rect 27620 28908 27672 28917
rect 27896 28908 27948 28960
rect 28632 28908 28684 28960
rect 48044 28908 48096 28960
rect 57428 28976 57480 29028
rect 56968 28908 57020 28960
rect 4214 28806 4266 28858
rect 4278 28806 4330 28858
rect 4342 28806 4394 28858
rect 4406 28806 4458 28858
rect 4470 28806 4522 28858
rect 34934 28806 34986 28858
rect 34998 28806 35050 28858
rect 35062 28806 35114 28858
rect 35126 28806 35178 28858
rect 35190 28806 35242 28858
rect 10600 28704 10652 28756
rect 10784 28704 10836 28756
rect 12164 28704 12216 28756
rect 12348 28704 12400 28756
rect 18788 28704 18840 28756
rect 24860 28704 24912 28756
rect 42524 28747 42576 28756
rect 9864 28636 9916 28688
rect 10692 28636 10744 28688
rect 22744 28636 22796 28688
rect 23848 28636 23900 28688
rect 24768 28636 24820 28688
rect 8944 28543 8996 28552
rect 8944 28509 8953 28543
rect 8953 28509 8987 28543
rect 8987 28509 8996 28543
rect 8944 28500 8996 28509
rect 9128 28543 9180 28552
rect 9128 28509 9137 28543
rect 9137 28509 9171 28543
rect 9171 28509 9180 28543
rect 9128 28500 9180 28509
rect 9680 28543 9732 28552
rect 9680 28509 9689 28543
rect 9689 28509 9723 28543
rect 9723 28509 9732 28543
rect 9680 28500 9732 28509
rect 11980 28611 12032 28620
rect 11980 28577 11989 28611
rect 11989 28577 12023 28611
rect 12023 28577 12032 28611
rect 11980 28568 12032 28577
rect 11152 28543 11204 28552
rect 11152 28509 11161 28543
rect 11161 28509 11195 28543
rect 11195 28509 11204 28543
rect 11152 28500 11204 28509
rect 11428 28500 11480 28552
rect 12164 28500 12216 28552
rect 6736 28432 6788 28484
rect 7012 28407 7064 28416
rect 7012 28373 7021 28407
rect 7021 28373 7055 28407
rect 7055 28373 7064 28407
rect 7012 28364 7064 28373
rect 10508 28432 10560 28484
rect 10692 28432 10744 28484
rect 17132 28568 17184 28620
rect 13452 28500 13504 28552
rect 13728 28500 13780 28552
rect 15016 28500 15068 28552
rect 14556 28407 14608 28416
rect 14556 28373 14565 28407
rect 14565 28373 14599 28407
rect 14599 28373 14608 28407
rect 14556 28364 14608 28373
rect 18604 28500 18656 28552
rect 19340 28500 19392 28552
rect 21088 28568 21140 28620
rect 22284 28568 22336 28620
rect 22468 28543 22520 28552
rect 19432 28432 19484 28484
rect 22468 28509 22477 28543
rect 22477 28509 22511 28543
rect 22511 28509 22520 28543
rect 22468 28500 22520 28509
rect 23664 28543 23716 28552
rect 23664 28509 23673 28543
rect 23673 28509 23707 28543
rect 23707 28509 23716 28543
rect 23664 28500 23716 28509
rect 24308 28500 24360 28552
rect 24584 28500 24636 28552
rect 22008 28432 22060 28484
rect 22100 28432 22152 28484
rect 22560 28432 22612 28484
rect 27620 28636 27672 28688
rect 32312 28636 32364 28688
rect 36636 28636 36688 28688
rect 39672 28636 39724 28688
rect 42524 28713 42533 28747
rect 42533 28713 42567 28747
rect 42567 28713 42576 28747
rect 42524 28704 42576 28713
rect 48504 28747 48556 28756
rect 48504 28713 48513 28747
rect 48513 28713 48547 28747
rect 48547 28713 48556 28747
rect 48504 28704 48556 28713
rect 51264 28704 51316 28756
rect 57888 28704 57940 28756
rect 58164 28747 58216 28756
rect 58164 28713 58173 28747
rect 58173 28713 58207 28747
rect 58207 28713 58216 28747
rect 58164 28704 58216 28713
rect 57796 28636 57848 28688
rect 27804 28568 27856 28620
rect 34612 28568 34664 28620
rect 37556 28611 37608 28620
rect 37556 28577 37565 28611
rect 37565 28577 37599 28611
rect 37599 28577 37608 28611
rect 37556 28568 37608 28577
rect 20076 28364 20128 28416
rect 22836 28407 22888 28416
rect 22836 28373 22845 28407
rect 22845 28373 22879 28407
rect 22879 28373 22888 28407
rect 22836 28364 22888 28373
rect 27252 28407 27304 28416
rect 27252 28373 27261 28407
rect 27261 28373 27295 28407
rect 27295 28373 27304 28407
rect 27252 28364 27304 28373
rect 27712 28364 27764 28416
rect 28264 28500 28316 28552
rect 35348 28500 35400 28552
rect 37740 28543 37792 28552
rect 37740 28509 37749 28543
rect 37749 28509 37783 28543
rect 37783 28509 37792 28543
rect 37740 28500 37792 28509
rect 28540 28407 28592 28416
rect 28540 28373 28549 28407
rect 28549 28373 28583 28407
rect 28583 28373 28592 28407
rect 28540 28364 28592 28373
rect 30380 28364 30432 28416
rect 31392 28475 31444 28484
rect 31392 28441 31401 28475
rect 31401 28441 31435 28475
rect 31435 28441 31444 28475
rect 31392 28432 31444 28441
rect 39120 28568 39172 28620
rect 42892 28568 42944 28620
rect 45192 28568 45244 28620
rect 39304 28500 39356 28552
rect 42340 28543 42392 28552
rect 42340 28509 42349 28543
rect 42349 28509 42383 28543
rect 42383 28509 42392 28543
rect 42340 28500 42392 28509
rect 45468 28543 45520 28552
rect 45468 28509 45477 28543
rect 45477 28509 45511 28543
rect 45511 28509 45520 28543
rect 45468 28500 45520 28509
rect 51356 28568 51408 28620
rect 48044 28543 48096 28552
rect 48044 28509 48053 28543
rect 48053 28509 48087 28543
rect 48087 28509 48096 28543
rect 48044 28500 48096 28509
rect 48320 28543 48372 28552
rect 48320 28509 48329 28543
rect 48329 28509 48363 28543
rect 48363 28509 48372 28543
rect 48320 28500 48372 28509
rect 49332 28500 49384 28552
rect 49608 28543 49660 28552
rect 49608 28509 49617 28543
rect 49617 28509 49651 28543
rect 49651 28509 49660 28543
rect 49608 28500 49660 28509
rect 57244 28500 57296 28552
rect 57428 28543 57480 28552
rect 57428 28509 57437 28543
rect 57437 28509 57471 28543
rect 57471 28509 57480 28543
rect 57428 28500 57480 28509
rect 47676 28432 47728 28484
rect 51264 28475 51316 28484
rect 51264 28441 51273 28475
rect 51273 28441 51307 28475
rect 51307 28441 51316 28475
rect 51264 28432 51316 28441
rect 41880 28407 41932 28416
rect 41880 28373 41889 28407
rect 41889 28373 41923 28407
rect 41923 28373 41932 28407
rect 41880 28364 41932 28373
rect 51632 28364 51684 28416
rect 56048 28364 56100 28416
rect 57980 28364 58032 28416
rect 19574 28262 19626 28314
rect 19638 28262 19690 28314
rect 19702 28262 19754 28314
rect 19766 28262 19818 28314
rect 19830 28262 19882 28314
rect 50294 28262 50346 28314
rect 50358 28262 50410 28314
rect 50422 28262 50474 28314
rect 50486 28262 50538 28314
rect 50550 28262 50602 28314
rect 7012 28092 7064 28144
rect 13728 28160 13780 28212
rect 13820 28160 13872 28212
rect 25412 28203 25464 28212
rect 25412 28169 25421 28203
rect 25421 28169 25455 28203
rect 25455 28169 25464 28203
rect 25412 28160 25464 28169
rect 32220 28160 32272 28212
rect 37740 28160 37792 28212
rect 43076 28160 43128 28212
rect 51356 28160 51408 28212
rect 55680 28160 55732 28212
rect 56968 28203 57020 28212
rect 56968 28169 56977 28203
rect 56977 28169 57011 28203
rect 57011 28169 57020 28203
rect 56968 28160 57020 28169
rect 8208 28092 8260 28144
rect 10416 28092 10468 28144
rect 2964 27956 3016 28008
rect 3056 27999 3108 28008
rect 3056 27965 3065 27999
rect 3065 27965 3099 27999
rect 3099 27965 3108 27999
rect 3056 27956 3108 27965
rect 3332 27956 3384 28008
rect 8484 28024 8536 28076
rect 9680 28024 9732 28076
rect 15108 28092 15160 28144
rect 19248 28092 19300 28144
rect 24768 28092 24820 28144
rect 27804 28092 27856 28144
rect 14004 28024 14056 28076
rect 8944 27956 8996 28008
rect 13728 27956 13780 28008
rect 15200 28024 15252 28076
rect 16212 28024 16264 28076
rect 17040 28024 17092 28076
rect 17224 28067 17276 28076
rect 17224 28033 17233 28067
rect 17233 28033 17267 28067
rect 17267 28033 17276 28067
rect 17224 28024 17276 28033
rect 22284 28024 22336 28076
rect 24124 28024 24176 28076
rect 4896 27888 4948 27940
rect 8024 27888 8076 27940
rect 10508 27888 10560 27940
rect 14464 27888 14516 27940
rect 6460 27820 6512 27872
rect 6736 27863 6788 27872
rect 6736 27829 6745 27863
rect 6745 27829 6779 27863
rect 6779 27829 6788 27863
rect 6736 27820 6788 27829
rect 7472 27863 7524 27872
rect 7472 27829 7481 27863
rect 7481 27829 7515 27863
rect 7515 27829 7524 27863
rect 7472 27820 7524 27829
rect 12256 27820 12308 27872
rect 15200 27820 15252 27872
rect 22008 27999 22060 28008
rect 22008 27965 22017 27999
rect 22017 27965 22051 27999
rect 22051 27965 22060 27999
rect 22008 27956 22060 27965
rect 23664 27956 23716 28008
rect 24216 27956 24268 28008
rect 25136 28024 25188 28076
rect 30748 28024 30800 28076
rect 31392 28024 31444 28076
rect 36360 28067 36412 28076
rect 36360 28033 36369 28067
rect 36369 28033 36403 28067
rect 36403 28033 36412 28067
rect 36360 28024 36412 28033
rect 36452 28024 36504 28076
rect 39120 28067 39172 28076
rect 39120 28033 39129 28067
rect 39129 28033 39163 28067
rect 39163 28033 39172 28067
rect 39120 28024 39172 28033
rect 39304 28067 39356 28076
rect 39304 28033 39313 28067
rect 39313 28033 39347 28067
rect 39347 28033 39356 28067
rect 39304 28024 39356 28033
rect 41052 28067 41104 28076
rect 41052 28033 41061 28067
rect 41061 28033 41095 28067
rect 41095 28033 41104 28067
rect 41052 28024 41104 28033
rect 41144 28067 41196 28076
rect 41144 28033 41153 28067
rect 41153 28033 41187 28067
rect 41187 28033 41196 28067
rect 41328 28067 41380 28076
rect 41144 28024 41196 28033
rect 41328 28033 41337 28067
rect 41337 28033 41371 28067
rect 41371 28033 41380 28067
rect 41328 28024 41380 28033
rect 30380 27956 30432 28008
rect 41236 27956 41288 28008
rect 41880 28024 41932 28076
rect 57244 28092 57296 28144
rect 57428 28092 57480 28144
rect 42340 27956 42392 28008
rect 42892 28024 42944 28076
rect 44916 28024 44968 28076
rect 51080 28067 51132 28076
rect 51080 28033 51089 28067
rect 51089 28033 51123 28067
rect 51123 28033 51132 28067
rect 51080 28024 51132 28033
rect 45008 27999 45060 28008
rect 45008 27965 45017 27999
rect 45017 27965 45051 27999
rect 45051 27965 45060 27999
rect 45008 27956 45060 27965
rect 17132 27888 17184 27940
rect 37648 27888 37700 27940
rect 45100 27888 45152 27940
rect 18052 27820 18104 27872
rect 24216 27863 24268 27872
rect 24216 27829 24225 27863
rect 24225 27829 24259 27863
rect 24259 27829 24268 27863
rect 24216 27820 24268 27829
rect 25044 27820 25096 27872
rect 29644 27863 29696 27872
rect 29644 27829 29653 27863
rect 29653 27829 29687 27863
rect 29687 27829 29696 27863
rect 29644 27820 29696 27829
rect 30380 27863 30432 27872
rect 30380 27829 30389 27863
rect 30389 27829 30423 27863
rect 30423 27829 30432 27863
rect 30380 27820 30432 27829
rect 46848 27820 46900 27872
rect 51356 28067 51408 28076
rect 51356 28033 51365 28067
rect 51365 28033 51399 28067
rect 51399 28033 51408 28067
rect 51356 28024 51408 28033
rect 51632 28024 51684 28076
rect 55312 28024 55364 28076
rect 55588 28067 55640 28076
rect 55588 28033 55597 28067
rect 55597 28033 55631 28067
rect 55631 28033 55640 28067
rect 55588 28024 55640 28033
rect 55864 28024 55916 28076
rect 55772 27999 55824 28008
rect 55772 27965 55781 27999
rect 55781 27965 55815 27999
rect 55815 27965 55824 27999
rect 55772 27956 55824 27965
rect 56968 27888 57020 27940
rect 51448 27820 51500 27872
rect 51724 27863 51776 27872
rect 51724 27829 51733 27863
rect 51733 27829 51767 27863
rect 51767 27829 51776 27863
rect 51724 27820 51776 27829
rect 57980 27820 58032 27872
rect 4214 27718 4266 27770
rect 4278 27718 4330 27770
rect 4342 27718 4394 27770
rect 4406 27718 4458 27770
rect 4470 27718 4522 27770
rect 34934 27718 34986 27770
rect 34998 27718 35050 27770
rect 35062 27718 35114 27770
rect 35126 27718 35178 27770
rect 35190 27718 35242 27770
rect 3056 27616 3108 27668
rect 27252 27616 27304 27668
rect 41052 27616 41104 27668
rect 45468 27659 45520 27668
rect 2044 27591 2096 27600
rect 2044 27557 2053 27591
rect 2053 27557 2087 27591
rect 2087 27557 2096 27591
rect 2044 27548 2096 27557
rect 2780 27480 2832 27532
rect 3976 27412 4028 27464
rect 5540 27412 5592 27464
rect 5632 27387 5684 27396
rect 5632 27353 5641 27387
rect 5641 27353 5675 27387
rect 5675 27353 5684 27387
rect 5632 27344 5684 27353
rect 7472 27548 7524 27600
rect 13268 27548 13320 27600
rect 14372 27548 14424 27600
rect 15292 27591 15344 27600
rect 15292 27557 15301 27591
rect 15301 27557 15335 27591
rect 15335 27557 15344 27591
rect 15292 27548 15344 27557
rect 17040 27591 17092 27600
rect 11244 27480 11296 27532
rect 6460 27455 6512 27464
rect 6460 27421 6469 27455
rect 6469 27421 6503 27455
rect 6503 27421 6512 27455
rect 6460 27412 6512 27421
rect 8024 27412 8076 27464
rect 8484 27412 8536 27464
rect 8944 27412 8996 27464
rect 11796 27412 11848 27464
rect 13084 27455 13136 27464
rect 6276 27276 6328 27328
rect 7196 27276 7248 27328
rect 8116 27276 8168 27328
rect 10692 27387 10744 27396
rect 10692 27353 10701 27387
rect 10701 27353 10735 27387
rect 10735 27353 10744 27387
rect 10692 27344 10744 27353
rect 13084 27421 13093 27455
rect 13093 27421 13127 27455
rect 13127 27421 13136 27455
rect 13084 27412 13136 27421
rect 14280 27455 14332 27464
rect 14280 27421 14289 27455
rect 14289 27421 14323 27455
rect 14323 27421 14332 27455
rect 14280 27412 14332 27421
rect 16764 27480 16816 27532
rect 14464 27455 14516 27464
rect 14464 27421 14473 27455
rect 14473 27421 14507 27455
rect 14507 27421 14516 27455
rect 14464 27412 14516 27421
rect 17040 27557 17049 27591
rect 17049 27557 17083 27591
rect 17083 27557 17092 27591
rect 17040 27548 17092 27557
rect 17592 27591 17644 27600
rect 17592 27557 17601 27591
rect 17601 27557 17635 27591
rect 17635 27557 17644 27591
rect 17592 27548 17644 27557
rect 22836 27548 22888 27600
rect 30932 27591 30984 27600
rect 16948 27480 17000 27532
rect 20352 27480 20404 27532
rect 22008 27480 22060 27532
rect 22284 27480 22336 27532
rect 20168 27412 20220 27464
rect 20812 27412 20864 27464
rect 25044 27523 25096 27532
rect 25044 27489 25053 27523
rect 25053 27489 25087 27523
rect 25087 27489 25096 27523
rect 25044 27480 25096 27489
rect 8944 27319 8996 27328
rect 8944 27285 8953 27319
rect 8953 27285 8987 27319
rect 8987 27285 8996 27319
rect 17960 27344 18012 27396
rect 23664 27455 23716 27464
rect 23664 27421 23673 27455
rect 23673 27421 23707 27455
rect 23707 27421 23716 27455
rect 23664 27412 23716 27421
rect 25136 27455 25188 27464
rect 25136 27421 25145 27455
rect 25145 27421 25179 27455
rect 25179 27421 25188 27455
rect 25136 27412 25188 27421
rect 26148 27455 26200 27464
rect 26148 27421 26157 27455
rect 26157 27421 26191 27455
rect 26191 27421 26200 27455
rect 26148 27412 26200 27421
rect 27436 27412 27488 27464
rect 28080 27455 28132 27464
rect 28080 27421 28089 27455
rect 28089 27421 28123 27455
rect 28123 27421 28132 27455
rect 28080 27412 28132 27421
rect 28540 27412 28592 27464
rect 30932 27557 30941 27591
rect 30941 27557 30975 27591
rect 30975 27557 30984 27591
rect 30932 27548 30984 27557
rect 32864 27548 32916 27600
rect 29644 27412 29696 27464
rect 30748 27455 30800 27464
rect 30748 27421 30757 27455
rect 30757 27421 30791 27455
rect 30791 27421 30800 27455
rect 30748 27412 30800 27421
rect 8944 27276 8996 27285
rect 17316 27276 17368 27328
rect 26884 27344 26936 27396
rect 34520 27480 34572 27532
rect 34704 27480 34756 27532
rect 36360 27548 36412 27600
rect 39304 27548 39356 27600
rect 45468 27625 45477 27659
rect 45477 27625 45511 27659
rect 45511 27625 45520 27659
rect 45468 27616 45520 27625
rect 48320 27616 48372 27668
rect 49148 27616 49200 27668
rect 51264 27616 51316 27668
rect 38108 27523 38160 27532
rect 38108 27489 38117 27523
rect 38117 27489 38151 27523
rect 38151 27489 38160 27523
rect 38108 27480 38160 27489
rect 36452 27455 36504 27464
rect 36452 27421 36461 27455
rect 36461 27421 36495 27455
rect 36495 27421 36504 27455
rect 38200 27455 38252 27464
rect 36452 27412 36504 27421
rect 38200 27421 38209 27455
rect 38209 27421 38243 27455
rect 38243 27421 38252 27455
rect 38200 27412 38252 27421
rect 41236 27523 41288 27532
rect 41236 27489 41245 27523
rect 41245 27489 41279 27523
rect 41279 27489 41288 27523
rect 41236 27480 41288 27489
rect 48044 27548 48096 27600
rect 45100 27523 45152 27532
rect 40868 27412 40920 27464
rect 41328 27455 41380 27464
rect 41328 27421 41337 27455
rect 41337 27421 41371 27455
rect 41371 27421 41380 27455
rect 41328 27412 41380 27421
rect 18880 27276 18932 27328
rect 19248 27276 19300 27328
rect 22744 27276 22796 27328
rect 22928 27276 22980 27328
rect 23388 27319 23440 27328
rect 23388 27285 23397 27319
rect 23397 27285 23431 27319
rect 23431 27285 23440 27319
rect 23388 27276 23440 27285
rect 26240 27319 26292 27328
rect 26240 27285 26249 27319
rect 26249 27285 26283 27319
rect 26283 27285 26292 27319
rect 26240 27276 26292 27285
rect 28632 27276 28684 27328
rect 28724 27276 28776 27328
rect 41144 27344 41196 27396
rect 45100 27489 45109 27523
rect 45109 27489 45143 27523
rect 45143 27489 45152 27523
rect 45100 27480 45152 27489
rect 46848 27480 46900 27532
rect 51908 27548 51960 27600
rect 52368 27591 52420 27600
rect 52368 27557 52377 27591
rect 52377 27557 52411 27591
rect 52411 27557 52420 27591
rect 52368 27548 52420 27557
rect 56968 27591 57020 27600
rect 44916 27412 44968 27464
rect 47400 27455 47452 27464
rect 47400 27421 47409 27455
rect 47409 27421 47443 27455
rect 47443 27421 47452 27455
rect 47400 27412 47452 27421
rect 49148 27455 49200 27464
rect 49148 27421 49157 27455
rect 49157 27421 49191 27455
rect 49191 27421 49200 27455
rect 49148 27412 49200 27421
rect 49332 27455 49384 27464
rect 49332 27421 49341 27455
rect 49341 27421 49375 27455
rect 49375 27421 49384 27455
rect 49332 27412 49384 27421
rect 50712 27412 50764 27464
rect 51264 27455 51316 27464
rect 37556 27276 37608 27328
rect 42340 27276 42392 27328
rect 47400 27276 47452 27328
rect 47952 27344 48004 27396
rect 51264 27421 51273 27455
rect 51273 27421 51307 27455
rect 51307 27421 51316 27455
rect 51264 27412 51316 27421
rect 51724 27412 51776 27464
rect 53932 27412 53984 27464
rect 55312 27455 55364 27464
rect 55312 27421 55321 27455
rect 55321 27421 55355 27455
rect 55355 27421 55364 27455
rect 55312 27412 55364 27421
rect 55956 27480 56008 27532
rect 56968 27557 56977 27591
rect 56977 27557 57011 27591
rect 57011 27557 57020 27591
rect 56968 27548 57020 27557
rect 55588 27412 55640 27464
rect 56600 27455 56652 27464
rect 51356 27344 51408 27396
rect 52644 27344 52696 27396
rect 55128 27344 55180 27396
rect 56600 27421 56609 27455
rect 56609 27421 56643 27455
rect 56643 27421 56652 27455
rect 56600 27412 56652 27421
rect 58164 27455 58216 27464
rect 58164 27421 58173 27455
rect 58173 27421 58207 27455
rect 58207 27421 58216 27455
rect 58164 27412 58216 27421
rect 51172 27276 51224 27328
rect 56876 27276 56928 27328
rect 19574 27174 19626 27226
rect 19638 27174 19690 27226
rect 19702 27174 19754 27226
rect 19766 27174 19818 27226
rect 19830 27174 19882 27226
rect 50294 27174 50346 27226
rect 50358 27174 50410 27226
rect 50422 27174 50474 27226
rect 50486 27174 50538 27226
rect 50550 27174 50602 27226
rect 5632 27072 5684 27124
rect 6644 27072 6696 27124
rect 7288 27072 7340 27124
rect 1860 27047 1912 27056
rect 1860 27013 1869 27047
rect 1869 27013 1903 27047
rect 1903 27013 1912 27047
rect 1860 27004 1912 27013
rect 6736 27004 6788 27056
rect 10140 27072 10192 27124
rect 14648 27072 14700 27124
rect 15108 27115 15160 27124
rect 15108 27081 15117 27115
rect 15117 27081 15151 27115
rect 15151 27081 15160 27115
rect 15108 27072 15160 27081
rect 15476 27072 15528 27124
rect 18420 27072 18472 27124
rect 19064 27115 19116 27124
rect 19064 27081 19073 27115
rect 19073 27081 19107 27115
rect 19107 27081 19116 27115
rect 19064 27072 19116 27081
rect 19984 27072 20036 27124
rect 30564 27072 30616 27124
rect 36452 27072 36504 27124
rect 40868 27072 40920 27124
rect 41328 27115 41380 27124
rect 41328 27081 41337 27115
rect 41337 27081 41371 27115
rect 41371 27081 41380 27115
rect 41328 27072 41380 27081
rect 44916 27072 44968 27124
rect 45008 27072 45060 27124
rect 51264 27072 51316 27124
rect 56600 27072 56652 27124
rect 58164 27115 58216 27124
rect 58164 27081 58173 27115
rect 58173 27081 58207 27115
rect 58207 27081 58216 27115
rect 58164 27072 58216 27081
rect 8024 27047 8076 27056
rect 6828 26979 6880 26988
rect 6828 26945 6837 26979
rect 6837 26945 6871 26979
rect 6871 26945 6880 26979
rect 6828 26936 6880 26945
rect 8024 27013 8051 27047
rect 8051 27013 8076 27047
rect 8024 27004 8076 27013
rect 10048 27047 10100 27056
rect 7104 26979 7156 26988
rect 7104 26945 7113 26979
rect 7113 26945 7147 26979
rect 7147 26945 7156 26979
rect 7104 26936 7156 26945
rect 8116 26936 8168 26988
rect 6276 26868 6328 26920
rect 10048 27013 10057 27047
rect 10057 27013 10091 27047
rect 10091 27013 10100 27047
rect 10048 27004 10100 27013
rect 9772 26936 9824 26988
rect 12256 27004 12308 27056
rect 13268 27004 13320 27056
rect 11428 26936 11480 26988
rect 13820 26979 13872 26988
rect 13820 26945 13829 26979
rect 13829 26945 13863 26979
rect 13863 26945 13872 26979
rect 14464 26979 14516 26988
rect 13820 26936 13872 26945
rect 14464 26945 14473 26979
rect 14473 26945 14507 26979
rect 14507 26945 14516 26979
rect 14464 26936 14516 26945
rect 14556 26979 14608 26988
rect 14556 26945 14566 26979
rect 14566 26945 14600 26979
rect 14600 26945 14608 26979
rect 16028 27004 16080 27056
rect 18696 27004 18748 27056
rect 24768 27004 24820 27056
rect 26240 27004 26292 27056
rect 27436 27047 27488 27056
rect 27436 27013 27445 27047
rect 27445 27013 27479 27047
rect 27479 27013 27488 27047
rect 27436 27004 27488 27013
rect 28632 27004 28684 27056
rect 38200 27004 38252 27056
rect 39948 27004 40000 27056
rect 14556 26936 14608 26945
rect 13544 26868 13596 26920
rect 14280 26868 14332 26920
rect 14648 26868 14700 26920
rect 14924 26936 14976 26988
rect 16488 26936 16540 26988
rect 20536 26936 20588 26988
rect 22192 26936 22244 26988
rect 22836 26936 22888 26988
rect 23664 26936 23716 26988
rect 15292 26868 15344 26920
rect 20168 26868 20220 26920
rect 20352 26911 20404 26920
rect 20352 26877 20361 26911
rect 20361 26877 20395 26911
rect 20395 26877 20404 26911
rect 20352 26868 20404 26877
rect 5448 26800 5500 26852
rect 11888 26843 11940 26852
rect 11888 26809 11897 26843
rect 11897 26809 11931 26843
rect 11931 26809 11940 26843
rect 11888 26800 11940 26809
rect 6644 26732 6696 26784
rect 9864 26732 9916 26784
rect 10324 26732 10376 26784
rect 15016 26800 15068 26852
rect 19248 26800 19300 26852
rect 17960 26732 18012 26784
rect 18420 26732 18472 26784
rect 21180 26868 21232 26920
rect 21640 26868 21692 26920
rect 26884 26868 26936 26920
rect 28540 26936 28592 26988
rect 32864 26936 32916 26988
rect 35348 26936 35400 26988
rect 37648 26936 37700 26988
rect 38108 26936 38160 26988
rect 40224 26979 40276 26988
rect 40224 26945 40233 26979
rect 40233 26945 40267 26979
rect 40267 26945 40276 26979
rect 40224 26936 40276 26945
rect 40500 26979 40552 26988
rect 40500 26945 40509 26979
rect 40509 26945 40543 26979
rect 40543 26945 40552 26979
rect 44272 26979 44324 26988
rect 40500 26936 40552 26945
rect 44272 26945 44281 26979
rect 44281 26945 44315 26979
rect 44315 26945 44324 26979
rect 51172 27004 51224 27056
rect 51356 27004 51408 27056
rect 55312 27004 55364 27056
rect 44272 26936 44324 26945
rect 50896 26979 50948 26988
rect 20720 26800 20772 26852
rect 30472 26868 30524 26920
rect 34520 26868 34572 26920
rect 44180 26911 44232 26920
rect 44180 26877 44189 26911
rect 44189 26877 44223 26911
rect 44223 26877 44232 26911
rect 50896 26945 50905 26979
rect 50905 26945 50939 26979
rect 50939 26945 50948 26979
rect 50896 26936 50948 26945
rect 53380 26979 53432 26988
rect 53380 26945 53389 26979
rect 53389 26945 53423 26979
rect 53423 26945 53432 26979
rect 53380 26936 53432 26945
rect 54024 26936 54076 26988
rect 55128 26936 55180 26988
rect 55956 26979 56008 26988
rect 55956 26945 55965 26979
rect 55965 26945 55999 26979
rect 55999 26945 56008 26979
rect 56968 26979 57020 26988
rect 55956 26936 56008 26945
rect 56968 26945 56977 26979
rect 56977 26945 57011 26979
rect 57011 26945 57020 26979
rect 56968 26936 57020 26945
rect 56876 26911 56928 26920
rect 44180 26868 44232 26877
rect 56876 26877 56885 26911
rect 56885 26877 56919 26911
rect 56919 26877 56928 26911
rect 56876 26868 56928 26877
rect 41052 26800 41104 26852
rect 55864 26800 55916 26852
rect 20628 26775 20680 26784
rect 20628 26741 20637 26775
rect 20637 26741 20671 26775
rect 20671 26741 20680 26775
rect 20628 26732 20680 26741
rect 20812 26732 20864 26784
rect 23572 26732 23624 26784
rect 27896 26732 27948 26784
rect 28080 26732 28132 26784
rect 29552 26775 29604 26784
rect 29552 26741 29561 26775
rect 29561 26741 29595 26775
rect 29595 26741 29604 26775
rect 29552 26732 29604 26741
rect 33600 26732 33652 26784
rect 34796 26732 34848 26784
rect 41144 26775 41196 26784
rect 41144 26741 41153 26775
rect 41153 26741 41187 26775
rect 41187 26741 41196 26775
rect 41144 26732 41196 26741
rect 57888 26732 57940 26784
rect 4214 26630 4266 26682
rect 4278 26630 4330 26682
rect 4342 26630 4394 26682
rect 4406 26630 4458 26682
rect 4470 26630 4522 26682
rect 34934 26630 34986 26682
rect 34998 26630 35050 26682
rect 35062 26630 35114 26682
rect 35126 26630 35178 26682
rect 35190 26630 35242 26682
rect 1860 26528 1912 26580
rect 3148 26528 3200 26580
rect 4068 26528 4120 26580
rect 6828 26528 6880 26580
rect 10968 26528 11020 26580
rect 13544 26528 13596 26580
rect 14096 26571 14148 26580
rect 14096 26537 14105 26571
rect 14105 26537 14139 26571
rect 14139 26537 14148 26571
rect 14096 26528 14148 26537
rect 8024 26460 8076 26512
rect 15200 26460 15252 26512
rect 6644 26392 6696 26444
rect 6276 26367 6328 26376
rect 6276 26333 6285 26367
rect 6285 26333 6319 26367
rect 6319 26333 6328 26367
rect 6276 26324 6328 26333
rect 8024 26324 8076 26376
rect 9864 26324 9916 26376
rect 10140 26367 10192 26376
rect 10140 26333 10149 26367
rect 10149 26333 10183 26367
rect 10183 26333 10192 26367
rect 10140 26324 10192 26333
rect 10324 26324 10376 26376
rect 11888 26392 11940 26444
rect 15016 26435 15068 26444
rect 15016 26401 15025 26435
rect 15025 26401 15059 26435
rect 15059 26401 15068 26435
rect 15016 26392 15068 26401
rect 16764 26324 16816 26376
rect 18144 26528 18196 26580
rect 18696 26571 18748 26580
rect 18696 26537 18705 26571
rect 18705 26537 18739 26571
rect 18739 26537 18748 26571
rect 18696 26528 18748 26537
rect 19064 26528 19116 26580
rect 19616 26528 19668 26580
rect 19984 26528 20036 26580
rect 21456 26528 21508 26580
rect 17684 26460 17736 26512
rect 21088 26460 21140 26512
rect 17316 26367 17368 26376
rect 17316 26333 17325 26367
rect 17325 26333 17359 26367
rect 17359 26333 17368 26367
rect 17316 26324 17368 26333
rect 17684 26324 17736 26376
rect 17776 26324 17828 26376
rect 18144 26367 18196 26376
rect 18144 26333 18154 26367
rect 18154 26333 18188 26367
rect 18188 26333 18196 26367
rect 18420 26367 18472 26376
rect 18144 26324 18196 26333
rect 18420 26333 18429 26367
rect 18429 26333 18463 26367
rect 18463 26333 18472 26367
rect 18420 26324 18472 26333
rect 18696 26324 18748 26376
rect 20628 26392 20680 26444
rect 22744 26460 22796 26512
rect 19340 26367 19392 26376
rect 19340 26333 19350 26367
rect 19350 26333 19384 26367
rect 19384 26333 19392 26367
rect 19340 26324 19392 26333
rect 19708 26324 19760 26376
rect 22836 26392 22888 26444
rect 23388 26392 23440 26444
rect 22192 26367 22244 26376
rect 11244 26299 11296 26308
rect 11244 26265 11253 26299
rect 11253 26265 11287 26299
rect 11287 26265 11296 26299
rect 11244 26256 11296 26265
rect 11428 26299 11480 26308
rect 11428 26265 11437 26299
rect 11437 26265 11471 26299
rect 11471 26265 11480 26299
rect 11428 26256 11480 26265
rect 15200 26256 15252 26308
rect 10232 26188 10284 26240
rect 17408 26188 17460 26240
rect 19616 26299 19668 26308
rect 19616 26265 19625 26299
rect 19625 26265 19659 26299
rect 19659 26265 19668 26299
rect 19616 26256 19668 26265
rect 22192 26333 22201 26367
rect 22201 26333 22235 26367
rect 22235 26333 22244 26367
rect 22192 26324 22244 26333
rect 23296 26367 23348 26376
rect 23296 26333 23305 26367
rect 23305 26333 23339 26367
rect 23339 26333 23348 26367
rect 23296 26324 23348 26333
rect 23572 26367 23624 26376
rect 23572 26333 23581 26367
rect 23581 26333 23615 26367
rect 23615 26333 23624 26367
rect 23572 26324 23624 26333
rect 23940 26324 23992 26376
rect 25136 26528 25188 26580
rect 34428 26528 34480 26580
rect 34796 26571 34848 26580
rect 34796 26537 34805 26571
rect 34805 26537 34839 26571
rect 34839 26537 34848 26571
rect 34796 26528 34848 26537
rect 38200 26528 38252 26580
rect 44272 26528 44324 26580
rect 50712 26571 50764 26580
rect 50712 26537 50721 26571
rect 50721 26537 50755 26571
rect 50755 26537 50764 26571
rect 50712 26528 50764 26537
rect 53380 26528 53432 26580
rect 55772 26528 55824 26580
rect 29552 26460 29604 26512
rect 33692 26435 33744 26444
rect 24400 26367 24452 26376
rect 24400 26333 24409 26367
rect 24409 26333 24443 26367
rect 24443 26333 24452 26367
rect 24400 26324 24452 26333
rect 27896 26367 27948 26376
rect 24124 26256 24176 26308
rect 27896 26333 27905 26367
rect 27905 26333 27939 26367
rect 27939 26333 27948 26367
rect 27896 26324 27948 26333
rect 30564 26367 30616 26376
rect 30564 26333 30573 26367
rect 30573 26333 30607 26367
rect 30607 26333 30616 26367
rect 30564 26324 30616 26333
rect 30748 26367 30800 26376
rect 30748 26333 30757 26367
rect 30757 26333 30791 26367
rect 30791 26333 30800 26367
rect 30748 26324 30800 26333
rect 33692 26401 33701 26435
rect 33701 26401 33735 26435
rect 33735 26401 33744 26435
rect 43168 26460 43220 26512
rect 33692 26392 33744 26401
rect 33140 26324 33192 26376
rect 33600 26324 33652 26376
rect 40500 26392 40552 26444
rect 49976 26392 50028 26444
rect 50896 26392 50948 26444
rect 37464 26324 37516 26376
rect 38108 26324 38160 26376
rect 38752 26324 38804 26376
rect 40224 26324 40276 26376
rect 41144 26367 41196 26376
rect 41144 26333 41153 26367
rect 41153 26333 41187 26367
rect 41187 26333 41196 26367
rect 41144 26324 41196 26333
rect 50068 26324 50120 26376
rect 51356 26367 51408 26376
rect 51356 26333 51365 26367
rect 51365 26333 51399 26367
rect 51399 26333 51408 26367
rect 51356 26324 51408 26333
rect 52828 26367 52880 26376
rect 52828 26333 52837 26367
rect 52837 26333 52871 26367
rect 52871 26333 52880 26367
rect 52828 26324 52880 26333
rect 55956 26367 56008 26376
rect 55956 26333 55965 26367
rect 55965 26333 55999 26367
rect 55999 26333 56008 26367
rect 55956 26324 56008 26333
rect 56600 26324 56652 26376
rect 37280 26256 37332 26308
rect 45100 26256 45152 26308
rect 52276 26256 52328 26308
rect 52460 26256 52512 26308
rect 53656 26256 53708 26308
rect 20628 26188 20680 26240
rect 21088 26188 21140 26240
rect 21916 26188 21968 26240
rect 24032 26188 24084 26240
rect 28080 26188 28132 26240
rect 39948 26188 40000 26240
rect 53196 26188 53248 26240
rect 19574 26086 19626 26138
rect 19638 26086 19690 26138
rect 19702 26086 19754 26138
rect 19766 26086 19818 26138
rect 19830 26086 19882 26138
rect 50294 26086 50346 26138
rect 50358 26086 50410 26138
rect 50422 26086 50474 26138
rect 50486 26086 50538 26138
rect 50550 26086 50602 26138
rect 2780 26027 2832 26036
rect 2780 25993 2789 26027
rect 2789 25993 2823 26027
rect 2823 25993 2832 26027
rect 2780 25984 2832 25993
rect 4068 25984 4120 26036
rect 6276 25984 6328 26036
rect 9956 26027 10008 26036
rect 9956 25993 9965 26027
rect 9965 25993 9999 26027
rect 9999 25993 10008 26027
rect 9956 25984 10008 25993
rect 10600 25984 10652 26036
rect 10692 25984 10744 26036
rect 3148 25891 3200 25900
rect 3148 25857 3157 25891
rect 3157 25857 3191 25891
rect 3191 25857 3200 25891
rect 3148 25848 3200 25857
rect 6920 25848 6972 25900
rect 3148 25712 3200 25764
rect 3976 25755 4028 25764
rect 3976 25721 3985 25755
rect 3985 25721 4019 25755
rect 4019 25721 4028 25755
rect 3976 25712 4028 25721
rect 6644 25712 6696 25764
rect 9404 25891 9456 25900
rect 9404 25857 9413 25891
rect 9413 25857 9447 25891
rect 9447 25857 9456 25891
rect 9404 25848 9456 25857
rect 9772 25848 9824 25900
rect 11244 25916 11296 25968
rect 12992 25916 13044 25968
rect 14464 25984 14516 26036
rect 17776 26027 17828 26036
rect 17776 25993 17785 26027
rect 17785 25993 17819 26027
rect 17819 25993 17828 26027
rect 17776 25984 17828 25993
rect 18236 25984 18288 26036
rect 19064 25984 19116 26036
rect 20628 25984 20680 26036
rect 28172 25984 28224 26036
rect 38752 26027 38804 26036
rect 38752 25993 38761 26027
rect 38761 25993 38795 26027
rect 38795 25993 38804 26027
rect 38752 25984 38804 25993
rect 44180 25984 44232 26036
rect 47952 26027 48004 26036
rect 47952 25993 47961 26027
rect 47961 25993 47995 26027
rect 47995 25993 48004 26027
rect 47952 25984 48004 25993
rect 10232 25891 10284 25900
rect 10232 25857 10241 25891
rect 10241 25857 10275 25891
rect 10275 25857 10284 25891
rect 10232 25848 10284 25857
rect 9680 25780 9732 25832
rect 10324 25780 10376 25832
rect 10600 25848 10652 25900
rect 10140 25712 10192 25764
rect 3424 25644 3476 25696
rect 9404 25644 9456 25696
rect 11060 25644 11112 25696
rect 11796 25891 11848 25900
rect 11796 25857 11805 25891
rect 11805 25857 11839 25891
rect 11839 25857 11848 25891
rect 13268 25891 13320 25900
rect 11796 25848 11848 25857
rect 13268 25857 13277 25891
rect 13277 25857 13311 25891
rect 13311 25857 13320 25891
rect 13268 25848 13320 25857
rect 13636 25891 13688 25900
rect 13176 25780 13228 25832
rect 13636 25857 13645 25891
rect 13645 25857 13679 25891
rect 13679 25857 13688 25891
rect 13636 25848 13688 25857
rect 15200 25916 15252 25968
rect 18144 25916 18196 25968
rect 21088 25959 21140 25968
rect 21088 25925 21097 25959
rect 21097 25925 21131 25959
rect 21131 25925 21140 25959
rect 21088 25916 21140 25925
rect 21732 25916 21784 25968
rect 14740 25848 14792 25900
rect 17224 25891 17276 25900
rect 17224 25857 17233 25891
rect 17233 25857 17267 25891
rect 17267 25857 17276 25891
rect 17224 25848 17276 25857
rect 17408 25891 17460 25900
rect 17408 25857 17417 25891
rect 17417 25857 17451 25891
rect 17451 25857 17460 25891
rect 17408 25848 17460 25857
rect 17684 25848 17736 25900
rect 13728 25780 13780 25832
rect 22284 25891 22336 25900
rect 22284 25857 22293 25891
rect 22293 25857 22327 25891
rect 22327 25857 22336 25891
rect 24032 25891 24084 25900
rect 22284 25848 22336 25857
rect 24032 25857 24041 25891
rect 24041 25857 24075 25891
rect 24075 25857 24084 25891
rect 24032 25848 24084 25857
rect 22928 25780 22980 25832
rect 24492 25891 24544 25900
rect 24492 25857 24506 25891
rect 24506 25857 24540 25891
rect 24540 25857 24544 25891
rect 24768 25916 24820 25968
rect 49332 25984 49384 26036
rect 50068 26027 50120 26036
rect 50068 25993 50077 26027
rect 50077 25993 50111 26027
rect 50111 25993 50120 26027
rect 50068 25984 50120 25993
rect 52828 25984 52880 26036
rect 53196 26027 53248 26036
rect 53196 25993 53205 26027
rect 53205 25993 53239 26027
rect 53239 25993 53248 26027
rect 53196 25984 53248 25993
rect 24492 25848 24544 25857
rect 24952 25848 25004 25900
rect 28080 25891 28132 25900
rect 28080 25857 28089 25891
rect 28089 25857 28123 25891
rect 28123 25857 28132 25891
rect 28080 25848 28132 25857
rect 24584 25780 24636 25832
rect 28264 25823 28316 25832
rect 28264 25789 28273 25823
rect 28273 25789 28307 25823
rect 28307 25789 28316 25823
rect 28264 25780 28316 25789
rect 54024 26027 54076 26036
rect 54024 25993 54033 26027
rect 54033 25993 54067 26027
rect 54067 25993 54076 26027
rect 54024 25984 54076 25993
rect 55956 25984 56008 26036
rect 53656 25959 53708 25968
rect 30748 25848 30800 25900
rect 37464 25891 37516 25900
rect 37464 25857 37473 25891
rect 37473 25857 37507 25891
rect 37507 25857 37516 25891
rect 37464 25848 37516 25857
rect 43812 25848 43864 25900
rect 46848 25891 46900 25900
rect 46848 25857 46857 25891
rect 46857 25857 46891 25891
rect 46891 25857 46900 25891
rect 46848 25848 46900 25857
rect 47032 25891 47084 25900
rect 47032 25857 47041 25891
rect 47041 25857 47075 25891
rect 47075 25857 47084 25891
rect 47032 25848 47084 25857
rect 47584 25891 47636 25900
rect 47584 25857 47593 25891
rect 47593 25857 47627 25891
rect 47627 25857 47636 25891
rect 47584 25848 47636 25857
rect 53656 25925 53665 25959
rect 53665 25925 53699 25959
rect 53699 25925 53708 25959
rect 53656 25916 53708 25925
rect 37280 25780 37332 25832
rect 38016 25780 38068 25832
rect 43720 25823 43772 25832
rect 43720 25789 43729 25823
rect 43729 25789 43763 25823
rect 43763 25789 43772 25823
rect 43720 25780 43772 25789
rect 49240 25823 49292 25832
rect 49240 25789 49249 25823
rect 49249 25789 49283 25823
rect 49283 25789 49292 25823
rect 50160 25891 50212 25900
rect 50160 25857 50169 25891
rect 50169 25857 50203 25891
rect 50203 25857 50212 25891
rect 50160 25848 50212 25857
rect 52368 25848 52420 25900
rect 49240 25780 49292 25789
rect 52276 25780 52328 25832
rect 53104 25848 53156 25900
rect 55956 25848 56008 25900
rect 52920 25780 52972 25832
rect 55772 25823 55824 25832
rect 55772 25789 55781 25823
rect 55781 25789 55815 25823
rect 55815 25789 55824 25823
rect 55772 25780 55824 25789
rect 13084 25712 13136 25764
rect 14096 25712 14148 25764
rect 20904 25712 20956 25764
rect 21548 25712 21600 25764
rect 34520 25712 34572 25764
rect 37188 25712 37240 25764
rect 18052 25644 18104 25696
rect 23940 25644 23992 25696
rect 40132 25644 40184 25696
rect 53196 25644 53248 25696
rect 4214 25542 4266 25594
rect 4278 25542 4330 25594
rect 4342 25542 4394 25594
rect 4406 25542 4458 25594
rect 4470 25542 4522 25594
rect 34934 25542 34986 25594
rect 34998 25542 35050 25594
rect 35062 25542 35114 25594
rect 35126 25542 35178 25594
rect 35190 25542 35242 25594
rect 6644 25440 6696 25492
rect 9864 25440 9916 25492
rect 10324 25483 10376 25492
rect 10324 25449 10333 25483
rect 10333 25449 10367 25483
rect 10367 25449 10376 25483
rect 10324 25440 10376 25449
rect 20720 25440 20772 25492
rect 21732 25483 21784 25492
rect 21732 25449 21741 25483
rect 21741 25449 21775 25483
rect 21775 25449 21784 25483
rect 21732 25440 21784 25449
rect 22192 25440 22244 25492
rect 43812 25483 43864 25492
rect 3056 25372 3108 25424
rect 3516 25372 3568 25424
rect 14556 25372 14608 25424
rect 2504 25236 2556 25288
rect 3976 25304 4028 25356
rect 4068 25304 4120 25356
rect 3148 25236 3200 25288
rect 3792 25279 3844 25288
rect 3792 25245 3801 25279
rect 3801 25245 3835 25279
rect 3835 25245 3844 25279
rect 3792 25236 3844 25245
rect 1860 25211 1912 25220
rect 1860 25177 1869 25211
rect 1869 25177 1903 25211
rect 1903 25177 1912 25211
rect 1860 25168 1912 25177
rect 2596 25168 2648 25220
rect 4252 25236 4304 25288
rect 9404 25304 9456 25356
rect 6276 25168 6328 25220
rect 12440 25236 12492 25288
rect 12992 25279 13044 25288
rect 12992 25245 13001 25279
rect 13001 25245 13035 25279
rect 13035 25245 13044 25279
rect 12992 25236 13044 25245
rect 13636 25304 13688 25356
rect 14004 25304 14056 25356
rect 6828 25168 6880 25220
rect 10048 25168 10100 25220
rect 10692 25168 10744 25220
rect 13176 25211 13228 25220
rect 13176 25177 13185 25211
rect 13185 25177 13219 25211
rect 13219 25177 13228 25211
rect 13176 25168 13228 25177
rect 7012 25100 7064 25152
rect 12716 25100 12768 25152
rect 14924 25236 14976 25288
rect 16764 25236 16816 25288
rect 17132 25236 17184 25288
rect 20168 25372 20220 25424
rect 21548 25372 21600 25424
rect 24492 25372 24544 25424
rect 17408 25304 17460 25356
rect 17960 25279 18012 25288
rect 17960 25245 17970 25279
rect 17970 25245 18004 25279
rect 18004 25245 18012 25279
rect 18236 25279 18288 25288
rect 17960 25236 18012 25245
rect 18236 25245 18245 25279
rect 18245 25245 18279 25279
rect 18279 25245 18288 25279
rect 18236 25236 18288 25245
rect 18328 25279 18380 25288
rect 18328 25245 18342 25279
rect 18342 25245 18376 25279
rect 18376 25245 18380 25279
rect 18328 25236 18380 25245
rect 20628 25236 20680 25288
rect 23388 25236 23440 25288
rect 23572 25279 23624 25288
rect 23572 25245 23581 25279
rect 23581 25245 23615 25279
rect 23615 25245 23624 25279
rect 23572 25236 23624 25245
rect 23756 25279 23808 25288
rect 23756 25245 23765 25279
rect 23765 25245 23799 25279
rect 23799 25245 23808 25279
rect 23756 25236 23808 25245
rect 24584 25279 24636 25288
rect 24584 25245 24591 25279
rect 24591 25245 24636 25279
rect 24584 25236 24636 25245
rect 27712 25304 27764 25356
rect 28264 25304 28316 25356
rect 30656 25415 30708 25424
rect 30656 25381 30665 25415
rect 30665 25381 30699 25415
rect 30699 25381 30708 25415
rect 30656 25372 30708 25381
rect 27620 25279 27672 25288
rect 27620 25245 27629 25279
rect 27629 25245 27663 25279
rect 27663 25245 27672 25279
rect 27620 25236 27672 25245
rect 28172 25236 28224 25288
rect 31300 25347 31352 25356
rect 31300 25313 31309 25347
rect 31309 25313 31343 25347
rect 31343 25313 31352 25347
rect 31300 25304 31352 25313
rect 33692 25372 33744 25424
rect 28724 25279 28776 25288
rect 28724 25245 28733 25279
rect 28733 25245 28767 25279
rect 28767 25245 28776 25279
rect 28724 25236 28776 25245
rect 31392 25279 31444 25288
rect 31392 25245 31401 25279
rect 31401 25245 31435 25279
rect 31435 25245 31444 25279
rect 31392 25236 31444 25245
rect 14096 25100 14148 25152
rect 14464 25211 14516 25220
rect 14464 25177 14473 25211
rect 14473 25177 14507 25211
rect 14507 25177 14516 25211
rect 16856 25211 16908 25220
rect 14464 25168 14516 25177
rect 16856 25177 16865 25211
rect 16865 25177 16899 25211
rect 16899 25177 16908 25211
rect 16856 25168 16908 25177
rect 17316 25168 17368 25220
rect 18144 25211 18196 25220
rect 18144 25177 18153 25211
rect 18153 25177 18187 25211
rect 18187 25177 18196 25211
rect 18144 25168 18196 25177
rect 18696 25168 18748 25220
rect 21732 25168 21784 25220
rect 24768 25211 24820 25220
rect 24768 25177 24777 25211
rect 24777 25177 24811 25211
rect 24811 25177 24820 25211
rect 34612 25372 34664 25424
rect 37464 25372 37516 25424
rect 38016 25415 38068 25424
rect 38016 25381 38025 25415
rect 38025 25381 38059 25415
rect 38059 25381 38068 25415
rect 38016 25372 38068 25381
rect 38108 25415 38160 25424
rect 38108 25381 38117 25415
rect 38117 25381 38151 25415
rect 38151 25381 38160 25415
rect 43812 25449 43821 25483
rect 43821 25449 43855 25483
rect 43855 25449 43864 25483
rect 43812 25440 43864 25449
rect 47584 25440 47636 25492
rect 50160 25483 50212 25492
rect 50160 25449 50169 25483
rect 50169 25449 50203 25483
rect 50203 25449 50212 25483
rect 50160 25440 50212 25449
rect 52828 25483 52880 25492
rect 52828 25449 52837 25483
rect 52837 25449 52871 25483
rect 52871 25449 52880 25483
rect 52828 25440 52880 25449
rect 55956 25483 56008 25492
rect 38108 25372 38160 25381
rect 52552 25372 52604 25424
rect 24768 25168 24820 25177
rect 14740 25143 14792 25152
rect 14740 25109 14749 25143
rect 14749 25109 14783 25143
rect 14783 25109 14792 25143
rect 14740 25100 14792 25109
rect 18236 25100 18288 25152
rect 18512 25100 18564 25152
rect 21364 25100 21416 25152
rect 34704 25236 34756 25288
rect 40132 25279 40184 25288
rect 40132 25245 40141 25279
rect 40141 25245 40175 25279
rect 40175 25245 40184 25279
rect 40132 25236 40184 25245
rect 40960 25279 41012 25288
rect 40960 25245 40969 25279
rect 40969 25245 41003 25279
rect 41003 25245 41012 25279
rect 40960 25236 41012 25245
rect 49240 25304 49292 25356
rect 52368 25304 52420 25356
rect 52920 25347 52972 25356
rect 52920 25313 52929 25347
rect 52929 25313 52963 25347
rect 52963 25313 52972 25347
rect 52920 25304 52972 25313
rect 55588 25347 55640 25356
rect 55588 25313 55597 25347
rect 55597 25313 55631 25347
rect 55631 25313 55640 25347
rect 55956 25449 55965 25483
rect 55965 25449 55999 25483
rect 55999 25449 56008 25483
rect 55956 25440 56008 25449
rect 55588 25304 55640 25313
rect 55864 25304 55916 25356
rect 41880 25236 41932 25288
rect 42800 25279 42852 25288
rect 42800 25245 42809 25279
rect 42809 25245 42843 25279
rect 42843 25245 42852 25279
rect 42800 25236 42852 25245
rect 43720 25279 43772 25288
rect 43720 25245 43729 25279
rect 43729 25245 43763 25279
rect 43763 25245 43772 25279
rect 43720 25236 43772 25245
rect 45744 25236 45796 25288
rect 45928 25236 45980 25288
rect 46112 25279 46164 25288
rect 46112 25245 46121 25279
rect 46121 25245 46155 25279
rect 46155 25245 46164 25279
rect 46112 25236 46164 25245
rect 46296 25236 46348 25288
rect 46848 25236 46900 25288
rect 50160 25279 50212 25288
rect 50160 25245 50169 25279
rect 50169 25245 50203 25279
rect 50203 25245 50212 25279
rect 50160 25236 50212 25245
rect 53196 25279 53248 25288
rect 53196 25245 53205 25279
rect 53205 25245 53239 25279
rect 53239 25245 53248 25279
rect 53196 25236 53248 25245
rect 53656 25236 53708 25288
rect 55404 25236 55456 25288
rect 57888 25279 57940 25288
rect 37188 25168 37240 25220
rect 40316 25211 40368 25220
rect 40316 25177 40325 25211
rect 40325 25177 40359 25211
rect 40359 25177 40368 25211
rect 40316 25168 40368 25177
rect 41604 25168 41656 25220
rect 57888 25245 57897 25279
rect 57897 25245 57931 25279
rect 57931 25245 57940 25279
rect 57888 25236 57940 25245
rect 26608 25100 26660 25152
rect 34060 25143 34112 25152
rect 34060 25109 34069 25143
rect 34069 25109 34103 25143
rect 34103 25109 34112 25143
rect 34060 25100 34112 25109
rect 44180 25143 44232 25152
rect 44180 25109 44189 25143
rect 44189 25109 44223 25143
rect 44223 25109 44232 25143
rect 44180 25100 44232 25109
rect 52276 25100 52328 25152
rect 55680 25100 55732 25152
rect 58072 25143 58124 25152
rect 58072 25109 58081 25143
rect 58081 25109 58115 25143
rect 58115 25109 58124 25143
rect 58072 25100 58124 25109
rect 19574 24998 19626 25050
rect 19638 24998 19690 25050
rect 19702 24998 19754 25050
rect 19766 24998 19818 25050
rect 19830 24998 19882 25050
rect 50294 24998 50346 25050
rect 50358 24998 50410 25050
rect 50422 24998 50474 25050
rect 50486 24998 50538 25050
rect 50550 24998 50602 25050
rect 1860 24896 1912 24948
rect 3056 24896 3108 24948
rect 3884 24896 3936 24948
rect 8300 24896 8352 24948
rect 8484 24896 8536 24948
rect 15660 24896 15712 24948
rect 17960 24896 18012 24948
rect 8208 24871 8260 24880
rect 8208 24837 8217 24871
rect 8217 24837 8251 24871
rect 8251 24837 8260 24871
rect 8208 24828 8260 24837
rect 11980 24828 12032 24880
rect 16488 24828 16540 24880
rect 17224 24828 17276 24880
rect 20168 24828 20220 24880
rect 2504 24803 2556 24812
rect 2504 24769 2513 24803
rect 2513 24769 2547 24803
rect 2547 24769 2556 24803
rect 2504 24760 2556 24769
rect 2596 24760 2648 24812
rect 3148 24803 3200 24812
rect 3148 24769 3157 24803
rect 3157 24769 3191 24803
rect 3191 24769 3200 24803
rect 3148 24760 3200 24769
rect 3424 24803 3476 24812
rect 3424 24769 3433 24803
rect 3433 24769 3467 24803
rect 3467 24769 3476 24803
rect 3424 24760 3476 24769
rect 3792 24692 3844 24744
rect 7012 24803 7064 24812
rect 7012 24769 7021 24803
rect 7021 24769 7055 24803
rect 7055 24769 7064 24803
rect 7196 24803 7248 24812
rect 7012 24760 7064 24769
rect 7196 24769 7205 24803
rect 7205 24769 7239 24803
rect 7239 24769 7248 24803
rect 7196 24760 7248 24769
rect 7288 24803 7340 24812
rect 7288 24769 7297 24803
rect 7297 24769 7331 24803
rect 7331 24769 7340 24803
rect 7472 24803 7524 24812
rect 7288 24760 7340 24769
rect 7472 24769 7481 24803
rect 7481 24769 7515 24803
rect 7515 24769 7524 24803
rect 7472 24760 7524 24769
rect 8024 24803 8076 24812
rect 8024 24769 8033 24803
rect 8033 24769 8067 24803
rect 8067 24769 8076 24803
rect 8024 24760 8076 24769
rect 8668 24760 8720 24812
rect 9680 24803 9732 24812
rect 9680 24769 9689 24803
rect 9689 24769 9723 24803
rect 9723 24769 9732 24803
rect 9680 24760 9732 24769
rect 10048 24760 10100 24812
rect 13544 24760 13596 24812
rect 8392 24692 8444 24744
rect 13360 24692 13412 24744
rect 15200 24760 15252 24812
rect 17040 24760 17092 24812
rect 20076 24803 20128 24812
rect 20076 24769 20085 24803
rect 20085 24769 20119 24803
rect 20119 24769 20128 24803
rect 20076 24760 20128 24769
rect 21272 24828 21324 24880
rect 21364 24828 21416 24880
rect 27620 24896 27672 24948
rect 31392 24896 31444 24948
rect 34520 24896 34572 24948
rect 34704 24896 34756 24948
rect 40960 24896 41012 24948
rect 50160 24896 50212 24948
rect 53932 24896 53984 24948
rect 57980 24939 58032 24948
rect 34060 24828 34112 24880
rect 23480 24803 23532 24812
rect 17408 24692 17460 24744
rect 18328 24692 18380 24744
rect 19340 24692 19392 24744
rect 20812 24692 20864 24744
rect 23480 24769 23489 24803
rect 23489 24769 23523 24803
rect 23523 24769 23532 24803
rect 23480 24760 23532 24769
rect 23756 24760 23808 24812
rect 24400 24803 24452 24812
rect 24400 24769 24409 24803
rect 24409 24769 24443 24803
rect 24443 24769 24452 24803
rect 24400 24760 24452 24769
rect 25136 24760 25188 24812
rect 26240 24760 26292 24812
rect 27712 24760 27764 24812
rect 28080 24803 28132 24812
rect 28080 24769 28089 24803
rect 28089 24769 28123 24803
rect 28123 24769 28132 24803
rect 28080 24760 28132 24769
rect 25320 24735 25372 24744
rect 25320 24701 25329 24735
rect 25329 24701 25363 24735
rect 25363 24701 25372 24735
rect 25320 24692 25372 24701
rect 25412 24692 25464 24744
rect 10784 24624 10836 24676
rect 14188 24624 14240 24676
rect 16764 24624 16816 24676
rect 17132 24624 17184 24676
rect 17684 24624 17736 24676
rect 18512 24624 18564 24676
rect 20260 24667 20312 24676
rect 20260 24633 20269 24667
rect 20269 24633 20303 24667
rect 20303 24633 20312 24667
rect 20260 24624 20312 24633
rect 23664 24624 23716 24676
rect 26240 24624 26292 24676
rect 26792 24624 26844 24676
rect 33784 24760 33836 24812
rect 33968 24803 34020 24812
rect 33968 24769 33977 24803
rect 33977 24769 34011 24803
rect 34011 24769 34020 24803
rect 33968 24760 34020 24769
rect 36544 24760 36596 24812
rect 39120 24760 39172 24812
rect 40132 24760 40184 24812
rect 31116 24735 31168 24744
rect 31116 24701 31125 24735
rect 31125 24701 31159 24735
rect 31159 24701 31168 24735
rect 31116 24692 31168 24701
rect 38568 24692 38620 24744
rect 40316 24760 40368 24812
rect 41604 24803 41656 24812
rect 41604 24769 41613 24803
rect 41613 24769 41647 24803
rect 41647 24769 41656 24803
rect 41604 24760 41656 24769
rect 41880 24760 41932 24812
rect 44180 24760 44232 24812
rect 44548 24803 44600 24812
rect 44548 24769 44557 24803
rect 44557 24769 44591 24803
rect 44591 24769 44600 24803
rect 44548 24760 44600 24769
rect 45376 24760 45428 24812
rect 45744 24803 45796 24812
rect 42800 24692 42852 24744
rect 45100 24735 45152 24744
rect 45100 24701 45109 24735
rect 45109 24701 45143 24735
rect 45143 24701 45152 24735
rect 45100 24692 45152 24701
rect 45744 24769 45753 24803
rect 45753 24769 45787 24803
rect 45787 24769 45796 24803
rect 45744 24760 45796 24769
rect 45836 24803 45888 24812
rect 45836 24769 45845 24803
rect 45845 24769 45879 24803
rect 45879 24769 45888 24803
rect 47032 24828 47084 24880
rect 52920 24828 52972 24880
rect 55588 24828 55640 24880
rect 57980 24905 57989 24939
rect 57989 24905 58023 24939
rect 58023 24905 58032 24939
rect 57980 24896 58032 24905
rect 45836 24760 45888 24769
rect 46296 24760 46348 24812
rect 45652 24692 45704 24744
rect 46112 24735 46164 24744
rect 46112 24701 46121 24735
rect 46121 24701 46155 24735
rect 46155 24701 46164 24735
rect 46112 24692 46164 24701
rect 51080 24803 51132 24812
rect 51080 24769 51089 24803
rect 51089 24769 51123 24803
rect 51123 24769 51132 24803
rect 51080 24760 51132 24769
rect 53196 24760 53248 24812
rect 55404 24803 55456 24812
rect 55404 24769 55413 24803
rect 55413 24769 55447 24803
rect 55447 24769 55456 24803
rect 55404 24760 55456 24769
rect 55496 24803 55548 24812
rect 55496 24769 55505 24803
rect 55505 24769 55539 24803
rect 55539 24769 55548 24803
rect 55496 24760 55548 24769
rect 55680 24692 55732 24744
rect 55864 24803 55916 24812
rect 55864 24769 55873 24803
rect 55873 24769 55907 24803
rect 55907 24769 55916 24803
rect 55864 24760 55916 24769
rect 56968 24803 57020 24812
rect 56968 24769 56977 24803
rect 56977 24769 57011 24803
rect 57011 24769 57020 24803
rect 56968 24760 57020 24769
rect 57060 24692 57112 24744
rect 57244 24760 57296 24812
rect 57888 24803 57940 24812
rect 57888 24769 57897 24803
rect 57897 24769 57931 24803
rect 57931 24769 57940 24803
rect 57888 24760 57940 24769
rect 56968 24624 57020 24676
rect 3608 24599 3660 24608
rect 3608 24565 3617 24599
rect 3617 24565 3651 24599
rect 3651 24565 3660 24599
rect 3608 24556 3660 24565
rect 7196 24556 7248 24608
rect 8668 24556 8720 24608
rect 9680 24556 9732 24608
rect 14096 24599 14148 24608
rect 14096 24565 14105 24599
rect 14105 24565 14139 24599
rect 14139 24565 14148 24599
rect 14096 24556 14148 24565
rect 15016 24556 15068 24608
rect 16488 24556 16540 24608
rect 20076 24556 20128 24608
rect 20536 24556 20588 24608
rect 28540 24599 28592 24608
rect 28540 24565 28549 24599
rect 28549 24565 28583 24599
rect 28583 24565 28592 24599
rect 28540 24556 28592 24565
rect 33232 24599 33284 24608
rect 33232 24565 33241 24599
rect 33241 24565 33275 24599
rect 33275 24565 33284 24599
rect 33232 24556 33284 24565
rect 33876 24556 33928 24608
rect 37372 24556 37424 24608
rect 37740 24599 37792 24608
rect 37740 24565 37749 24599
rect 37749 24565 37783 24599
rect 37783 24565 37792 24599
rect 37740 24556 37792 24565
rect 39948 24556 40000 24608
rect 40960 24556 41012 24608
rect 45836 24556 45888 24608
rect 49516 24599 49568 24608
rect 49516 24565 49525 24599
rect 49525 24565 49559 24599
rect 49559 24565 49568 24599
rect 49516 24556 49568 24565
rect 57152 24556 57204 24608
rect 4214 24454 4266 24506
rect 4278 24454 4330 24506
rect 4342 24454 4394 24506
rect 4406 24454 4458 24506
rect 4470 24454 4522 24506
rect 34934 24454 34986 24506
rect 34998 24454 35050 24506
rect 35062 24454 35114 24506
rect 35126 24454 35178 24506
rect 35190 24454 35242 24506
rect 3884 24395 3936 24404
rect 3884 24361 3893 24395
rect 3893 24361 3927 24395
rect 3927 24361 3936 24395
rect 3884 24352 3936 24361
rect 8208 24352 8260 24404
rect 8392 24352 8444 24404
rect 10876 24352 10928 24404
rect 12808 24352 12860 24404
rect 17040 24352 17092 24404
rect 17960 24395 18012 24404
rect 17960 24361 17969 24395
rect 17969 24361 18003 24395
rect 18003 24361 18012 24395
rect 17960 24352 18012 24361
rect 7656 24284 7708 24336
rect 13360 24284 13412 24336
rect 14740 24327 14792 24336
rect 14740 24293 14749 24327
rect 14749 24293 14783 24327
rect 14783 24293 14792 24327
rect 14740 24284 14792 24293
rect 6920 24148 6972 24200
rect 8392 24148 8444 24200
rect 9220 24148 9272 24200
rect 10324 24148 10376 24200
rect 9312 24080 9364 24132
rect 9772 24080 9824 24132
rect 12992 24148 13044 24200
rect 14188 24191 14240 24200
rect 14188 24157 14198 24191
rect 14198 24157 14232 24191
rect 14232 24157 14240 24191
rect 14648 24216 14700 24268
rect 14464 24191 14516 24200
rect 14188 24148 14240 24157
rect 14464 24157 14473 24191
rect 14473 24157 14507 24191
rect 14507 24157 14516 24191
rect 14464 24148 14516 24157
rect 14556 24191 14608 24200
rect 16488 24216 16540 24268
rect 14556 24157 14570 24191
rect 14570 24157 14604 24191
rect 14604 24157 14608 24191
rect 14556 24148 14608 24157
rect 16580 24191 16632 24200
rect 10784 24080 10836 24132
rect 13544 24123 13596 24132
rect 13544 24089 13553 24123
rect 13553 24089 13587 24123
rect 13587 24089 13596 24123
rect 13544 24080 13596 24089
rect 16580 24157 16589 24191
rect 16589 24157 16623 24191
rect 16623 24157 16632 24191
rect 16580 24148 16632 24157
rect 16764 24148 16816 24200
rect 17224 24148 17276 24200
rect 17408 24191 17460 24200
rect 17408 24157 17418 24191
rect 17418 24157 17452 24191
rect 17452 24157 17460 24191
rect 17408 24148 17460 24157
rect 16488 24123 16540 24132
rect 16488 24089 16497 24123
rect 16497 24089 16531 24123
rect 16531 24089 16540 24123
rect 19064 24216 19116 24268
rect 17776 24191 17828 24200
rect 17776 24157 17790 24191
rect 17790 24157 17824 24191
rect 17824 24157 17828 24191
rect 17776 24148 17828 24157
rect 18512 24148 18564 24200
rect 20720 24352 20772 24404
rect 21456 24395 21508 24404
rect 21456 24361 21465 24395
rect 21465 24361 21499 24395
rect 21499 24361 21508 24395
rect 21456 24352 21508 24361
rect 20076 24191 20128 24200
rect 20076 24157 20085 24191
rect 20085 24157 20119 24191
rect 20119 24157 20128 24191
rect 20076 24148 20128 24157
rect 20168 24191 20220 24200
rect 20168 24157 20177 24191
rect 20177 24157 20211 24191
rect 20211 24157 20220 24191
rect 24952 24352 25004 24404
rect 25136 24395 25188 24404
rect 25136 24361 25145 24395
rect 25145 24361 25179 24395
rect 25179 24361 25188 24395
rect 25136 24352 25188 24361
rect 25596 24352 25648 24404
rect 27712 24395 27764 24404
rect 23388 24284 23440 24336
rect 27712 24361 27721 24395
rect 27721 24361 27755 24395
rect 27755 24361 27764 24395
rect 27712 24352 27764 24361
rect 27804 24352 27856 24404
rect 28724 24352 28776 24404
rect 31116 24395 31168 24404
rect 31116 24361 31125 24395
rect 31125 24361 31159 24395
rect 31159 24361 31168 24395
rect 31116 24352 31168 24361
rect 33968 24395 34020 24404
rect 33968 24361 33977 24395
rect 33977 24361 34011 24395
rect 34011 24361 34020 24395
rect 33968 24352 34020 24361
rect 20168 24148 20220 24157
rect 20904 24148 20956 24200
rect 23664 24216 23716 24268
rect 24768 24216 24820 24268
rect 21456 24148 21508 24200
rect 23572 24148 23624 24200
rect 24492 24191 24544 24200
rect 24492 24157 24501 24191
rect 24501 24157 24535 24191
rect 24535 24157 24544 24191
rect 24492 24148 24544 24157
rect 24584 24191 24636 24200
rect 24584 24157 24594 24191
rect 24594 24157 24628 24191
rect 24628 24157 24636 24191
rect 24584 24148 24636 24157
rect 25044 24148 25096 24200
rect 16488 24080 16540 24089
rect 13268 24012 13320 24064
rect 13820 24012 13872 24064
rect 14096 24012 14148 24064
rect 14188 24012 14240 24064
rect 19984 24123 20036 24132
rect 17868 24012 17920 24064
rect 19984 24089 19993 24123
rect 19993 24089 20027 24123
rect 20027 24089 20036 24123
rect 19984 24080 20036 24089
rect 20444 24080 20496 24132
rect 21180 24123 21232 24132
rect 21180 24089 21189 24123
rect 21189 24089 21223 24123
rect 21223 24089 21232 24123
rect 21180 24080 21232 24089
rect 23020 24080 23072 24132
rect 23940 24080 23992 24132
rect 28540 24191 28592 24200
rect 28540 24157 28549 24191
rect 28549 24157 28583 24191
rect 28583 24157 28592 24191
rect 28540 24148 28592 24157
rect 28816 24191 28868 24200
rect 28816 24157 28825 24191
rect 28825 24157 28859 24191
rect 28859 24157 28868 24191
rect 28816 24148 28868 24157
rect 33876 24191 33928 24200
rect 33876 24157 33885 24191
rect 33885 24157 33919 24191
rect 33919 24157 33928 24191
rect 33876 24148 33928 24157
rect 38568 24395 38620 24404
rect 38568 24361 38577 24395
rect 38577 24361 38611 24395
rect 38611 24361 38620 24395
rect 38568 24352 38620 24361
rect 39120 24395 39172 24404
rect 39120 24361 39129 24395
rect 39129 24361 39163 24395
rect 39163 24361 39172 24395
rect 39120 24352 39172 24361
rect 40224 24352 40276 24404
rect 44548 24352 44600 24404
rect 45652 24395 45704 24404
rect 45652 24361 45661 24395
rect 45661 24361 45695 24395
rect 45695 24361 45704 24395
rect 45652 24352 45704 24361
rect 55496 24352 55548 24404
rect 37648 24327 37700 24336
rect 37648 24293 37657 24327
rect 37657 24293 37691 24327
rect 37691 24293 37700 24327
rect 37648 24284 37700 24293
rect 43812 24284 43864 24336
rect 40592 24216 40644 24268
rect 38108 24191 38160 24200
rect 38108 24157 38117 24191
rect 38117 24157 38151 24191
rect 38151 24157 38160 24191
rect 38108 24148 38160 24157
rect 41052 24191 41104 24200
rect 20260 24012 20312 24064
rect 20996 24012 21048 24064
rect 21364 24012 21416 24064
rect 22744 24012 22796 24064
rect 24584 24012 24636 24064
rect 25964 24012 26016 24064
rect 29460 24012 29512 24064
rect 29644 24012 29696 24064
rect 31300 24055 31352 24064
rect 31300 24021 31309 24055
rect 31309 24021 31343 24055
rect 31343 24021 31352 24055
rect 31300 24012 31352 24021
rect 33784 24012 33836 24064
rect 34336 24012 34388 24064
rect 37740 24080 37792 24132
rect 41052 24157 41061 24191
rect 41061 24157 41095 24191
rect 41095 24157 41104 24191
rect 41052 24148 41104 24157
rect 45100 24216 45152 24268
rect 43812 24148 43864 24200
rect 44180 24148 44232 24200
rect 49240 24216 49292 24268
rect 52828 24216 52880 24268
rect 57888 24216 57940 24268
rect 43996 24080 44048 24132
rect 44548 24080 44600 24132
rect 45376 24191 45428 24200
rect 45376 24157 45385 24191
rect 45385 24157 45419 24191
rect 45419 24157 45428 24191
rect 47860 24191 47912 24200
rect 45376 24148 45428 24157
rect 47860 24157 47869 24191
rect 47869 24157 47903 24191
rect 47903 24157 47912 24191
rect 47860 24148 47912 24157
rect 48044 24191 48096 24200
rect 48044 24157 48053 24191
rect 48053 24157 48087 24191
rect 48087 24157 48096 24191
rect 48044 24148 48096 24157
rect 52276 24148 52328 24200
rect 52736 24148 52788 24200
rect 53656 24148 53708 24200
rect 55312 24191 55364 24200
rect 55312 24157 55321 24191
rect 55321 24157 55355 24191
rect 55355 24157 55364 24191
rect 55312 24148 55364 24157
rect 55404 24191 55456 24200
rect 55404 24157 55413 24191
rect 55413 24157 55447 24191
rect 55447 24157 55456 24191
rect 55588 24191 55640 24200
rect 55404 24148 55456 24157
rect 55588 24157 55597 24191
rect 55597 24157 55631 24191
rect 55631 24157 55640 24191
rect 55588 24148 55640 24157
rect 55680 24191 55732 24200
rect 55680 24157 55689 24191
rect 55689 24157 55723 24191
rect 55723 24157 55732 24191
rect 55680 24148 55732 24157
rect 56692 24123 56744 24132
rect 56692 24089 56701 24123
rect 56701 24089 56735 24123
rect 56735 24089 56744 24123
rect 56692 24080 56744 24089
rect 56784 24080 56836 24132
rect 37372 24012 37424 24064
rect 38384 24012 38436 24064
rect 43536 24012 43588 24064
rect 56324 24012 56376 24064
rect 19574 23910 19626 23962
rect 19638 23910 19690 23962
rect 19702 23910 19754 23962
rect 19766 23910 19818 23962
rect 19830 23910 19882 23962
rect 50294 23910 50346 23962
rect 50358 23910 50410 23962
rect 50422 23910 50474 23962
rect 50486 23910 50538 23962
rect 50550 23910 50602 23962
rect 9404 23851 9456 23860
rect 2596 23740 2648 23792
rect 4068 23740 4120 23792
rect 9404 23817 9413 23851
rect 9413 23817 9447 23851
rect 9447 23817 9456 23851
rect 9404 23808 9456 23817
rect 10324 23851 10376 23860
rect 10324 23817 10333 23851
rect 10333 23817 10367 23851
rect 10367 23817 10376 23851
rect 10324 23808 10376 23817
rect 10784 23851 10836 23860
rect 10784 23817 10793 23851
rect 10793 23817 10827 23851
rect 10827 23817 10836 23851
rect 10784 23808 10836 23817
rect 12808 23808 12860 23860
rect 14556 23808 14608 23860
rect 17224 23851 17276 23860
rect 17224 23817 17233 23851
rect 17233 23817 17267 23851
rect 17267 23817 17276 23851
rect 17224 23808 17276 23817
rect 18144 23808 18196 23860
rect 19248 23808 19300 23860
rect 19340 23808 19392 23860
rect 20168 23808 20220 23860
rect 20352 23808 20404 23860
rect 20536 23808 20588 23860
rect 2504 23715 2556 23724
rect 2504 23681 2513 23715
rect 2513 23681 2547 23715
rect 2547 23681 2556 23715
rect 2504 23672 2556 23681
rect 5448 23715 5500 23724
rect 5448 23681 5457 23715
rect 5457 23681 5491 23715
rect 5491 23681 5500 23715
rect 5448 23672 5500 23681
rect 7656 23740 7708 23792
rect 9956 23783 10008 23792
rect 9956 23749 9965 23783
rect 9965 23749 9999 23783
rect 9999 23749 10008 23783
rect 9956 23740 10008 23749
rect 7748 23715 7800 23724
rect 7748 23681 7757 23715
rect 7757 23681 7791 23715
rect 7791 23681 7800 23715
rect 7748 23672 7800 23681
rect 9312 23672 9364 23724
rect 10140 23672 10192 23724
rect 12440 23715 12492 23724
rect 12440 23681 12449 23715
rect 12449 23681 12483 23715
rect 12483 23681 12492 23715
rect 12440 23672 12492 23681
rect 7012 23604 7064 23656
rect 12532 23604 12584 23656
rect 9220 23579 9272 23588
rect 9220 23545 9229 23579
rect 9229 23545 9263 23579
rect 9263 23545 9272 23579
rect 9220 23536 9272 23545
rect 12992 23579 13044 23588
rect 4804 23511 4856 23520
rect 4804 23477 4813 23511
rect 4813 23477 4847 23511
rect 4847 23477 4856 23511
rect 4804 23468 4856 23477
rect 8024 23468 8076 23520
rect 12992 23545 13001 23579
rect 13001 23545 13035 23579
rect 13035 23545 13044 23579
rect 12992 23536 13044 23545
rect 10600 23468 10652 23520
rect 12532 23468 12584 23520
rect 16764 23740 16816 23792
rect 17868 23740 17920 23792
rect 20720 23808 20772 23860
rect 21180 23808 21232 23860
rect 21364 23808 21416 23860
rect 23020 23851 23072 23860
rect 23020 23817 23029 23851
rect 23029 23817 23063 23851
rect 23063 23817 23072 23851
rect 23020 23808 23072 23817
rect 13636 23715 13688 23724
rect 13636 23681 13645 23715
rect 13645 23681 13679 23715
rect 13679 23681 13688 23715
rect 13636 23672 13688 23681
rect 14556 23672 14608 23724
rect 13544 23604 13596 23656
rect 16580 23672 16632 23724
rect 16948 23715 17000 23724
rect 16948 23681 16957 23715
rect 16957 23681 16991 23715
rect 16991 23681 17000 23715
rect 16948 23672 17000 23681
rect 17040 23715 17092 23724
rect 17040 23681 17049 23715
rect 17049 23681 17083 23715
rect 17083 23681 17092 23715
rect 17040 23672 17092 23681
rect 14096 23468 14148 23520
rect 17776 23604 17828 23656
rect 18420 23672 18472 23724
rect 18972 23672 19024 23724
rect 19432 23672 19484 23724
rect 20168 23672 20220 23724
rect 20904 23740 20956 23792
rect 20996 23672 21048 23724
rect 18328 23604 18380 23656
rect 19984 23604 20036 23656
rect 23572 23740 23624 23792
rect 24952 23783 25004 23792
rect 24952 23749 24961 23783
rect 24961 23749 24995 23783
rect 24995 23749 25004 23783
rect 24952 23740 25004 23749
rect 25964 23783 26016 23792
rect 23756 23672 23808 23724
rect 23940 23715 23992 23724
rect 23940 23681 23949 23715
rect 23949 23681 23983 23715
rect 23983 23681 23992 23715
rect 23940 23672 23992 23681
rect 18052 23536 18104 23588
rect 18420 23536 18472 23588
rect 20536 23536 20588 23588
rect 18972 23468 19024 23520
rect 19340 23468 19392 23520
rect 21640 23536 21692 23588
rect 23664 23604 23716 23656
rect 24308 23536 24360 23588
rect 24768 23604 24820 23656
rect 25044 23715 25096 23724
rect 25044 23681 25058 23715
rect 25058 23681 25092 23715
rect 25092 23681 25096 23715
rect 25044 23672 25096 23681
rect 25964 23749 25973 23783
rect 25973 23749 26007 23783
rect 26007 23749 26016 23783
rect 25964 23740 26016 23749
rect 31300 23808 31352 23860
rect 23572 23468 23624 23520
rect 25412 23468 25464 23520
rect 27712 23468 27764 23520
rect 28816 23468 28868 23520
rect 29644 23511 29696 23520
rect 29644 23477 29653 23511
rect 29653 23477 29687 23511
rect 29687 23477 29696 23511
rect 31116 23604 31168 23656
rect 35440 23740 35492 23792
rect 34704 23672 34756 23724
rect 34888 23715 34940 23724
rect 34888 23681 34897 23715
rect 34897 23681 34931 23715
rect 34931 23681 34940 23715
rect 37280 23715 37332 23724
rect 34888 23672 34940 23681
rect 37280 23681 37289 23715
rect 37289 23681 37323 23715
rect 37323 23681 37332 23715
rect 37280 23672 37332 23681
rect 37464 23715 37516 23724
rect 37464 23681 37473 23715
rect 37473 23681 37507 23715
rect 37507 23681 37516 23715
rect 37464 23672 37516 23681
rect 37740 23715 37792 23724
rect 37740 23681 37749 23715
rect 37749 23681 37783 23715
rect 37783 23681 37792 23715
rect 37740 23672 37792 23681
rect 41052 23740 41104 23792
rect 43536 23740 43588 23792
rect 43996 23740 44048 23792
rect 47308 23808 47360 23860
rect 47860 23808 47912 23860
rect 48044 23851 48096 23860
rect 48044 23817 48053 23851
rect 48053 23817 48087 23851
rect 48087 23817 48096 23851
rect 48044 23808 48096 23817
rect 53196 23851 53248 23860
rect 53196 23817 53205 23851
rect 53205 23817 53239 23851
rect 53239 23817 53248 23851
rect 53196 23808 53248 23817
rect 55772 23808 55824 23860
rect 40132 23715 40184 23724
rect 40132 23681 40141 23715
rect 40141 23681 40175 23715
rect 40175 23681 40184 23715
rect 40132 23672 40184 23681
rect 49516 23740 49568 23792
rect 50252 23672 50304 23724
rect 50620 23672 50672 23724
rect 51080 23672 51132 23724
rect 55312 23740 55364 23792
rect 52276 23672 52328 23724
rect 55680 23672 55732 23724
rect 47584 23647 47636 23656
rect 47584 23613 47593 23647
rect 47593 23613 47627 23647
rect 47627 23613 47636 23647
rect 47584 23604 47636 23613
rect 52736 23647 52788 23656
rect 52736 23613 52745 23647
rect 52745 23613 52779 23647
rect 52779 23613 52788 23647
rect 52736 23604 52788 23613
rect 45376 23536 45428 23588
rect 47400 23536 47452 23588
rect 52276 23536 52328 23588
rect 29644 23468 29696 23477
rect 36544 23468 36596 23520
rect 36728 23511 36780 23520
rect 36728 23477 36737 23511
rect 36737 23477 36771 23511
rect 36771 23477 36780 23511
rect 36728 23468 36780 23477
rect 37464 23468 37516 23520
rect 41604 23468 41656 23520
rect 43904 23511 43956 23520
rect 43904 23477 43913 23511
rect 43913 23477 43947 23511
rect 43947 23477 43956 23511
rect 43904 23468 43956 23477
rect 52092 23468 52144 23520
rect 52828 23511 52880 23520
rect 52828 23477 52837 23511
rect 52837 23477 52871 23511
rect 52871 23477 52880 23511
rect 52828 23468 52880 23477
rect 57888 23468 57940 23520
rect 4214 23366 4266 23418
rect 4278 23366 4330 23418
rect 4342 23366 4394 23418
rect 4406 23366 4458 23418
rect 4470 23366 4522 23418
rect 34934 23366 34986 23418
rect 34998 23366 35050 23418
rect 35062 23366 35114 23418
rect 35126 23366 35178 23418
rect 35190 23366 35242 23418
rect 6828 23264 6880 23316
rect 7288 23264 7340 23316
rect 7748 23196 7800 23248
rect 9312 23264 9364 23316
rect 9496 23264 9548 23316
rect 15476 23264 15528 23316
rect 20812 23264 20864 23316
rect 23756 23264 23808 23316
rect 24492 23264 24544 23316
rect 31116 23264 31168 23316
rect 35440 23264 35492 23316
rect 55312 23264 55364 23316
rect 55496 23307 55548 23316
rect 55496 23273 55505 23307
rect 55505 23273 55539 23307
rect 55539 23273 55548 23307
rect 55496 23264 55548 23273
rect 12808 23196 12860 23248
rect 13820 23196 13872 23248
rect 6184 23171 6236 23180
rect 6184 23137 6193 23171
rect 6193 23137 6227 23171
rect 6227 23137 6236 23171
rect 6184 23128 6236 23137
rect 7012 23171 7064 23180
rect 7012 23137 7021 23171
rect 7021 23137 7055 23171
rect 7055 23137 7064 23171
rect 7012 23128 7064 23137
rect 1860 23103 1912 23112
rect 1860 23069 1869 23103
rect 1869 23069 1903 23103
rect 1903 23069 1912 23103
rect 1860 23060 1912 23069
rect 4620 23060 4672 23112
rect 8024 23103 8076 23112
rect 2044 23035 2096 23044
rect 2044 23001 2053 23035
rect 2053 23001 2087 23035
rect 2087 23001 2096 23035
rect 2044 22992 2096 23001
rect 4804 22992 4856 23044
rect 8024 23069 8033 23103
rect 8033 23069 8067 23103
rect 8067 23069 8076 23103
rect 8024 23060 8076 23069
rect 9864 23103 9916 23112
rect 9864 23069 9873 23103
rect 9873 23069 9907 23103
rect 9907 23069 9916 23103
rect 9864 23060 9916 23069
rect 10140 23103 10192 23112
rect 10140 23069 10149 23103
rect 10149 23069 10183 23103
rect 10183 23069 10192 23103
rect 10140 23060 10192 23069
rect 12624 23060 12676 23112
rect 13636 23060 13688 23112
rect 15016 23128 15068 23180
rect 20260 23196 20312 23248
rect 21640 23196 21692 23248
rect 23020 23196 23072 23248
rect 24768 23196 24820 23248
rect 37740 23196 37792 23248
rect 52736 23196 52788 23248
rect 16488 23128 16540 23180
rect 15384 23060 15436 23112
rect 16396 23060 16448 23112
rect 18328 23128 18380 23180
rect 19984 23128 20036 23180
rect 17684 23103 17736 23112
rect 17684 23069 17693 23103
rect 17693 23069 17727 23103
rect 17727 23069 17736 23103
rect 17684 23060 17736 23069
rect 11520 22924 11572 22976
rect 13728 22924 13780 22976
rect 16120 22992 16172 23044
rect 16764 23035 16816 23044
rect 16764 23001 16773 23035
rect 16773 23001 16807 23035
rect 16807 23001 16816 23035
rect 16764 22992 16816 23001
rect 17592 23035 17644 23044
rect 17592 23001 17601 23035
rect 17601 23001 17635 23035
rect 17635 23001 17644 23035
rect 17592 22992 17644 23001
rect 20076 23060 20128 23112
rect 20996 23060 21048 23112
rect 23480 23060 23532 23112
rect 23756 23060 23808 23112
rect 24860 23103 24912 23112
rect 24860 23069 24869 23103
rect 24869 23069 24903 23103
rect 24903 23069 24912 23103
rect 24860 23060 24912 23069
rect 26424 23060 26476 23112
rect 26792 23103 26844 23112
rect 26792 23069 26801 23103
rect 26801 23069 26835 23103
rect 26835 23069 26844 23103
rect 26792 23060 26844 23069
rect 27804 23060 27856 23112
rect 28816 23103 28868 23112
rect 28816 23069 28825 23103
rect 28825 23069 28859 23103
rect 28859 23069 28868 23103
rect 28816 23060 28868 23069
rect 20168 22992 20220 23044
rect 21456 22992 21508 23044
rect 30380 23060 30432 23112
rect 43996 23171 44048 23180
rect 43996 23137 44005 23171
rect 44005 23137 44039 23171
rect 44039 23137 44048 23171
rect 43996 23128 44048 23137
rect 51080 23128 51132 23180
rect 52092 23171 52144 23180
rect 52092 23137 52101 23171
rect 52101 23137 52135 23171
rect 52135 23137 52144 23171
rect 52092 23128 52144 23137
rect 53288 23128 53340 23180
rect 14464 22967 14516 22976
rect 14464 22933 14473 22967
rect 14473 22933 14507 22967
rect 14507 22933 14516 22967
rect 14464 22924 14516 22933
rect 19156 22924 19208 22976
rect 20076 22924 20128 22976
rect 20904 22924 20956 22976
rect 24952 22967 25004 22976
rect 24952 22933 24961 22967
rect 24961 22933 24995 22967
rect 24995 22933 25004 22967
rect 24952 22924 25004 22933
rect 30288 22992 30340 23044
rect 31576 23060 31628 23112
rect 42800 23060 42852 23112
rect 43904 23103 43956 23112
rect 43904 23069 43913 23103
rect 43913 23069 43947 23103
rect 43947 23069 43956 23103
rect 43904 23060 43956 23069
rect 46020 23103 46072 23112
rect 46020 23069 46029 23103
rect 46029 23069 46063 23103
rect 46063 23069 46072 23103
rect 46020 23060 46072 23069
rect 46296 23103 46348 23112
rect 46296 23069 46305 23103
rect 46305 23069 46339 23103
rect 46339 23069 46348 23103
rect 46296 23060 46348 23069
rect 47308 23103 47360 23112
rect 47308 23069 47317 23103
rect 47317 23069 47351 23103
rect 47351 23069 47360 23103
rect 47308 23060 47360 23069
rect 47400 23103 47452 23112
rect 47400 23069 47409 23103
rect 47409 23069 47443 23103
rect 47443 23069 47452 23103
rect 47584 23103 47636 23112
rect 47400 23060 47452 23069
rect 47584 23069 47593 23103
rect 47593 23069 47627 23103
rect 47627 23069 47636 23103
rect 47584 23060 47636 23069
rect 50252 23103 50304 23112
rect 50252 23069 50261 23103
rect 50261 23069 50295 23103
rect 50295 23069 50304 23103
rect 50252 23060 50304 23069
rect 50620 23060 50672 23112
rect 52276 23060 52328 23112
rect 53012 23060 53064 23112
rect 34704 22992 34756 23044
rect 34888 22992 34940 23044
rect 54484 23103 54536 23112
rect 54484 23069 54493 23103
rect 54493 23069 54527 23103
rect 54527 23069 54536 23103
rect 54484 23060 54536 23069
rect 55496 23060 55548 23112
rect 56508 23103 56560 23112
rect 56508 23069 56517 23103
rect 56517 23069 56551 23103
rect 56551 23069 56560 23103
rect 56508 23060 56560 23069
rect 57060 23103 57112 23112
rect 57060 23069 57069 23103
rect 57069 23069 57103 23103
rect 57103 23069 57112 23103
rect 57060 23060 57112 23069
rect 53748 22992 53800 23044
rect 57704 22992 57756 23044
rect 27712 22924 27764 22976
rect 29828 22924 29880 22976
rect 33508 22967 33560 22976
rect 33508 22933 33517 22967
rect 33517 22933 33551 22967
rect 33551 22933 33560 22967
rect 33508 22924 33560 22933
rect 34612 22924 34664 22976
rect 35624 22967 35676 22976
rect 35624 22933 35633 22967
rect 35633 22933 35667 22967
rect 35667 22933 35676 22967
rect 35624 22924 35676 22933
rect 43536 22967 43588 22976
rect 43536 22933 43545 22967
rect 43545 22933 43579 22967
rect 43579 22933 43588 22967
rect 43536 22924 43588 22933
rect 46112 22967 46164 22976
rect 46112 22933 46121 22967
rect 46121 22933 46155 22967
rect 46155 22933 46164 22967
rect 46112 22924 46164 22933
rect 54484 22924 54536 22976
rect 55680 22967 55732 22976
rect 55680 22933 55689 22967
rect 55689 22933 55723 22967
rect 55723 22933 55732 22967
rect 55680 22924 55732 22933
rect 19574 22822 19626 22874
rect 19638 22822 19690 22874
rect 19702 22822 19754 22874
rect 19766 22822 19818 22874
rect 19830 22822 19882 22874
rect 50294 22822 50346 22874
rect 50358 22822 50410 22874
rect 50422 22822 50474 22874
rect 50486 22822 50538 22874
rect 50550 22822 50602 22874
rect 1860 22720 1912 22772
rect 4620 22720 4672 22772
rect 5264 22720 5316 22772
rect 6184 22720 6236 22772
rect 8484 22720 8536 22772
rect 4068 22652 4120 22704
rect 8760 22695 8812 22704
rect 8760 22661 8769 22695
rect 8769 22661 8803 22695
rect 8803 22661 8812 22695
rect 8760 22652 8812 22661
rect 9864 22652 9916 22704
rect 3608 22584 3660 22636
rect 6828 22584 6880 22636
rect 7656 22627 7708 22636
rect 7656 22593 7665 22627
rect 7665 22593 7699 22627
rect 7699 22593 7708 22627
rect 7656 22584 7708 22593
rect 8300 22584 8352 22636
rect 12900 22652 12952 22704
rect 10600 22584 10652 22636
rect 12808 22627 12860 22636
rect 12808 22593 12817 22627
rect 12817 22593 12851 22627
rect 12851 22593 12860 22627
rect 12808 22584 12860 22593
rect 12992 22627 13044 22636
rect 12992 22593 13001 22627
rect 13001 22593 13035 22627
rect 13035 22593 13044 22627
rect 12992 22584 13044 22593
rect 13084 22516 13136 22568
rect 4620 22423 4672 22432
rect 4620 22389 4629 22423
rect 4629 22389 4663 22423
rect 4663 22389 4672 22423
rect 4620 22380 4672 22389
rect 9772 22380 9824 22432
rect 15384 22720 15436 22772
rect 17500 22720 17552 22772
rect 19248 22720 19300 22772
rect 14464 22652 14516 22704
rect 14004 22627 14056 22636
rect 14004 22593 14011 22627
rect 14011 22593 14056 22627
rect 14004 22584 14056 22593
rect 14188 22627 14240 22636
rect 14188 22593 14197 22627
rect 14197 22593 14231 22627
rect 14231 22593 14240 22627
rect 14188 22584 14240 22593
rect 14924 22584 14976 22636
rect 15016 22584 15068 22636
rect 16488 22584 16540 22636
rect 14280 22448 14332 22500
rect 14464 22491 14516 22500
rect 14464 22457 14473 22491
rect 14473 22457 14507 22491
rect 14507 22457 14516 22491
rect 14464 22448 14516 22457
rect 15108 22448 15160 22500
rect 17040 22627 17092 22636
rect 17040 22593 17049 22627
rect 17049 22593 17083 22627
rect 17083 22593 17092 22627
rect 19156 22627 19208 22636
rect 17040 22584 17092 22593
rect 19156 22593 19165 22627
rect 19165 22593 19199 22627
rect 19199 22593 19208 22627
rect 19156 22584 19208 22593
rect 19340 22627 19392 22636
rect 19340 22593 19347 22627
rect 19347 22593 19392 22627
rect 19340 22584 19392 22593
rect 19984 22720 20036 22772
rect 20720 22720 20772 22772
rect 20812 22652 20864 22704
rect 20996 22584 21048 22636
rect 21824 22627 21876 22636
rect 21824 22593 21833 22627
rect 21833 22593 21867 22627
rect 21867 22593 21876 22627
rect 21824 22584 21876 22593
rect 23480 22720 23532 22772
rect 28816 22720 28868 22772
rect 30288 22763 30340 22772
rect 30288 22729 30297 22763
rect 30297 22729 30331 22763
rect 30331 22729 30340 22763
rect 30288 22720 30340 22729
rect 34704 22720 34756 22772
rect 34796 22720 34848 22772
rect 35440 22763 35492 22772
rect 35440 22729 35449 22763
rect 35449 22729 35483 22763
rect 35483 22729 35492 22763
rect 35440 22720 35492 22729
rect 38108 22720 38160 22772
rect 43536 22720 43588 22772
rect 46020 22720 46072 22772
rect 47584 22720 47636 22772
rect 52828 22720 52880 22772
rect 57060 22763 57112 22772
rect 57060 22729 57069 22763
rect 57069 22729 57103 22763
rect 57103 22729 57112 22763
rect 57060 22720 57112 22729
rect 33508 22652 33560 22704
rect 20352 22516 20404 22568
rect 20628 22516 20680 22568
rect 22192 22627 22244 22636
rect 22192 22593 22201 22627
rect 22201 22593 22235 22627
rect 22235 22593 22244 22627
rect 22192 22584 22244 22593
rect 23572 22584 23624 22636
rect 24032 22584 24084 22636
rect 24216 22584 24268 22636
rect 24492 22584 24544 22636
rect 23664 22448 23716 22500
rect 29828 22584 29880 22636
rect 30380 22627 30432 22636
rect 30380 22593 30389 22627
rect 30389 22593 30423 22627
rect 30423 22593 30432 22627
rect 30380 22584 30432 22593
rect 32956 22584 33008 22636
rect 35624 22652 35676 22704
rect 46296 22695 46348 22704
rect 46296 22661 46305 22695
rect 46305 22661 46339 22695
rect 46339 22661 46348 22695
rect 46296 22652 46348 22661
rect 50620 22652 50672 22704
rect 52276 22652 52328 22704
rect 34612 22627 34664 22636
rect 34612 22593 34621 22627
rect 34621 22593 34655 22627
rect 34655 22593 34664 22627
rect 34612 22584 34664 22593
rect 35440 22627 35492 22636
rect 33324 22516 33376 22568
rect 35440 22593 35449 22627
rect 35449 22593 35483 22627
rect 35483 22593 35492 22627
rect 35440 22584 35492 22593
rect 33508 22448 33560 22500
rect 15936 22380 15988 22432
rect 22008 22380 22060 22432
rect 24400 22380 24452 22432
rect 34520 22448 34572 22500
rect 34612 22448 34664 22500
rect 35808 22584 35860 22636
rect 38936 22584 38988 22636
rect 40224 22627 40276 22636
rect 40224 22593 40233 22627
rect 40233 22593 40267 22627
rect 40267 22593 40276 22627
rect 40224 22584 40276 22593
rect 42524 22627 42576 22636
rect 42524 22593 42533 22627
rect 42533 22593 42567 22627
rect 42567 22593 42576 22627
rect 42524 22584 42576 22593
rect 42984 22584 43036 22636
rect 49332 22627 49384 22636
rect 49332 22593 49341 22627
rect 49341 22593 49375 22627
rect 49375 22593 49384 22627
rect 49332 22584 49384 22593
rect 49700 22584 49752 22636
rect 52092 22584 52144 22636
rect 53748 22652 53800 22704
rect 56508 22695 56560 22704
rect 56508 22661 56517 22695
rect 56517 22661 56551 22695
rect 56551 22661 56560 22695
rect 56508 22652 56560 22661
rect 53012 22627 53064 22636
rect 53012 22593 53021 22627
rect 53021 22593 53055 22627
rect 53055 22593 53064 22627
rect 53012 22584 53064 22593
rect 53288 22584 53340 22636
rect 53656 22584 53708 22636
rect 56232 22627 56284 22636
rect 40132 22559 40184 22568
rect 36636 22491 36688 22500
rect 36636 22457 36645 22491
rect 36645 22457 36679 22491
rect 36679 22457 36688 22491
rect 40132 22525 40141 22559
rect 40141 22525 40175 22559
rect 40175 22525 40184 22559
rect 40132 22516 40184 22525
rect 40592 22559 40644 22568
rect 40592 22525 40601 22559
rect 40601 22525 40635 22559
rect 40635 22525 40644 22559
rect 40592 22516 40644 22525
rect 56232 22593 56241 22627
rect 56241 22593 56275 22627
rect 56275 22593 56284 22627
rect 56232 22584 56284 22593
rect 56324 22627 56376 22636
rect 56324 22593 56333 22627
rect 56333 22593 56367 22627
rect 56367 22593 56376 22627
rect 56324 22584 56376 22593
rect 56692 22584 56744 22636
rect 57152 22627 57204 22636
rect 57152 22593 57161 22627
rect 57161 22593 57195 22627
rect 57195 22593 57204 22627
rect 57152 22584 57204 22593
rect 55496 22516 55548 22568
rect 36636 22448 36688 22457
rect 54484 22448 54536 22500
rect 36728 22380 36780 22432
rect 42892 22423 42944 22432
rect 42892 22389 42901 22423
rect 42901 22389 42935 22423
rect 42935 22389 42944 22423
rect 42892 22380 42944 22389
rect 46112 22380 46164 22432
rect 46572 22380 46624 22432
rect 4214 22278 4266 22330
rect 4278 22278 4330 22330
rect 4342 22278 4394 22330
rect 4406 22278 4458 22330
rect 4470 22278 4522 22330
rect 34934 22278 34986 22330
rect 34998 22278 35050 22330
rect 35062 22278 35114 22330
rect 35126 22278 35178 22330
rect 35190 22278 35242 22330
rect 10600 22176 10652 22228
rect 13084 22176 13136 22228
rect 13360 22176 13412 22228
rect 13728 22176 13780 22228
rect 15752 22219 15804 22228
rect 15752 22185 15761 22219
rect 15761 22185 15795 22219
rect 15795 22185 15804 22219
rect 15752 22176 15804 22185
rect 16488 22176 16540 22228
rect 20628 22176 20680 22228
rect 21824 22176 21876 22228
rect 23112 22176 23164 22228
rect 7472 22151 7524 22160
rect 7472 22117 7481 22151
rect 7481 22117 7515 22151
rect 7515 22117 7524 22151
rect 7472 22108 7524 22117
rect 2136 21972 2188 22024
rect 2780 21972 2832 22024
rect 9864 22040 9916 22092
rect 12900 22108 12952 22160
rect 17592 22108 17644 22160
rect 19432 22108 19484 22160
rect 33600 22176 33652 22228
rect 35440 22176 35492 22228
rect 35808 22176 35860 22228
rect 37188 22219 37240 22228
rect 37188 22185 37197 22219
rect 37197 22185 37231 22219
rect 37231 22185 37240 22219
rect 37188 22176 37240 22185
rect 40132 22176 40184 22228
rect 42524 22219 42576 22228
rect 42524 22185 42533 22219
rect 42533 22185 42567 22219
rect 42567 22185 42576 22219
rect 42524 22176 42576 22185
rect 42800 22219 42852 22228
rect 42800 22185 42809 22219
rect 42809 22185 42843 22219
rect 42843 22185 42852 22219
rect 42800 22176 42852 22185
rect 46020 22176 46072 22228
rect 46572 22219 46624 22228
rect 46572 22185 46581 22219
rect 46581 22185 46615 22219
rect 46615 22185 46624 22219
rect 46572 22176 46624 22185
rect 2872 21904 2924 21956
rect 4896 21972 4948 22024
rect 5080 22015 5132 22024
rect 5080 21981 5089 22015
rect 5089 21981 5123 22015
rect 5123 21981 5132 22015
rect 5080 21972 5132 21981
rect 7104 21972 7156 22024
rect 7656 21972 7708 22024
rect 8024 21972 8076 22024
rect 9404 21972 9456 22024
rect 9956 22015 10008 22024
rect 9956 21981 9965 22015
rect 9965 21981 9999 22015
rect 9999 21981 10008 22015
rect 9956 21972 10008 21981
rect 10048 22015 10100 22024
rect 10048 21981 10057 22015
rect 10057 21981 10091 22015
rect 10091 21981 10100 22015
rect 10876 22040 10928 22092
rect 14280 22040 14332 22092
rect 14924 22040 14976 22092
rect 15016 22040 15068 22092
rect 21824 22040 21876 22092
rect 27804 22108 27856 22160
rect 33508 22108 33560 22160
rect 34796 22108 34848 22160
rect 35348 22108 35400 22160
rect 30564 22083 30616 22092
rect 10048 21972 10100 21981
rect 10784 21972 10836 22024
rect 11060 22015 11112 22024
rect 11060 21981 11069 22015
rect 11069 21981 11103 22015
rect 11103 21981 11112 22015
rect 11060 21972 11112 21981
rect 13176 21972 13228 22024
rect 13544 21972 13596 22024
rect 16304 22015 16356 22024
rect 16304 21981 16313 22015
rect 16313 21981 16347 22015
rect 16347 21981 16356 22015
rect 16304 21972 16356 21981
rect 2688 21836 2740 21888
rect 3148 21879 3200 21888
rect 3148 21845 3157 21879
rect 3157 21845 3191 21879
rect 3191 21845 3200 21879
rect 15752 21904 15804 21956
rect 19892 21972 19944 22024
rect 20628 21972 20680 22024
rect 20720 22015 20772 22024
rect 20720 21981 20729 22015
rect 20729 21981 20763 22015
rect 20763 21981 20772 22015
rect 20720 21972 20772 21981
rect 21456 22015 21508 22024
rect 16488 21904 16540 21956
rect 4160 21879 4212 21888
rect 3148 21836 3200 21845
rect 4160 21845 4169 21879
rect 4169 21845 4203 21879
rect 4203 21845 4212 21879
rect 4160 21836 4212 21845
rect 6736 21836 6788 21888
rect 9312 21879 9364 21888
rect 9312 21845 9337 21879
rect 9337 21845 9364 21879
rect 9312 21836 9364 21845
rect 10048 21836 10100 21888
rect 10508 21879 10560 21888
rect 10508 21845 10517 21879
rect 10517 21845 10551 21879
rect 10551 21845 10560 21879
rect 10508 21836 10560 21845
rect 11244 21879 11296 21888
rect 11244 21845 11253 21879
rect 11253 21845 11287 21879
rect 11287 21845 11296 21879
rect 11244 21836 11296 21845
rect 13176 21836 13228 21888
rect 15200 21836 15252 21888
rect 19340 21879 19392 21888
rect 19340 21845 19349 21879
rect 19349 21845 19383 21879
rect 19383 21845 19392 21879
rect 19340 21836 19392 21845
rect 20168 21836 20220 21888
rect 21088 21836 21140 21888
rect 21456 21981 21465 22015
rect 21465 21981 21499 22015
rect 21499 21981 21508 22015
rect 21456 21972 21508 21981
rect 21548 22015 21600 22024
rect 21548 21981 21557 22015
rect 21557 21981 21591 22015
rect 21591 21981 21600 22015
rect 21548 21972 21600 21981
rect 23664 21972 23716 22024
rect 24400 22015 24452 22024
rect 21364 21947 21416 21956
rect 21364 21913 21373 21947
rect 21373 21913 21407 21947
rect 21407 21913 21416 21947
rect 21364 21904 21416 21913
rect 21732 21904 21784 21956
rect 21640 21836 21692 21888
rect 22100 21836 22152 21888
rect 24124 21904 24176 21956
rect 24400 21981 24409 22015
rect 24409 21981 24443 22015
rect 24443 21981 24452 22015
rect 24400 21972 24452 21981
rect 30564 22049 30573 22083
rect 30573 22049 30607 22083
rect 30607 22049 30616 22083
rect 30564 22040 30616 22049
rect 30840 22040 30892 22092
rect 36820 22083 36872 22092
rect 36820 22049 36829 22083
rect 36829 22049 36863 22083
rect 36863 22049 36872 22083
rect 36820 22040 36872 22049
rect 38200 22040 38252 22092
rect 24768 22015 24820 22024
rect 24768 21981 24777 22015
rect 24777 21981 24811 22015
rect 24811 21981 24820 22015
rect 24768 21972 24820 21981
rect 34520 21972 34572 22024
rect 37280 21972 37332 22024
rect 38936 22015 38988 22024
rect 38936 21981 38945 22015
rect 38945 21981 38979 22015
rect 38979 21981 38988 22015
rect 38936 21972 38988 21981
rect 39028 21972 39080 22024
rect 42892 21972 42944 22024
rect 42984 22015 43036 22024
rect 42984 21981 42993 22015
rect 42993 21981 43027 22015
rect 43027 21981 43036 22015
rect 45652 22015 45704 22024
rect 42984 21972 43036 21981
rect 45652 21981 45661 22015
rect 45661 21981 45695 22015
rect 45695 21981 45704 22015
rect 45652 21972 45704 21981
rect 46480 21972 46532 22024
rect 57060 22040 57112 22092
rect 23572 21836 23624 21888
rect 25320 21836 25372 21888
rect 32680 21904 32732 21956
rect 40316 21947 40368 21956
rect 40316 21913 40325 21947
rect 40325 21913 40359 21947
rect 40359 21913 40368 21947
rect 40316 21904 40368 21913
rect 26792 21879 26844 21888
rect 26792 21845 26801 21879
rect 26801 21845 26835 21879
rect 26835 21845 26844 21879
rect 26792 21836 26844 21845
rect 29828 21836 29880 21888
rect 33048 21836 33100 21888
rect 33324 21879 33376 21888
rect 33324 21845 33333 21879
rect 33333 21845 33367 21879
rect 33367 21845 33376 21879
rect 33324 21836 33376 21845
rect 34704 21836 34756 21888
rect 38200 21879 38252 21888
rect 38200 21845 38209 21879
rect 38209 21845 38243 21879
rect 38243 21845 38252 21879
rect 38200 21836 38252 21845
rect 45836 21836 45888 21888
rect 57152 21972 57204 22024
rect 57980 21904 58032 21956
rect 55680 21836 55732 21888
rect 19574 21734 19626 21786
rect 19638 21734 19690 21786
rect 19702 21734 19754 21786
rect 19766 21734 19818 21786
rect 19830 21734 19882 21786
rect 50294 21734 50346 21786
rect 50358 21734 50410 21786
rect 50422 21734 50474 21786
rect 50486 21734 50538 21786
rect 50550 21734 50602 21786
rect 2872 21632 2924 21684
rect 1400 21539 1452 21548
rect 1400 21505 1409 21539
rect 1409 21505 1443 21539
rect 1443 21505 1452 21539
rect 1400 21496 1452 21505
rect 2228 21496 2280 21548
rect 2780 21471 2832 21480
rect 2780 21437 2789 21471
rect 2789 21437 2823 21471
rect 2823 21437 2832 21471
rect 2780 21428 2832 21437
rect 4620 21632 4672 21684
rect 5172 21632 5224 21684
rect 9956 21632 10008 21684
rect 11520 21675 11572 21684
rect 5080 21564 5132 21616
rect 9496 21607 9548 21616
rect 4160 21539 4212 21548
rect 4160 21505 4169 21539
rect 4169 21505 4203 21539
rect 4203 21505 4212 21539
rect 4160 21496 4212 21505
rect 4620 21539 4672 21548
rect 4620 21505 4629 21539
rect 4629 21505 4663 21539
rect 4663 21505 4672 21539
rect 4620 21496 4672 21505
rect 6736 21496 6788 21548
rect 7564 21496 7616 21548
rect 9496 21573 9505 21607
rect 9505 21573 9539 21607
rect 9539 21573 9548 21607
rect 9496 21564 9548 21573
rect 9680 21607 9732 21616
rect 9680 21573 9689 21607
rect 9689 21573 9723 21607
rect 9723 21573 9732 21607
rect 11520 21641 11529 21675
rect 11529 21641 11563 21675
rect 11563 21641 11572 21675
rect 11520 21632 11572 21641
rect 13544 21675 13596 21684
rect 13544 21641 13553 21675
rect 13553 21641 13587 21675
rect 13587 21641 13596 21675
rect 13544 21632 13596 21641
rect 15936 21632 15988 21684
rect 16488 21632 16540 21684
rect 20076 21632 20128 21684
rect 9680 21564 9732 21573
rect 9772 21539 9824 21548
rect 9772 21505 9781 21539
rect 9781 21505 9815 21539
rect 9815 21505 9824 21539
rect 9772 21496 9824 21505
rect 9864 21496 9916 21548
rect 14188 21564 14240 21616
rect 17592 21564 17644 21616
rect 18696 21564 18748 21616
rect 12900 21496 12952 21548
rect 13176 21539 13228 21548
rect 13176 21505 13185 21539
rect 13185 21505 13219 21539
rect 13219 21505 13228 21539
rect 13176 21496 13228 21505
rect 11060 21428 11112 21480
rect 11244 21428 11296 21480
rect 13360 21539 13412 21548
rect 13360 21505 13369 21539
rect 13369 21505 13403 21539
rect 13403 21505 13412 21539
rect 13360 21496 13412 21505
rect 14924 21496 14976 21548
rect 19064 21539 19116 21548
rect 19064 21505 19073 21539
rect 19073 21505 19107 21539
rect 19107 21505 19116 21539
rect 19064 21496 19116 21505
rect 19984 21564 20036 21616
rect 20536 21632 20588 21684
rect 20904 21632 20956 21684
rect 21548 21632 21600 21684
rect 23112 21675 23164 21684
rect 23112 21641 23121 21675
rect 23121 21641 23155 21675
rect 23155 21641 23164 21675
rect 23112 21632 23164 21641
rect 23664 21675 23716 21684
rect 23664 21641 23673 21675
rect 23673 21641 23707 21675
rect 23707 21641 23716 21675
rect 23664 21632 23716 21641
rect 25596 21675 25648 21684
rect 20352 21607 20404 21616
rect 20352 21573 20361 21607
rect 20361 21573 20395 21607
rect 20395 21573 20404 21607
rect 20352 21564 20404 21573
rect 21088 21564 21140 21616
rect 8024 21360 8076 21412
rect 1584 21335 1636 21344
rect 1584 21301 1593 21335
rect 1593 21301 1627 21335
rect 1627 21301 1636 21335
rect 1584 21292 1636 21301
rect 5816 21335 5868 21344
rect 5816 21301 5825 21335
rect 5825 21301 5859 21335
rect 5859 21301 5868 21335
rect 5816 21292 5868 21301
rect 18052 21428 18104 21480
rect 19616 21496 19668 21548
rect 12992 21360 13044 21412
rect 22836 21496 22888 21548
rect 24216 21607 24268 21616
rect 24216 21573 24225 21607
rect 24225 21573 24259 21607
rect 24259 21573 24268 21607
rect 24216 21564 24268 21573
rect 25596 21641 25605 21675
rect 25605 21641 25639 21675
rect 25639 21641 25648 21675
rect 25596 21632 25648 21641
rect 31576 21675 31628 21684
rect 31576 21641 31585 21675
rect 31585 21641 31619 21675
rect 31619 21641 31628 21675
rect 31576 21632 31628 21641
rect 31668 21632 31720 21684
rect 32680 21632 32732 21684
rect 32956 21632 33008 21684
rect 34520 21632 34572 21684
rect 34612 21632 34664 21684
rect 39028 21632 39080 21684
rect 24308 21496 24360 21548
rect 26792 21564 26844 21616
rect 27988 21564 28040 21616
rect 25044 21539 25096 21548
rect 25044 21505 25053 21539
rect 25053 21505 25087 21539
rect 25087 21505 25096 21539
rect 25044 21496 25096 21505
rect 25136 21539 25188 21548
rect 25136 21505 25145 21539
rect 25145 21505 25179 21539
rect 25179 21505 25188 21539
rect 25320 21539 25372 21548
rect 25136 21496 25188 21505
rect 25320 21505 25329 21539
rect 25329 21505 25363 21539
rect 25363 21505 25372 21539
rect 25320 21496 25372 21505
rect 25412 21539 25464 21548
rect 25412 21505 25421 21539
rect 25421 21505 25455 21539
rect 25455 21505 25464 21539
rect 25412 21496 25464 21505
rect 26332 21496 26384 21548
rect 27804 21496 27856 21548
rect 30564 21539 30616 21548
rect 30564 21505 30573 21539
rect 30573 21505 30607 21539
rect 30607 21505 30616 21539
rect 30564 21496 30616 21505
rect 35348 21564 35400 21616
rect 45008 21564 45060 21616
rect 49332 21632 49384 21684
rect 53012 21632 53064 21684
rect 53288 21675 53340 21684
rect 53288 21641 53297 21675
rect 53297 21641 53331 21675
rect 53331 21641 53340 21675
rect 53288 21632 53340 21641
rect 54484 21632 54536 21684
rect 56692 21632 56744 21684
rect 57152 21632 57204 21684
rect 57980 21675 58032 21684
rect 57980 21641 57989 21675
rect 57989 21641 58023 21675
rect 58023 21641 58032 21675
rect 57980 21632 58032 21641
rect 16304 21292 16356 21344
rect 17224 21335 17276 21344
rect 17224 21301 17233 21335
rect 17233 21301 17267 21335
rect 17267 21301 17276 21335
rect 17224 21292 17276 21301
rect 18420 21292 18472 21344
rect 18604 21292 18656 21344
rect 25688 21428 25740 21480
rect 34796 21496 34848 21548
rect 45652 21496 45704 21548
rect 48412 21539 48464 21548
rect 48412 21505 48421 21539
rect 48421 21505 48455 21539
rect 48455 21505 48464 21539
rect 48412 21496 48464 21505
rect 49700 21539 49752 21548
rect 49700 21505 49709 21539
rect 49709 21505 49743 21539
rect 49743 21505 49752 21539
rect 49700 21496 49752 21505
rect 53748 21564 53800 21616
rect 37280 21428 37332 21480
rect 45836 21471 45888 21480
rect 45836 21437 45845 21471
rect 45845 21437 45879 21471
rect 45879 21437 45888 21471
rect 45836 21428 45888 21437
rect 46480 21471 46532 21480
rect 46480 21437 46489 21471
rect 46489 21437 46523 21471
rect 46523 21437 46532 21471
rect 46480 21428 46532 21437
rect 48320 21471 48372 21480
rect 48320 21437 48329 21471
rect 48329 21437 48363 21471
rect 48363 21437 48372 21471
rect 48320 21428 48372 21437
rect 51724 21471 51776 21480
rect 51724 21437 51733 21471
rect 51733 21437 51767 21471
rect 51767 21437 51776 21471
rect 51724 21428 51776 21437
rect 20352 21360 20404 21412
rect 21456 21360 21508 21412
rect 21824 21360 21876 21412
rect 26516 21360 26568 21412
rect 36820 21360 36872 21412
rect 49240 21360 49292 21412
rect 54116 21539 54168 21548
rect 54116 21505 54125 21539
rect 54125 21505 54159 21539
rect 54159 21505 54168 21539
rect 54116 21496 54168 21505
rect 54208 21539 54260 21548
rect 54208 21505 54217 21539
rect 54217 21505 54251 21539
rect 54251 21505 54260 21539
rect 54208 21496 54260 21505
rect 56968 21539 57020 21548
rect 56968 21505 56977 21539
rect 56977 21505 57011 21539
rect 57011 21505 57020 21539
rect 56968 21496 57020 21505
rect 57336 21496 57388 21548
rect 20628 21292 20680 21344
rect 20720 21292 20772 21344
rect 22744 21292 22796 21344
rect 23756 21292 23808 21344
rect 24308 21292 24360 21344
rect 25136 21292 25188 21344
rect 25964 21292 26016 21344
rect 29092 21292 29144 21344
rect 30380 21292 30432 21344
rect 37004 21292 37056 21344
rect 43352 21335 43404 21344
rect 43352 21301 43361 21335
rect 43361 21301 43395 21335
rect 43395 21301 43404 21335
rect 43352 21292 43404 21301
rect 51080 21292 51132 21344
rect 51816 21335 51868 21344
rect 51816 21301 51825 21335
rect 51825 21301 51859 21335
rect 51859 21301 51868 21335
rect 55680 21428 55732 21480
rect 51816 21292 51868 21301
rect 4214 21190 4266 21242
rect 4278 21190 4330 21242
rect 4342 21190 4394 21242
rect 4406 21190 4458 21242
rect 4470 21190 4522 21242
rect 34934 21190 34986 21242
rect 34998 21190 35050 21242
rect 35062 21190 35114 21242
rect 35126 21190 35178 21242
rect 35190 21190 35242 21242
rect 1400 21131 1452 21140
rect 1400 21097 1409 21131
rect 1409 21097 1443 21131
rect 1443 21097 1452 21131
rect 1400 21088 1452 21097
rect 3148 21088 3200 21140
rect 9496 21131 9548 21140
rect 9496 21097 9505 21131
rect 9505 21097 9539 21131
rect 9539 21097 9548 21131
rect 9496 21088 9548 21097
rect 9772 21088 9824 21140
rect 13360 21088 13412 21140
rect 14648 21088 14700 21140
rect 14832 21088 14884 21140
rect 5816 21020 5868 21072
rect 14556 21020 14608 21072
rect 2504 20927 2556 20936
rect 2504 20893 2513 20927
rect 2513 20893 2547 20927
rect 2547 20893 2556 20927
rect 2504 20884 2556 20893
rect 2688 20927 2740 20936
rect 2688 20893 2697 20927
rect 2697 20893 2731 20927
rect 2731 20893 2740 20927
rect 2688 20884 2740 20893
rect 4620 20952 4672 21004
rect 5080 20952 5132 21004
rect 6736 20995 6788 21004
rect 6736 20961 6745 20995
rect 6745 20961 6779 20995
rect 6779 20961 6788 20995
rect 6736 20952 6788 20961
rect 7472 20952 7524 21004
rect 13820 20952 13872 21004
rect 4896 20884 4948 20936
rect 7564 20884 7616 20936
rect 8300 20884 8352 20936
rect 9312 20884 9364 20936
rect 10784 20927 10836 20936
rect 10784 20893 10793 20927
rect 10793 20893 10827 20927
rect 10827 20893 10836 20927
rect 10784 20884 10836 20893
rect 13728 20884 13780 20936
rect 14832 20927 14884 20936
rect 14832 20893 14841 20927
rect 14841 20893 14875 20927
rect 14875 20893 14884 20927
rect 14832 20884 14884 20893
rect 14924 20884 14976 20936
rect 7840 20816 7892 20868
rect 8116 20816 8168 20868
rect 12992 20816 13044 20868
rect 13176 20816 13228 20868
rect 15016 20859 15068 20868
rect 15016 20825 15025 20859
rect 15025 20825 15059 20859
rect 15059 20825 15068 20859
rect 15016 20816 15068 20825
rect 16120 21020 16172 21072
rect 17224 21020 17276 21072
rect 19524 21020 19576 21072
rect 18052 20995 18104 21004
rect 18052 20961 18061 20995
rect 18061 20961 18095 20995
rect 18095 20961 18104 20995
rect 18052 20952 18104 20961
rect 16304 20927 16356 20936
rect 16304 20893 16318 20927
rect 16318 20893 16352 20927
rect 16352 20893 16356 20927
rect 18604 20952 18656 21004
rect 19800 21088 19852 21140
rect 24768 21088 24820 21140
rect 25044 21088 25096 21140
rect 30748 21131 30800 21140
rect 30748 21097 30757 21131
rect 30757 21097 30791 21131
rect 30791 21097 30800 21131
rect 30748 21088 30800 21097
rect 16304 20884 16356 20893
rect 16120 20859 16172 20868
rect 6460 20791 6512 20800
rect 6460 20757 6469 20791
rect 6469 20757 6503 20791
rect 6503 20757 6512 20791
rect 6460 20748 6512 20757
rect 16120 20825 16129 20859
rect 16129 20825 16163 20859
rect 16163 20825 16172 20859
rect 16120 20816 16172 20825
rect 18328 20884 18380 20936
rect 18144 20859 18196 20868
rect 18144 20825 18153 20859
rect 18153 20825 18187 20859
rect 18187 20825 18196 20859
rect 18144 20816 18196 20825
rect 16488 20791 16540 20800
rect 16488 20757 16497 20791
rect 16497 20757 16531 20791
rect 16531 20757 16540 20791
rect 16488 20748 16540 20757
rect 18420 20748 18472 20800
rect 19432 20927 19484 20936
rect 19432 20893 19439 20927
rect 19439 20893 19484 20927
rect 19432 20884 19484 20893
rect 19892 20884 19944 20936
rect 20076 20884 20128 20936
rect 20352 20884 20404 20936
rect 21364 20952 21416 21004
rect 20904 20927 20956 20936
rect 20904 20893 20913 20927
rect 20913 20893 20947 20927
rect 20947 20893 20956 20927
rect 20904 20884 20956 20893
rect 19432 20748 19484 20800
rect 20444 20816 20496 20868
rect 20628 20816 20680 20868
rect 20812 20859 20864 20868
rect 20812 20825 20821 20859
rect 20821 20825 20855 20859
rect 20855 20825 20864 20859
rect 20812 20816 20864 20825
rect 20260 20748 20312 20800
rect 21640 20927 21692 20936
rect 21640 20893 21677 20927
rect 21677 20893 21692 20927
rect 21640 20884 21692 20893
rect 21824 20927 21876 20936
rect 21824 20893 21833 20927
rect 21833 20893 21867 20927
rect 21867 20893 21876 20927
rect 21824 20884 21876 20893
rect 22836 21020 22888 21072
rect 24216 21020 24268 21072
rect 27620 21020 27672 21072
rect 28816 21020 28868 21072
rect 31668 21088 31720 21140
rect 31760 21088 31812 21140
rect 34612 21088 34664 21140
rect 35348 21088 35400 21140
rect 42984 21088 43036 21140
rect 45652 21088 45704 21140
rect 48412 21131 48464 21140
rect 48412 21097 48421 21131
rect 48421 21097 48455 21131
rect 48455 21097 48464 21131
rect 48412 21088 48464 21097
rect 49700 21088 49752 21140
rect 51724 21088 51776 21140
rect 45284 21020 45336 21072
rect 53748 21088 53800 21140
rect 46480 20952 46532 21004
rect 23572 20884 23624 20936
rect 24676 20927 24728 20936
rect 24676 20893 24685 20927
rect 24685 20893 24719 20927
rect 24719 20893 24728 20927
rect 24676 20884 24728 20893
rect 25412 20884 25464 20936
rect 25688 20927 25740 20936
rect 25688 20893 25697 20927
rect 25697 20893 25731 20927
rect 25731 20893 25740 20927
rect 25688 20884 25740 20893
rect 22376 20816 22428 20868
rect 25964 20859 26016 20868
rect 25964 20825 25973 20859
rect 25973 20825 26007 20859
rect 26007 20825 26016 20859
rect 25964 20816 26016 20825
rect 26516 20884 26568 20936
rect 27528 20927 27580 20936
rect 27528 20893 27537 20927
rect 27537 20893 27571 20927
rect 27571 20893 27580 20927
rect 27528 20884 27580 20893
rect 27344 20816 27396 20868
rect 21732 20748 21784 20800
rect 25320 20748 25372 20800
rect 26240 20748 26292 20800
rect 28080 20884 28132 20936
rect 29552 20927 29604 20936
rect 29552 20893 29561 20927
rect 29561 20893 29595 20927
rect 29595 20893 29604 20927
rect 29552 20884 29604 20893
rect 29644 20927 29696 20936
rect 29644 20893 29653 20927
rect 29653 20893 29687 20927
rect 29687 20893 29696 20927
rect 29828 20927 29880 20936
rect 29644 20884 29696 20893
rect 29828 20893 29837 20927
rect 29837 20893 29871 20927
rect 29871 20893 29880 20927
rect 29828 20884 29880 20893
rect 28816 20816 28868 20868
rect 30380 20884 30432 20936
rect 30840 20927 30892 20936
rect 30840 20893 30849 20927
rect 30849 20893 30883 20927
rect 30883 20893 30892 20927
rect 30840 20884 30892 20893
rect 31760 20927 31812 20936
rect 31760 20893 31769 20927
rect 31769 20893 31803 20927
rect 31803 20893 31812 20927
rect 31760 20884 31812 20893
rect 34796 20884 34848 20936
rect 37004 20927 37056 20936
rect 37004 20893 37013 20927
rect 37013 20893 37047 20927
rect 37047 20893 37056 20927
rect 37004 20884 37056 20893
rect 40224 20884 40276 20936
rect 41972 20927 42024 20936
rect 41972 20893 41981 20927
rect 41981 20893 42015 20927
rect 42015 20893 42024 20927
rect 41972 20884 42024 20893
rect 42156 20927 42208 20936
rect 42156 20893 42165 20927
rect 42165 20893 42199 20927
rect 42199 20893 42208 20927
rect 42156 20884 42208 20893
rect 43444 20927 43496 20936
rect 43444 20893 43453 20927
rect 43453 20893 43487 20927
rect 43487 20893 43496 20927
rect 43444 20884 43496 20893
rect 43628 20927 43680 20936
rect 43628 20893 43637 20927
rect 43637 20893 43671 20927
rect 43671 20893 43680 20927
rect 43628 20884 43680 20893
rect 45008 20927 45060 20936
rect 32680 20816 32732 20868
rect 34520 20816 34572 20868
rect 34888 20859 34940 20868
rect 34888 20825 34897 20859
rect 34897 20825 34931 20859
rect 34931 20825 34940 20859
rect 34888 20816 34940 20825
rect 40500 20859 40552 20868
rect 40500 20825 40509 20859
rect 40509 20825 40543 20859
rect 40543 20825 40552 20859
rect 40500 20816 40552 20825
rect 43996 20859 44048 20868
rect 43996 20825 44005 20859
rect 44005 20825 44039 20859
rect 44039 20825 44048 20859
rect 43996 20816 44048 20825
rect 45008 20893 45017 20927
rect 45017 20893 45051 20927
rect 45051 20893 45060 20927
rect 45008 20884 45060 20893
rect 45284 20927 45336 20936
rect 45284 20893 45293 20927
rect 45293 20893 45327 20927
rect 45327 20893 45336 20927
rect 45284 20884 45336 20893
rect 48320 20927 48372 20936
rect 48320 20893 48329 20927
rect 48329 20893 48363 20927
rect 48363 20893 48372 20927
rect 48320 20884 48372 20893
rect 51080 20995 51132 21004
rect 49240 20927 49292 20936
rect 49240 20893 49249 20927
rect 49249 20893 49283 20927
rect 49283 20893 49292 20927
rect 49240 20884 49292 20893
rect 51080 20961 51089 20995
rect 51089 20961 51123 20995
rect 51123 20961 51132 20995
rect 51080 20952 51132 20961
rect 51724 20952 51776 21004
rect 51356 20927 51408 20936
rect 47492 20816 47544 20868
rect 51356 20893 51365 20927
rect 51365 20893 51399 20927
rect 51399 20893 51408 20927
rect 51356 20884 51408 20893
rect 52000 20927 52052 20936
rect 52000 20893 52009 20927
rect 52009 20893 52043 20927
rect 52043 20893 52052 20927
rect 52000 20884 52052 20893
rect 56324 21020 56376 21072
rect 56692 21020 56744 21072
rect 54116 20995 54168 21004
rect 54116 20961 54125 20995
rect 54125 20961 54159 20995
rect 54159 20961 54168 20995
rect 54116 20952 54168 20961
rect 54392 20952 54444 21004
rect 54208 20927 54260 20936
rect 54208 20893 54217 20927
rect 54217 20893 54251 20927
rect 54251 20893 54260 20927
rect 55680 20927 55732 20936
rect 54208 20884 54260 20893
rect 55680 20893 55689 20927
rect 55689 20893 55723 20927
rect 55723 20893 55732 20927
rect 55680 20884 55732 20893
rect 56232 20884 56284 20936
rect 56784 20927 56836 20936
rect 56784 20893 56792 20927
rect 56792 20893 56826 20927
rect 56826 20893 56836 20927
rect 56784 20884 56836 20893
rect 57704 20952 57756 21004
rect 58164 20927 58216 20936
rect 58164 20893 58173 20927
rect 58173 20893 58207 20927
rect 58207 20893 58216 20927
rect 58164 20884 58216 20893
rect 55496 20859 55548 20868
rect 55496 20825 55505 20859
rect 55505 20825 55539 20859
rect 55539 20825 55548 20859
rect 56600 20859 56652 20868
rect 55496 20816 55548 20825
rect 37372 20791 37424 20800
rect 37372 20757 37381 20791
rect 37381 20757 37415 20791
rect 37415 20757 37424 20791
rect 37372 20748 37424 20757
rect 45100 20791 45152 20800
rect 45100 20757 45109 20791
rect 45109 20757 45143 20791
rect 45143 20757 45152 20791
rect 45100 20748 45152 20757
rect 56232 20791 56284 20800
rect 56232 20757 56241 20791
rect 56241 20757 56275 20791
rect 56275 20757 56284 20791
rect 56232 20748 56284 20757
rect 56600 20825 56609 20859
rect 56609 20825 56643 20859
rect 56643 20825 56652 20859
rect 56600 20816 56652 20825
rect 56692 20816 56744 20868
rect 56968 20816 57020 20868
rect 19574 20646 19626 20698
rect 19638 20646 19690 20698
rect 19702 20646 19754 20698
rect 19766 20646 19818 20698
rect 19830 20646 19882 20698
rect 50294 20646 50346 20698
rect 50358 20646 50410 20698
rect 50422 20646 50474 20698
rect 50486 20646 50538 20698
rect 50550 20646 50602 20698
rect 1492 20476 1544 20528
rect 2228 20476 2280 20528
rect 5264 20587 5316 20596
rect 5264 20553 5273 20587
rect 5273 20553 5307 20587
rect 5307 20553 5316 20587
rect 5264 20544 5316 20553
rect 7472 20544 7524 20596
rect 8208 20544 8260 20596
rect 14648 20587 14700 20596
rect 14648 20553 14657 20587
rect 14657 20553 14691 20587
rect 14691 20553 14700 20587
rect 14648 20544 14700 20553
rect 18236 20544 18288 20596
rect 19064 20544 19116 20596
rect 19156 20544 19208 20596
rect 21732 20544 21784 20596
rect 21916 20544 21968 20596
rect 22376 20544 22428 20596
rect 24308 20544 24360 20596
rect 26516 20544 26568 20596
rect 29644 20544 29696 20596
rect 31760 20544 31812 20596
rect 34888 20544 34940 20596
rect 41972 20544 42024 20596
rect 47492 20544 47544 20596
rect 51816 20587 51868 20596
rect 51816 20553 51825 20587
rect 51825 20553 51859 20587
rect 51859 20553 51868 20587
rect 51816 20544 51868 20553
rect 57060 20544 57112 20596
rect 10416 20519 10468 20528
rect 2136 20451 2188 20460
rect 2136 20417 2145 20451
rect 2145 20417 2179 20451
rect 2179 20417 2188 20451
rect 10416 20485 10425 20519
rect 10425 20485 10459 20519
rect 10459 20485 10468 20519
rect 10416 20476 10468 20485
rect 13820 20476 13872 20528
rect 2136 20408 2188 20417
rect 2504 20451 2556 20460
rect 2504 20417 2513 20451
rect 2513 20417 2547 20451
rect 2547 20417 2556 20451
rect 2504 20408 2556 20417
rect 6460 20408 6512 20460
rect 7840 20451 7892 20460
rect 7840 20417 7849 20451
rect 7849 20417 7883 20451
rect 7883 20417 7892 20451
rect 7840 20408 7892 20417
rect 8024 20408 8076 20460
rect 9496 20408 9548 20460
rect 9956 20451 10008 20460
rect 9956 20417 9965 20451
rect 9965 20417 9999 20451
rect 9999 20417 10008 20451
rect 9956 20408 10008 20417
rect 10324 20408 10376 20460
rect 12624 20408 12676 20460
rect 13360 20451 13412 20460
rect 13360 20417 13369 20451
rect 13369 20417 13403 20451
rect 13403 20417 13412 20451
rect 13360 20408 13412 20417
rect 3976 20383 4028 20392
rect 3976 20349 3985 20383
rect 3985 20349 4019 20383
rect 4019 20349 4028 20383
rect 3976 20340 4028 20349
rect 4068 20272 4120 20324
rect 1952 20204 2004 20256
rect 4896 20204 4948 20256
rect 9680 20272 9732 20324
rect 13084 20315 13136 20324
rect 13084 20281 13093 20315
rect 13093 20281 13127 20315
rect 13127 20281 13136 20315
rect 13084 20272 13136 20281
rect 13728 20451 13780 20460
rect 13728 20417 13737 20451
rect 13737 20417 13771 20451
rect 13771 20417 13780 20451
rect 18328 20476 18380 20528
rect 24216 20476 24268 20528
rect 25320 20519 25372 20528
rect 25320 20485 25329 20519
rect 25329 20485 25363 20519
rect 25363 20485 25372 20519
rect 25320 20476 25372 20485
rect 25688 20476 25740 20528
rect 27344 20476 27396 20528
rect 13728 20408 13780 20417
rect 18604 20408 18656 20460
rect 19984 20408 20036 20460
rect 20444 20408 20496 20460
rect 18420 20340 18472 20392
rect 29000 20519 29052 20528
rect 29000 20485 29025 20519
rect 29025 20485 29052 20519
rect 29000 20476 29052 20485
rect 29644 20451 29696 20460
rect 29644 20417 29653 20451
rect 29653 20417 29687 20451
rect 29687 20417 29696 20451
rect 29644 20408 29696 20417
rect 30104 20408 30156 20460
rect 30748 20408 30800 20460
rect 30380 20383 30432 20392
rect 13636 20272 13688 20324
rect 15200 20272 15252 20324
rect 18144 20272 18196 20324
rect 19156 20272 19208 20324
rect 29552 20272 29604 20324
rect 30380 20349 30389 20383
rect 30389 20349 30423 20383
rect 30423 20349 30432 20383
rect 30380 20340 30432 20349
rect 30840 20340 30892 20392
rect 33416 20476 33468 20528
rect 42156 20476 42208 20528
rect 33508 20451 33560 20460
rect 33508 20417 33517 20451
rect 33517 20417 33551 20451
rect 33551 20417 33560 20451
rect 33508 20408 33560 20417
rect 34520 20408 34572 20460
rect 34704 20451 34756 20460
rect 34704 20417 34713 20451
rect 34713 20417 34747 20451
rect 34747 20417 34756 20451
rect 34704 20408 34756 20417
rect 37372 20408 37424 20460
rect 38292 20408 38344 20460
rect 40500 20451 40552 20460
rect 40500 20417 40509 20451
rect 40509 20417 40543 20451
rect 40543 20417 40552 20451
rect 40500 20408 40552 20417
rect 43352 20451 43404 20460
rect 34796 20340 34848 20392
rect 38476 20383 38528 20392
rect 38476 20349 38485 20383
rect 38485 20349 38519 20383
rect 38519 20349 38528 20383
rect 38476 20340 38528 20349
rect 39764 20340 39816 20392
rect 31760 20272 31812 20324
rect 43352 20417 43361 20451
rect 43361 20417 43395 20451
rect 43395 20417 43404 20451
rect 43352 20408 43404 20417
rect 43996 20408 44048 20460
rect 45008 20476 45060 20528
rect 57244 20519 57296 20528
rect 57244 20485 57253 20519
rect 57253 20485 57287 20519
rect 57287 20485 57296 20519
rect 57244 20476 57296 20485
rect 58164 20519 58216 20528
rect 58164 20485 58173 20519
rect 58173 20485 58207 20519
rect 58207 20485 58216 20519
rect 58164 20476 58216 20485
rect 45100 20451 45152 20460
rect 45100 20417 45109 20451
rect 45109 20417 45143 20451
rect 45143 20417 45152 20451
rect 45100 20408 45152 20417
rect 45284 20408 45336 20460
rect 51080 20408 51132 20460
rect 51356 20451 51408 20460
rect 51356 20417 51365 20451
rect 51365 20417 51399 20451
rect 51399 20417 51408 20451
rect 51356 20408 51408 20417
rect 43444 20383 43496 20392
rect 43444 20349 43453 20383
rect 43453 20349 43487 20383
rect 43487 20349 43496 20383
rect 43444 20340 43496 20349
rect 51724 20408 51776 20460
rect 56968 20451 57020 20460
rect 56968 20417 56977 20451
rect 56977 20417 57011 20451
rect 57011 20417 57020 20451
rect 56968 20408 57020 20417
rect 52000 20340 52052 20392
rect 41972 20272 42024 20324
rect 45836 20272 45888 20324
rect 11152 20204 11204 20256
rect 13544 20204 13596 20256
rect 15752 20247 15804 20256
rect 15752 20213 15761 20247
rect 15761 20213 15795 20247
rect 15795 20213 15804 20247
rect 15752 20204 15804 20213
rect 18328 20204 18380 20256
rect 25964 20247 26016 20256
rect 25964 20213 25973 20247
rect 25973 20213 26007 20247
rect 26007 20213 26016 20247
rect 25964 20204 26016 20213
rect 26056 20204 26108 20256
rect 27712 20204 27764 20256
rect 28264 20204 28316 20256
rect 29092 20204 29144 20256
rect 29736 20204 29788 20256
rect 30380 20204 30432 20256
rect 39764 20247 39816 20256
rect 39764 20213 39773 20247
rect 39773 20213 39807 20247
rect 39807 20213 39816 20247
rect 39764 20204 39816 20213
rect 43628 20204 43680 20256
rect 54024 20204 54076 20256
rect 4214 20102 4266 20154
rect 4278 20102 4330 20154
rect 4342 20102 4394 20154
rect 4406 20102 4458 20154
rect 4470 20102 4522 20154
rect 34934 20102 34986 20154
rect 34998 20102 35050 20154
rect 35062 20102 35114 20154
rect 35126 20102 35178 20154
rect 35190 20102 35242 20154
rect 3976 20000 4028 20052
rect 5448 20000 5500 20052
rect 8208 20043 8260 20052
rect 2872 19771 2924 19780
rect 2872 19737 2881 19771
rect 2881 19737 2915 19771
rect 2915 19737 2924 19771
rect 2872 19728 2924 19737
rect 5264 19864 5316 19916
rect 4068 19796 4120 19848
rect 5540 19839 5592 19848
rect 5540 19805 5549 19839
rect 5549 19805 5583 19839
rect 5583 19805 5592 19839
rect 8208 20009 8217 20043
rect 8217 20009 8251 20043
rect 8251 20009 8260 20043
rect 8208 20000 8260 20009
rect 6920 19932 6972 19984
rect 8116 19932 8168 19984
rect 12992 20000 13044 20052
rect 13544 20043 13596 20052
rect 13544 20009 13553 20043
rect 13553 20009 13587 20043
rect 13587 20009 13596 20043
rect 13544 20000 13596 20009
rect 14648 20000 14700 20052
rect 16764 20000 16816 20052
rect 26056 20000 26108 20052
rect 26516 20000 26568 20052
rect 11152 19907 11204 19916
rect 7104 19839 7156 19848
rect 5540 19796 5592 19805
rect 7104 19805 7113 19839
rect 7113 19805 7147 19839
rect 7147 19805 7156 19839
rect 7104 19796 7156 19805
rect 11152 19873 11161 19907
rect 11161 19873 11195 19907
rect 11195 19873 11204 19907
rect 11152 19864 11204 19873
rect 11980 19907 12032 19916
rect 11980 19873 11989 19907
rect 11989 19873 12023 19907
rect 12023 19873 12032 19907
rect 11980 19864 12032 19873
rect 7840 19796 7892 19848
rect 9680 19839 9732 19848
rect 8024 19771 8076 19780
rect 8024 19737 8033 19771
rect 8033 19737 8067 19771
rect 8067 19737 8076 19771
rect 8024 19728 8076 19737
rect 9680 19805 9689 19839
rect 9689 19805 9723 19839
rect 9723 19805 9732 19839
rect 9680 19796 9732 19805
rect 9496 19771 9548 19780
rect 9496 19737 9505 19771
rect 9505 19737 9539 19771
rect 9539 19737 9548 19771
rect 9496 19728 9548 19737
rect 10232 19728 10284 19780
rect 13636 19728 13688 19780
rect 6276 19703 6328 19712
rect 6276 19669 6285 19703
rect 6285 19669 6319 19703
rect 6319 19669 6328 19703
rect 6276 19660 6328 19669
rect 7840 19660 7892 19712
rect 14188 19703 14240 19712
rect 14188 19669 14197 19703
rect 14197 19669 14231 19703
rect 14231 19669 14240 19703
rect 14188 19660 14240 19669
rect 20076 19932 20128 19984
rect 19984 19864 20036 19916
rect 34520 20000 34572 20052
rect 42800 20000 42852 20052
rect 54208 20000 54260 20052
rect 54392 20043 54444 20052
rect 54392 20009 54401 20043
rect 54401 20009 54435 20043
rect 54435 20009 54444 20043
rect 54392 20000 54444 20009
rect 18696 19796 18748 19848
rect 16028 19771 16080 19780
rect 16028 19737 16037 19771
rect 16037 19737 16071 19771
rect 16071 19737 16080 19771
rect 16028 19728 16080 19737
rect 17776 19728 17828 19780
rect 18236 19660 18288 19712
rect 19248 19728 19300 19780
rect 26332 19796 26384 19848
rect 26516 19796 26568 19848
rect 27160 19839 27212 19848
rect 27160 19805 27169 19839
rect 27169 19805 27203 19839
rect 27203 19805 27212 19839
rect 27160 19796 27212 19805
rect 28080 19839 28132 19848
rect 28080 19805 28089 19839
rect 28089 19805 28123 19839
rect 28123 19805 28132 19839
rect 28080 19796 28132 19805
rect 29000 19864 29052 19916
rect 30840 19907 30892 19916
rect 30840 19873 30849 19907
rect 30849 19873 30883 19907
rect 30883 19873 30892 19907
rect 30840 19864 30892 19873
rect 39764 19932 39816 19984
rect 33508 19864 33560 19916
rect 38292 19907 38344 19916
rect 28264 19839 28316 19848
rect 28264 19805 28273 19839
rect 28273 19805 28307 19839
rect 28307 19805 28316 19839
rect 28264 19796 28316 19805
rect 28816 19796 28868 19848
rect 38292 19873 38301 19907
rect 38301 19873 38335 19907
rect 38335 19873 38344 19907
rect 38292 19864 38344 19873
rect 43444 19864 43496 19916
rect 46940 19864 46992 19916
rect 48320 19864 48372 19916
rect 48964 19864 49016 19916
rect 20904 19728 20956 19780
rect 25964 19728 26016 19780
rect 28172 19771 28224 19780
rect 20076 19660 20128 19712
rect 20996 19660 21048 19712
rect 22192 19660 22244 19712
rect 23204 19703 23256 19712
rect 23204 19669 23213 19703
rect 23213 19669 23247 19703
rect 23247 19669 23256 19703
rect 23204 19660 23256 19669
rect 28172 19737 28181 19771
rect 28181 19737 28215 19771
rect 28215 19737 28224 19771
rect 28172 19728 28224 19737
rect 29644 19728 29696 19780
rect 31852 19728 31904 19780
rect 32864 19728 32916 19780
rect 33416 19728 33468 19780
rect 34796 19796 34848 19848
rect 35992 19839 36044 19848
rect 35992 19805 36001 19839
rect 36001 19805 36035 19839
rect 36035 19805 36044 19839
rect 35992 19796 36044 19805
rect 36176 19839 36228 19848
rect 36176 19805 36185 19839
rect 36185 19805 36219 19839
rect 36219 19805 36228 19839
rect 36176 19796 36228 19805
rect 38476 19839 38528 19848
rect 38476 19805 38485 19839
rect 38485 19805 38519 19839
rect 38519 19805 38528 19839
rect 38476 19796 38528 19805
rect 44180 19796 44232 19848
rect 29920 19660 29972 19712
rect 42708 19728 42760 19780
rect 47768 19796 47820 19848
rect 49884 19796 49936 19848
rect 50620 19796 50672 19848
rect 50712 19839 50764 19848
rect 50712 19805 50721 19839
rect 50721 19805 50755 19839
rect 50755 19805 50764 19839
rect 53472 19839 53524 19848
rect 50712 19796 50764 19805
rect 53472 19805 53481 19839
rect 53481 19805 53515 19839
rect 53515 19805 53524 19839
rect 53472 19796 53524 19805
rect 57336 19864 57388 19916
rect 53932 19796 53984 19848
rect 56692 19839 56744 19848
rect 56692 19805 56701 19839
rect 56701 19805 56735 19839
rect 56735 19805 56744 19839
rect 56692 19796 56744 19805
rect 56876 19839 56928 19848
rect 56876 19805 56885 19839
rect 56885 19805 56919 19839
rect 56919 19805 56928 19839
rect 56876 19796 56928 19805
rect 57152 19796 57204 19848
rect 50988 19728 51040 19780
rect 54668 19771 54720 19780
rect 38844 19660 38896 19712
rect 41788 19660 41840 19712
rect 48780 19660 48832 19712
rect 52000 19660 52052 19712
rect 53564 19703 53616 19712
rect 53564 19669 53573 19703
rect 53573 19669 53607 19703
rect 53607 19669 53616 19703
rect 54668 19737 54677 19771
rect 54677 19737 54711 19771
rect 54711 19737 54720 19771
rect 54668 19728 54720 19737
rect 56508 19703 56560 19712
rect 53564 19660 53616 19669
rect 56508 19669 56517 19703
rect 56517 19669 56551 19703
rect 56551 19669 56560 19703
rect 56508 19660 56560 19669
rect 19574 19558 19626 19610
rect 19638 19558 19690 19610
rect 19702 19558 19754 19610
rect 19766 19558 19818 19610
rect 19830 19558 19882 19610
rect 50294 19558 50346 19610
rect 50358 19558 50410 19610
rect 50422 19558 50474 19610
rect 50486 19558 50538 19610
rect 50550 19558 50602 19610
rect 2872 19456 2924 19508
rect 1400 19320 1452 19372
rect 5448 19456 5500 19508
rect 14372 19456 14424 19508
rect 18604 19456 18656 19508
rect 7748 19388 7800 19440
rect 9956 19388 10008 19440
rect 14188 19388 14240 19440
rect 15936 19431 15988 19440
rect 5540 19320 5592 19372
rect 6276 19320 6328 19372
rect 7196 19363 7248 19372
rect 7196 19329 7205 19363
rect 7205 19329 7239 19363
rect 7239 19329 7248 19363
rect 7196 19320 7248 19329
rect 7472 19363 7524 19372
rect 7472 19329 7481 19363
rect 7481 19329 7515 19363
rect 7515 19329 7524 19363
rect 7472 19320 7524 19329
rect 8024 19320 8076 19372
rect 13636 19363 13688 19372
rect 13636 19329 13645 19363
rect 13645 19329 13679 19363
rect 13679 19329 13688 19363
rect 13636 19320 13688 19329
rect 14648 19363 14700 19372
rect 14648 19329 14657 19363
rect 14657 19329 14691 19363
rect 14691 19329 14700 19363
rect 14648 19320 14700 19329
rect 14832 19363 14884 19372
rect 14832 19329 14841 19363
rect 14841 19329 14875 19363
rect 14875 19329 14884 19363
rect 14832 19320 14884 19329
rect 15936 19397 15945 19431
rect 15945 19397 15979 19431
rect 15979 19397 15988 19431
rect 15936 19388 15988 19397
rect 18052 19388 18104 19440
rect 18512 19431 18564 19440
rect 15200 19363 15252 19372
rect 15200 19329 15209 19363
rect 15209 19329 15243 19363
rect 15243 19329 15252 19363
rect 15200 19320 15252 19329
rect 3976 19252 4028 19304
rect 6920 19252 6972 19304
rect 7748 19295 7800 19304
rect 7748 19261 7757 19295
rect 7757 19261 7791 19295
rect 7791 19261 7800 19295
rect 7748 19252 7800 19261
rect 11152 19252 11204 19304
rect 13544 19295 13596 19304
rect 13544 19261 13553 19295
rect 13553 19261 13587 19295
rect 13587 19261 13596 19295
rect 13544 19252 13596 19261
rect 14740 19252 14792 19304
rect 16028 19320 16080 19372
rect 17776 19363 17828 19372
rect 17776 19329 17785 19363
rect 17785 19329 17819 19363
rect 17819 19329 17828 19363
rect 17776 19320 17828 19329
rect 18236 19363 18288 19372
rect 18236 19329 18245 19363
rect 18245 19329 18279 19363
rect 18279 19329 18288 19363
rect 18236 19320 18288 19329
rect 18512 19397 18521 19431
rect 18521 19397 18555 19431
rect 18555 19397 18564 19431
rect 18512 19388 18564 19397
rect 18696 19320 18748 19372
rect 18880 19456 18932 19508
rect 19156 19388 19208 19440
rect 19524 19363 19576 19372
rect 19524 19329 19533 19363
rect 19533 19329 19567 19363
rect 19567 19329 19576 19363
rect 19524 19320 19576 19329
rect 19984 19456 20036 19508
rect 21456 19388 21508 19440
rect 16212 19252 16264 19304
rect 16764 19295 16816 19304
rect 16764 19261 16773 19295
rect 16773 19261 16807 19295
rect 16807 19261 16816 19295
rect 16764 19252 16816 19261
rect 19708 19363 19760 19372
rect 19708 19329 19722 19363
rect 19722 19329 19756 19363
rect 19756 19329 19760 19363
rect 19708 19320 19760 19329
rect 19984 19252 20036 19304
rect 7656 19184 7708 19236
rect 10508 19184 10560 19236
rect 16396 19184 16448 19236
rect 21456 19252 21508 19304
rect 22376 19456 22428 19508
rect 23388 19456 23440 19508
rect 22100 19431 22152 19440
rect 22100 19397 22109 19431
rect 22109 19397 22143 19431
rect 22143 19397 22152 19431
rect 22100 19388 22152 19397
rect 22744 19388 22796 19440
rect 22192 19363 22244 19372
rect 22192 19329 22201 19363
rect 22201 19329 22235 19363
rect 22235 19329 22244 19363
rect 22192 19320 22244 19329
rect 21916 19184 21968 19236
rect 23020 19320 23072 19372
rect 23296 19363 23348 19372
rect 23296 19329 23305 19363
rect 23305 19329 23339 19363
rect 23339 19329 23348 19363
rect 23480 19363 23532 19372
rect 23296 19320 23348 19329
rect 23480 19329 23489 19363
rect 23489 19329 23523 19363
rect 23523 19329 23532 19363
rect 23480 19320 23532 19329
rect 24952 19456 25004 19508
rect 28080 19456 28132 19508
rect 29736 19456 29788 19508
rect 32680 19499 32732 19508
rect 32680 19465 32689 19499
rect 32689 19465 32723 19499
rect 32723 19465 32732 19499
rect 32680 19456 32732 19465
rect 34796 19456 34848 19508
rect 44180 19499 44232 19508
rect 44180 19465 44189 19499
rect 44189 19465 44223 19499
rect 44223 19465 44232 19499
rect 44180 19456 44232 19465
rect 50620 19456 50672 19508
rect 24676 19388 24728 19440
rect 29000 19388 29052 19440
rect 35992 19388 36044 19440
rect 24492 19320 24544 19372
rect 24768 19320 24820 19372
rect 31760 19320 31812 19372
rect 34336 19363 34388 19372
rect 23112 19252 23164 19304
rect 24308 19252 24360 19304
rect 26240 19252 26292 19304
rect 31024 19252 31076 19304
rect 32312 19295 32364 19304
rect 32312 19261 32321 19295
rect 32321 19261 32355 19295
rect 32355 19261 32364 19295
rect 32312 19252 32364 19261
rect 29000 19184 29052 19236
rect 31392 19184 31444 19236
rect 2688 19116 2740 19168
rect 4068 19159 4120 19168
rect 4068 19125 4077 19159
rect 4077 19125 4111 19159
rect 4111 19125 4120 19159
rect 4068 19116 4120 19125
rect 12992 19116 13044 19168
rect 16120 19116 16172 19168
rect 16488 19116 16540 19168
rect 18144 19116 18196 19168
rect 23388 19116 23440 19168
rect 29460 19116 29512 19168
rect 31484 19159 31536 19168
rect 31484 19125 31493 19159
rect 31493 19125 31527 19159
rect 31527 19125 31536 19159
rect 31484 19116 31536 19125
rect 31760 19116 31812 19168
rect 34336 19329 34345 19363
rect 34345 19329 34379 19363
rect 34379 19329 34388 19363
rect 34336 19320 34388 19329
rect 36176 19320 36228 19372
rect 37004 19320 37056 19372
rect 37188 19320 37240 19372
rect 42708 19320 42760 19372
rect 38016 19295 38068 19304
rect 38016 19261 38025 19295
rect 38025 19261 38059 19295
rect 38059 19261 38068 19295
rect 38016 19252 38068 19261
rect 42800 19295 42852 19304
rect 42800 19261 42809 19295
rect 42809 19261 42843 19295
rect 42843 19261 42852 19295
rect 43996 19363 44048 19372
rect 43996 19329 44005 19363
rect 44005 19329 44039 19363
rect 44039 19329 44048 19363
rect 43996 19320 44048 19329
rect 42800 19252 42852 19261
rect 45100 19252 45152 19304
rect 46020 19320 46072 19372
rect 46940 19320 46992 19372
rect 47768 19363 47820 19372
rect 47768 19329 47777 19363
rect 47777 19329 47811 19363
rect 47811 19329 47820 19363
rect 47768 19320 47820 19329
rect 50988 19456 51040 19508
rect 56232 19456 56284 19508
rect 57244 19456 57296 19508
rect 48780 19363 48832 19372
rect 48780 19329 48789 19363
rect 48789 19329 48823 19363
rect 48823 19329 48832 19363
rect 48780 19320 48832 19329
rect 48964 19363 49016 19372
rect 48964 19329 48973 19363
rect 48973 19329 49007 19363
rect 49007 19329 49016 19363
rect 48964 19320 49016 19329
rect 49516 19363 49568 19372
rect 49516 19329 49525 19363
rect 49525 19329 49559 19363
rect 49559 19329 49568 19363
rect 49700 19363 49752 19372
rect 49516 19320 49568 19329
rect 49700 19329 49709 19363
rect 49709 19329 49743 19363
rect 49743 19329 49752 19363
rect 49700 19320 49752 19329
rect 50160 19320 50212 19372
rect 50436 19363 50488 19372
rect 50436 19329 50445 19363
rect 50445 19329 50479 19363
rect 50479 19329 50488 19363
rect 50436 19320 50488 19329
rect 56600 19388 56652 19440
rect 53472 19320 53524 19372
rect 54668 19320 54720 19372
rect 56876 19320 56928 19372
rect 57888 19320 57940 19372
rect 49608 19252 49660 19304
rect 50620 19252 50672 19304
rect 52736 19252 52788 19304
rect 53564 19295 53616 19304
rect 53564 19261 53573 19295
rect 53573 19261 53607 19295
rect 53607 19261 53616 19295
rect 53564 19252 53616 19261
rect 53932 19295 53984 19304
rect 53932 19261 53941 19295
rect 53941 19261 53975 19295
rect 53975 19261 53984 19295
rect 53932 19252 53984 19261
rect 49884 19184 49936 19236
rect 40316 19116 40368 19168
rect 41788 19159 41840 19168
rect 41788 19125 41797 19159
rect 41797 19125 41831 19159
rect 41831 19125 41840 19159
rect 41788 19116 41840 19125
rect 50712 19116 50764 19168
rect 51724 19159 51776 19168
rect 51724 19125 51733 19159
rect 51733 19125 51767 19159
rect 51767 19125 51776 19159
rect 51724 19116 51776 19125
rect 56600 19116 56652 19168
rect 57152 19159 57204 19168
rect 57152 19125 57161 19159
rect 57161 19125 57195 19159
rect 57195 19125 57204 19159
rect 57152 19116 57204 19125
rect 57704 19116 57756 19168
rect 4214 19014 4266 19066
rect 4278 19014 4330 19066
rect 4342 19014 4394 19066
rect 4406 19014 4458 19066
rect 4470 19014 4522 19066
rect 34934 19014 34986 19066
rect 34998 19014 35050 19066
rect 35062 19014 35114 19066
rect 35126 19014 35178 19066
rect 35190 19014 35242 19066
rect 1400 18955 1452 18964
rect 1400 18921 1409 18955
rect 1409 18921 1443 18955
rect 1443 18921 1452 18955
rect 1400 18912 1452 18921
rect 4068 18912 4120 18964
rect 7748 18912 7800 18964
rect 11060 18912 11112 18964
rect 10508 18844 10560 18896
rect 17868 18912 17920 18964
rect 18052 18955 18104 18964
rect 18052 18921 18061 18955
rect 18061 18921 18095 18955
rect 18095 18921 18104 18955
rect 18052 18912 18104 18921
rect 19708 18912 19760 18964
rect 20628 18912 20680 18964
rect 22376 18912 22428 18964
rect 23480 18912 23532 18964
rect 27160 18912 27212 18964
rect 29000 18955 29052 18964
rect 29000 18921 29009 18955
rect 29009 18921 29043 18955
rect 29043 18921 29052 18955
rect 29000 18912 29052 18921
rect 30656 18912 30708 18964
rect 31024 18955 31076 18964
rect 31024 18921 31033 18955
rect 31033 18921 31067 18955
rect 31067 18921 31076 18955
rect 31024 18912 31076 18921
rect 32864 18955 32916 18964
rect 32864 18921 32873 18955
rect 32873 18921 32907 18955
rect 32907 18921 32916 18955
rect 32864 18912 32916 18921
rect 34704 18912 34756 18964
rect 43996 18912 44048 18964
rect 49516 18912 49568 18964
rect 50436 18912 50488 18964
rect 51724 18912 51776 18964
rect 53196 18912 53248 18964
rect 53472 18912 53524 18964
rect 1584 18708 1636 18760
rect 4068 18708 4120 18760
rect 4896 18751 4948 18760
rect 4896 18717 4905 18751
rect 4905 18717 4939 18751
rect 4939 18717 4948 18751
rect 4896 18708 4948 18717
rect 7196 18751 7248 18760
rect 7196 18717 7205 18751
rect 7205 18717 7239 18751
rect 7239 18717 7248 18751
rect 7196 18708 7248 18717
rect 7472 18776 7524 18828
rect 8024 18776 8076 18828
rect 7564 18751 7616 18760
rect 7564 18717 7573 18751
rect 7573 18717 7607 18751
rect 7607 18717 7616 18751
rect 7564 18708 7616 18717
rect 4988 18640 5040 18692
rect 6276 18640 6328 18692
rect 13544 18819 13596 18828
rect 11060 18708 11112 18760
rect 8668 18572 8720 18624
rect 13544 18785 13553 18819
rect 13553 18785 13587 18819
rect 13587 18785 13596 18819
rect 13544 18776 13596 18785
rect 15200 18819 15252 18828
rect 15200 18785 15209 18819
rect 15209 18785 15243 18819
rect 15243 18785 15252 18819
rect 15200 18776 15252 18785
rect 14372 18751 14424 18760
rect 14372 18717 14381 18751
rect 14381 18717 14415 18751
rect 14415 18717 14424 18751
rect 14372 18708 14424 18717
rect 14924 18751 14976 18760
rect 14924 18717 14933 18751
rect 14933 18717 14967 18751
rect 14967 18717 14976 18751
rect 14924 18708 14976 18717
rect 15292 18751 15344 18760
rect 15292 18717 15301 18751
rect 15301 18717 15335 18751
rect 15335 18717 15344 18751
rect 15292 18708 15344 18717
rect 16212 18751 16264 18760
rect 14740 18640 14792 18692
rect 16212 18717 16221 18751
rect 16221 18717 16255 18751
rect 16255 18717 16264 18751
rect 16212 18708 16264 18717
rect 20720 18844 20772 18896
rect 21272 18844 21324 18896
rect 27620 18887 27672 18896
rect 21456 18776 21508 18828
rect 17868 18708 17920 18760
rect 19248 18751 19300 18760
rect 16120 18640 16172 18692
rect 16948 18640 17000 18692
rect 17776 18640 17828 18692
rect 19248 18717 19257 18751
rect 19257 18717 19291 18751
rect 19291 18717 19300 18751
rect 19248 18708 19300 18717
rect 18880 18640 18932 18692
rect 20812 18708 20864 18760
rect 21732 18708 21784 18760
rect 22100 18776 22152 18828
rect 23204 18708 23256 18760
rect 25688 18751 25740 18760
rect 21364 18640 21416 18692
rect 21824 18683 21876 18692
rect 21824 18649 21833 18683
rect 21833 18649 21867 18683
rect 21867 18649 21876 18683
rect 21824 18640 21876 18649
rect 12808 18572 12860 18624
rect 17960 18572 18012 18624
rect 18144 18572 18196 18624
rect 24216 18640 24268 18692
rect 24492 18572 24544 18624
rect 25688 18717 25697 18751
rect 25697 18717 25731 18751
rect 25731 18717 25740 18751
rect 25688 18708 25740 18717
rect 26424 18708 26476 18760
rect 27620 18853 27629 18887
rect 27629 18853 27663 18887
rect 27663 18853 27672 18887
rect 27620 18844 27672 18853
rect 27712 18844 27764 18896
rect 31208 18844 31260 18896
rect 31484 18844 31536 18896
rect 34520 18844 34572 18896
rect 35992 18844 36044 18896
rect 42800 18844 42852 18896
rect 27804 18776 27856 18828
rect 40316 18819 40368 18828
rect 27712 18708 27764 18760
rect 29184 18708 29236 18760
rect 29736 18751 29788 18760
rect 29736 18717 29745 18751
rect 29745 18717 29779 18751
rect 29779 18717 29788 18751
rect 29736 18708 29788 18717
rect 29920 18751 29972 18760
rect 29920 18717 29929 18751
rect 29929 18717 29963 18751
rect 29963 18717 29972 18751
rect 29920 18708 29972 18717
rect 30104 18751 30156 18760
rect 30104 18717 30113 18751
rect 30113 18717 30147 18751
rect 30147 18717 30156 18751
rect 30104 18708 30156 18717
rect 30196 18708 30248 18760
rect 27528 18640 27580 18692
rect 27620 18640 27672 18692
rect 29644 18640 29696 18692
rect 29368 18572 29420 18624
rect 31392 18640 31444 18692
rect 31852 18751 31904 18760
rect 31852 18717 31861 18751
rect 31861 18717 31895 18751
rect 31895 18717 31904 18751
rect 33600 18751 33652 18760
rect 31852 18708 31904 18717
rect 33600 18717 33609 18751
rect 33609 18717 33643 18751
rect 33643 18717 33652 18751
rect 33600 18708 33652 18717
rect 32312 18640 32364 18692
rect 33968 18751 34020 18760
rect 33968 18717 33977 18751
rect 33977 18717 34011 18751
rect 34011 18717 34020 18751
rect 33968 18708 34020 18717
rect 35716 18708 35768 18760
rect 36360 18708 36412 18760
rect 40316 18785 40325 18819
rect 40325 18785 40359 18819
rect 40359 18785 40368 18819
rect 40316 18776 40368 18785
rect 40684 18708 40736 18760
rect 41696 18751 41748 18760
rect 41696 18717 41705 18751
rect 41705 18717 41739 18751
rect 41739 18717 41748 18751
rect 41696 18708 41748 18717
rect 49608 18776 49660 18828
rect 45100 18708 45152 18760
rect 46020 18751 46072 18760
rect 46020 18717 46029 18751
rect 46029 18717 46063 18751
rect 46063 18717 46072 18751
rect 46020 18708 46072 18717
rect 50160 18751 50212 18760
rect 50160 18717 50169 18751
rect 50169 18717 50203 18751
rect 50203 18717 50212 18751
rect 50160 18708 50212 18717
rect 52552 18844 52604 18896
rect 52552 18751 52604 18760
rect 31300 18572 31352 18624
rect 31760 18615 31812 18624
rect 31760 18581 31769 18615
rect 31769 18581 31803 18615
rect 31803 18581 31812 18615
rect 31760 18572 31812 18581
rect 32404 18572 32456 18624
rect 33140 18572 33192 18624
rect 34336 18640 34388 18692
rect 36268 18683 36320 18692
rect 36268 18649 36277 18683
rect 36277 18649 36311 18683
rect 36311 18649 36320 18683
rect 36268 18640 36320 18649
rect 49700 18640 49752 18692
rect 52552 18717 52561 18751
rect 52561 18717 52595 18751
rect 52595 18717 52604 18751
rect 52552 18708 52604 18717
rect 53196 18751 53248 18760
rect 50620 18640 50672 18692
rect 53196 18717 53205 18751
rect 53205 18717 53239 18751
rect 53239 18717 53248 18751
rect 53196 18708 53248 18717
rect 56784 18819 56836 18828
rect 56784 18785 56793 18819
rect 56793 18785 56827 18819
rect 56827 18785 56836 18819
rect 56784 18776 56836 18785
rect 57336 18819 57388 18828
rect 57336 18785 57345 18819
rect 57345 18785 57379 18819
rect 57379 18785 57388 18819
rect 57336 18776 57388 18785
rect 53472 18751 53524 18760
rect 53472 18717 53481 18751
rect 53481 18717 53515 18751
rect 53515 18717 53524 18751
rect 53472 18708 53524 18717
rect 56600 18751 56652 18760
rect 53380 18640 53432 18692
rect 56600 18717 56609 18751
rect 56609 18717 56643 18751
rect 56643 18717 56652 18751
rect 56600 18708 56652 18717
rect 57888 18751 57940 18760
rect 57888 18717 57897 18751
rect 57897 18717 57931 18751
rect 57931 18717 57940 18751
rect 57888 18708 57940 18717
rect 56692 18640 56744 18692
rect 34520 18572 34572 18624
rect 35900 18572 35952 18624
rect 52736 18615 52788 18624
rect 52736 18581 52745 18615
rect 52745 18581 52779 18615
rect 52779 18581 52788 18615
rect 52736 18572 52788 18581
rect 57796 18572 57848 18624
rect 19574 18470 19626 18522
rect 19638 18470 19690 18522
rect 19702 18470 19754 18522
rect 19766 18470 19818 18522
rect 19830 18470 19882 18522
rect 50294 18470 50346 18522
rect 50358 18470 50410 18522
rect 50422 18470 50474 18522
rect 50486 18470 50538 18522
rect 50550 18470 50602 18522
rect 2412 18368 2464 18420
rect 7564 18368 7616 18420
rect 1584 18300 1636 18352
rect 2044 18275 2096 18284
rect 2044 18241 2053 18275
rect 2053 18241 2087 18275
rect 2087 18241 2096 18275
rect 2044 18232 2096 18241
rect 2780 18275 2832 18284
rect 2780 18241 2789 18275
rect 2789 18241 2823 18275
rect 2823 18241 2832 18275
rect 3056 18275 3108 18284
rect 2780 18232 2832 18241
rect 3056 18241 3065 18275
rect 3065 18241 3099 18275
rect 3099 18241 3108 18275
rect 3056 18232 3108 18241
rect 7196 18232 7248 18284
rect 7656 18275 7708 18284
rect 7656 18241 7665 18275
rect 7665 18241 7699 18275
rect 7699 18241 7708 18275
rect 7656 18232 7708 18241
rect 7840 18275 7892 18284
rect 7840 18241 7849 18275
rect 7849 18241 7883 18275
rect 7883 18241 7892 18275
rect 7840 18232 7892 18241
rect 8024 18232 8076 18284
rect 10692 18232 10744 18284
rect 12808 18232 12860 18284
rect 15200 18368 15252 18420
rect 15292 18368 15344 18420
rect 15936 18368 15988 18420
rect 16120 18368 16172 18420
rect 18236 18368 18288 18420
rect 18420 18368 18472 18420
rect 22008 18368 22060 18420
rect 22100 18368 22152 18420
rect 23112 18368 23164 18420
rect 14648 18343 14700 18352
rect 14648 18309 14657 18343
rect 14657 18309 14691 18343
rect 14691 18309 14700 18343
rect 14648 18300 14700 18309
rect 15108 18300 15160 18352
rect 18052 18300 18104 18352
rect 14740 18275 14792 18284
rect 14740 18241 14749 18275
rect 14749 18241 14783 18275
rect 14783 18241 14792 18275
rect 14740 18232 14792 18241
rect 14832 18275 14884 18284
rect 14832 18241 14841 18275
rect 14841 18241 14875 18275
rect 14875 18241 14884 18275
rect 14832 18232 14884 18241
rect 17960 18232 18012 18284
rect 18328 18232 18380 18284
rect 20168 18300 20220 18352
rect 24124 18300 24176 18352
rect 26240 18368 26292 18420
rect 29184 18411 29236 18420
rect 29184 18377 29193 18411
rect 29193 18377 29227 18411
rect 29227 18377 29236 18411
rect 29184 18368 29236 18377
rect 30656 18368 30708 18420
rect 32864 18368 32916 18420
rect 34336 18368 34388 18420
rect 34520 18411 34572 18420
rect 34520 18377 34529 18411
rect 34529 18377 34563 18411
rect 34563 18377 34572 18411
rect 34520 18368 34572 18377
rect 35716 18368 35768 18420
rect 37372 18368 37424 18420
rect 42708 18368 42760 18420
rect 50160 18368 50212 18420
rect 53380 18411 53432 18420
rect 53380 18377 53389 18411
rect 53389 18377 53423 18411
rect 53423 18377 53432 18411
rect 53380 18368 53432 18377
rect 56692 18411 56744 18420
rect 56692 18377 56701 18411
rect 56701 18377 56735 18411
rect 56735 18377 56744 18411
rect 56692 18368 56744 18377
rect 57980 18411 58032 18420
rect 57980 18377 57989 18411
rect 57989 18377 58023 18411
rect 58023 18377 58032 18411
rect 57980 18368 58032 18377
rect 9956 18164 10008 18216
rect 16028 18164 16080 18216
rect 18880 18164 18932 18216
rect 19892 18232 19944 18284
rect 21824 18232 21876 18284
rect 24308 18232 24360 18284
rect 25044 18300 25096 18352
rect 29368 18343 29420 18352
rect 29368 18309 29377 18343
rect 29377 18309 29411 18343
rect 29411 18309 29420 18343
rect 29368 18300 29420 18309
rect 12992 18096 13044 18148
rect 13452 18096 13504 18148
rect 6000 18028 6052 18080
rect 7472 18028 7524 18080
rect 8300 18028 8352 18080
rect 12808 18028 12860 18080
rect 15200 18028 15252 18080
rect 19432 18096 19484 18148
rect 20444 18164 20496 18216
rect 24216 18164 24268 18216
rect 24952 18275 25004 18284
rect 24952 18241 24961 18275
rect 24961 18241 24995 18275
rect 24995 18241 25004 18275
rect 24952 18232 25004 18241
rect 28172 18232 28224 18284
rect 29000 18232 29052 18284
rect 26976 18164 27028 18216
rect 31024 18232 31076 18284
rect 31392 18275 31444 18284
rect 31392 18241 31401 18275
rect 31401 18241 31435 18275
rect 31435 18241 31444 18275
rect 31392 18232 31444 18241
rect 31760 18300 31812 18352
rect 33324 18232 33376 18284
rect 34336 18275 34388 18284
rect 34336 18241 34345 18275
rect 34345 18241 34379 18275
rect 34379 18241 34388 18275
rect 34336 18232 34388 18241
rect 34428 18232 34480 18284
rect 35992 18275 36044 18284
rect 35992 18241 36001 18275
rect 36001 18241 36035 18275
rect 36035 18241 36044 18275
rect 35992 18232 36044 18241
rect 36084 18275 36136 18284
rect 36084 18241 36093 18275
rect 36093 18241 36127 18275
rect 36127 18241 36136 18275
rect 36084 18232 36136 18241
rect 23480 18028 23532 18080
rect 25688 18028 25740 18080
rect 26976 18071 27028 18080
rect 26976 18037 26985 18071
rect 26985 18037 27019 18071
rect 27019 18037 27028 18071
rect 26976 18028 27028 18037
rect 30012 18028 30064 18080
rect 31484 18071 31536 18080
rect 31484 18037 31493 18071
rect 31493 18037 31527 18071
rect 31527 18037 31536 18071
rect 33600 18096 33652 18148
rect 31484 18028 31536 18037
rect 33968 18028 34020 18080
rect 35716 18164 35768 18216
rect 35808 18096 35860 18148
rect 38844 18232 38896 18284
rect 40316 18232 40368 18284
rect 40684 18275 40736 18284
rect 40684 18241 40693 18275
rect 40693 18241 40727 18275
rect 40727 18241 40736 18275
rect 40684 18232 40736 18241
rect 46020 18300 46072 18352
rect 44732 18232 44784 18284
rect 48780 18232 48832 18284
rect 48964 18275 49016 18284
rect 48964 18241 48973 18275
rect 48973 18241 49007 18275
rect 49007 18241 49016 18275
rect 48964 18232 49016 18241
rect 49148 18275 49200 18284
rect 49148 18241 49157 18275
rect 49157 18241 49191 18275
rect 49191 18241 49200 18275
rect 53472 18275 53524 18284
rect 49148 18232 49200 18241
rect 53472 18241 53481 18275
rect 53481 18241 53515 18275
rect 53515 18241 53524 18275
rect 53472 18232 53524 18241
rect 53656 18275 53708 18284
rect 53656 18241 53665 18275
rect 53665 18241 53699 18275
rect 53699 18241 53708 18275
rect 53656 18232 53708 18241
rect 56600 18275 56652 18284
rect 56600 18241 56609 18275
rect 56609 18241 56643 18275
rect 56643 18241 56652 18275
rect 56600 18232 56652 18241
rect 56784 18275 56836 18284
rect 56784 18241 56793 18275
rect 56793 18241 56827 18275
rect 56827 18241 56836 18275
rect 56784 18232 56836 18241
rect 57704 18232 57756 18284
rect 57060 18164 57112 18216
rect 57796 18164 57848 18216
rect 45100 18096 45152 18148
rect 37464 18071 37516 18080
rect 37464 18037 37473 18071
rect 37473 18037 37507 18071
rect 37507 18037 37516 18071
rect 37464 18028 37516 18037
rect 53380 18028 53432 18080
rect 4214 17926 4266 17978
rect 4278 17926 4330 17978
rect 4342 17926 4394 17978
rect 4406 17926 4458 17978
rect 4470 17926 4522 17978
rect 34934 17926 34986 17978
rect 34998 17926 35050 17978
rect 35062 17926 35114 17978
rect 35126 17926 35178 17978
rect 35190 17926 35242 17978
rect 3976 17824 4028 17876
rect 7012 17867 7064 17876
rect 7012 17833 7021 17867
rect 7021 17833 7055 17867
rect 7055 17833 7064 17867
rect 7012 17824 7064 17833
rect 7656 17867 7708 17876
rect 7656 17833 7665 17867
rect 7665 17833 7699 17867
rect 7699 17833 7708 17867
rect 7656 17824 7708 17833
rect 12624 17824 12676 17876
rect 14464 17824 14516 17876
rect 20720 17824 20772 17876
rect 22100 17824 22152 17876
rect 23204 17824 23256 17876
rect 23756 17824 23808 17876
rect 24952 17867 25004 17876
rect 24952 17833 24961 17867
rect 24961 17833 24995 17867
rect 24995 17833 25004 17867
rect 24952 17824 25004 17833
rect 30196 17824 30248 17876
rect 33232 17824 33284 17876
rect 33416 17867 33468 17876
rect 33416 17833 33425 17867
rect 33425 17833 33459 17867
rect 33459 17833 33468 17867
rect 33416 17824 33468 17833
rect 36268 17824 36320 17876
rect 45100 17867 45152 17876
rect 45100 17833 45109 17867
rect 45109 17833 45143 17867
rect 45143 17833 45152 17867
rect 45100 17824 45152 17833
rect 49700 17824 49752 17876
rect 52736 17824 52788 17876
rect 53472 17824 53524 17876
rect 56968 17867 57020 17876
rect 56968 17833 56977 17867
rect 56977 17833 57011 17867
rect 57011 17833 57020 17867
rect 56968 17824 57020 17833
rect 7196 17799 7248 17808
rect 7196 17765 7205 17799
rect 7205 17765 7239 17799
rect 7239 17765 7248 17799
rect 7196 17756 7248 17765
rect 3976 17688 4028 17740
rect 4988 17663 5040 17672
rect 4988 17629 4997 17663
rect 4997 17629 5031 17663
rect 5031 17629 5040 17663
rect 4988 17620 5040 17629
rect 6000 17663 6052 17672
rect 1584 17552 1636 17604
rect 2044 17552 2096 17604
rect 6000 17629 6009 17663
rect 6009 17629 6043 17663
rect 6043 17629 6052 17663
rect 6000 17620 6052 17629
rect 7748 17620 7800 17672
rect 8024 17620 8076 17672
rect 14372 17756 14424 17808
rect 19984 17756 20036 17808
rect 12440 17731 12492 17740
rect 12440 17697 12449 17731
rect 12449 17697 12483 17731
rect 12483 17697 12492 17731
rect 12440 17688 12492 17697
rect 13360 17688 13412 17740
rect 16672 17688 16724 17740
rect 19432 17688 19484 17740
rect 20536 17688 20588 17740
rect 12624 17663 12676 17672
rect 7288 17552 7340 17604
rect 12624 17629 12633 17663
rect 12633 17629 12667 17663
rect 12667 17629 12676 17663
rect 12624 17620 12676 17629
rect 13728 17620 13780 17672
rect 15200 17663 15252 17672
rect 15200 17629 15209 17663
rect 15209 17629 15243 17663
rect 15243 17629 15252 17663
rect 15200 17620 15252 17629
rect 18512 17620 18564 17672
rect 18604 17620 18656 17672
rect 20076 17620 20128 17672
rect 15016 17595 15068 17604
rect 15016 17561 15025 17595
rect 15025 17561 15059 17595
rect 15059 17561 15068 17595
rect 15016 17552 15068 17561
rect 15568 17595 15620 17604
rect 15568 17561 15577 17595
rect 15577 17561 15611 17595
rect 15611 17561 15620 17595
rect 15568 17552 15620 17561
rect 18236 17552 18288 17604
rect 20628 17663 20680 17672
rect 20628 17629 20642 17663
rect 20642 17629 20676 17663
rect 20676 17629 20680 17663
rect 20628 17620 20680 17629
rect 21916 17620 21968 17672
rect 24768 17756 24820 17808
rect 36084 17756 36136 17808
rect 41696 17756 41748 17808
rect 24676 17688 24728 17740
rect 26240 17688 26292 17740
rect 40224 17688 40276 17740
rect 43996 17688 44048 17740
rect 45376 17688 45428 17740
rect 53656 17731 53708 17740
rect 53656 17697 53665 17731
rect 53665 17697 53699 17731
rect 53699 17697 53708 17731
rect 53656 17688 53708 17697
rect 57060 17731 57112 17740
rect 57060 17697 57069 17731
rect 57069 17697 57103 17731
rect 57103 17697 57112 17731
rect 57060 17688 57112 17697
rect 20444 17595 20496 17604
rect 20444 17561 20453 17595
rect 20453 17561 20487 17595
rect 20487 17561 20496 17595
rect 20444 17552 20496 17561
rect 20720 17552 20772 17604
rect 23756 17620 23808 17672
rect 23480 17595 23532 17604
rect 23480 17561 23489 17595
rect 23489 17561 23523 17595
rect 23523 17561 23532 17595
rect 23480 17552 23532 17561
rect 24860 17620 24912 17672
rect 26424 17620 26476 17672
rect 30104 17620 30156 17672
rect 30656 17663 30708 17672
rect 30656 17629 30665 17663
rect 30665 17629 30699 17663
rect 30699 17629 30708 17663
rect 30656 17620 30708 17629
rect 32404 17620 32456 17672
rect 24584 17595 24636 17604
rect 24584 17561 24593 17595
rect 24593 17561 24627 17595
rect 24627 17561 24636 17595
rect 24584 17552 24636 17561
rect 24952 17552 25004 17604
rect 25964 17552 26016 17604
rect 26976 17552 27028 17604
rect 28632 17552 28684 17604
rect 32588 17552 32640 17604
rect 33416 17620 33468 17672
rect 40500 17620 40552 17672
rect 44180 17663 44232 17672
rect 44180 17629 44189 17663
rect 44189 17629 44223 17663
rect 44223 17629 44232 17663
rect 44180 17620 44232 17629
rect 44732 17620 44784 17672
rect 35900 17552 35952 17604
rect 36544 17552 36596 17604
rect 44088 17552 44140 17604
rect 48964 17620 49016 17672
rect 48320 17595 48372 17604
rect 48320 17561 48329 17595
rect 48329 17561 48363 17595
rect 48363 17561 48372 17595
rect 48320 17552 48372 17561
rect 48504 17595 48556 17604
rect 48504 17561 48513 17595
rect 48513 17561 48547 17595
rect 48547 17561 48556 17595
rect 48504 17552 48556 17561
rect 49148 17552 49200 17604
rect 53380 17620 53432 17672
rect 56692 17620 56744 17672
rect 56968 17620 57020 17672
rect 58072 17663 58124 17672
rect 58072 17629 58081 17663
rect 58081 17629 58115 17663
rect 58115 17629 58124 17663
rect 58072 17620 58124 17629
rect 56324 17552 56376 17604
rect 8208 17484 8260 17536
rect 8944 17527 8996 17536
rect 8944 17493 8953 17527
rect 8953 17493 8987 17527
rect 8987 17493 8996 17527
rect 8944 17484 8996 17493
rect 14004 17484 14056 17536
rect 16948 17484 17000 17536
rect 18328 17527 18380 17536
rect 18328 17493 18337 17527
rect 18337 17493 18371 17527
rect 18371 17493 18380 17527
rect 18328 17484 18380 17493
rect 20812 17527 20864 17536
rect 20812 17493 20821 17527
rect 20821 17493 20855 17527
rect 20855 17493 20864 17527
rect 20812 17484 20864 17493
rect 23204 17484 23256 17536
rect 23848 17527 23900 17536
rect 23848 17493 23857 17527
rect 23857 17493 23891 17527
rect 23891 17493 23900 17527
rect 23848 17484 23900 17493
rect 26332 17527 26384 17536
rect 26332 17493 26341 17527
rect 26341 17493 26375 17527
rect 26375 17493 26384 17527
rect 26332 17484 26384 17493
rect 28724 17484 28776 17536
rect 30840 17527 30892 17536
rect 30840 17493 30849 17527
rect 30849 17493 30883 17527
rect 30883 17493 30892 17527
rect 30840 17484 30892 17493
rect 33784 17484 33836 17536
rect 34428 17484 34480 17536
rect 40224 17527 40276 17536
rect 40224 17493 40233 17527
rect 40233 17493 40267 17527
rect 40267 17493 40276 17527
rect 40224 17484 40276 17493
rect 48780 17484 48832 17536
rect 52552 17484 52604 17536
rect 53564 17484 53616 17536
rect 19574 17382 19626 17434
rect 19638 17382 19690 17434
rect 19702 17382 19754 17434
rect 19766 17382 19818 17434
rect 19830 17382 19882 17434
rect 50294 17382 50346 17434
rect 50358 17382 50410 17434
rect 50422 17382 50474 17434
rect 50486 17382 50538 17434
rect 50550 17382 50602 17434
rect 3056 17280 3108 17332
rect 3516 17280 3568 17332
rect 8944 17280 8996 17332
rect 9128 17280 9180 17332
rect 16580 17280 16632 17332
rect 20076 17323 20128 17332
rect 20076 17289 20085 17323
rect 20085 17289 20119 17323
rect 20119 17289 20128 17323
rect 20076 17280 20128 17289
rect 20352 17280 20404 17332
rect 24584 17280 24636 17332
rect 28356 17280 28408 17332
rect 4988 17212 5040 17264
rect 7472 17255 7524 17264
rect 7472 17221 7481 17255
rect 7481 17221 7515 17255
rect 7515 17221 7524 17255
rect 7472 17212 7524 17221
rect 8024 17212 8076 17264
rect 8208 17212 8260 17264
rect 10416 17212 10468 17264
rect 2872 17119 2924 17128
rect 2872 17085 2881 17119
rect 2881 17085 2915 17119
rect 2915 17085 2924 17119
rect 2872 17076 2924 17085
rect 7288 17119 7340 17128
rect 7288 17085 7297 17119
rect 7297 17085 7331 17119
rect 7331 17085 7340 17119
rect 9956 17187 10008 17196
rect 9956 17153 9965 17187
rect 9965 17153 9999 17187
rect 9999 17153 10008 17187
rect 9956 17144 10008 17153
rect 10140 17144 10192 17196
rect 12900 17212 12952 17264
rect 13728 17212 13780 17264
rect 14096 17187 14148 17196
rect 14096 17153 14105 17187
rect 14105 17153 14139 17187
rect 14139 17153 14148 17187
rect 14096 17144 14148 17153
rect 14372 17187 14424 17196
rect 14372 17153 14381 17187
rect 14381 17153 14415 17187
rect 14415 17153 14424 17187
rect 14372 17144 14424 17153
rect 14556 17144 14608 17196
rect 14740 17144 14792 17196
rect 15200 17144 15252 17196
rect 7288 17076 7340 17085
rect 9036 17076 9088 17128
rect 12440 17076 12492 17128
rect 3424 17008 3476 17060
rect 8208 17008 8260 17060
rect 1860 16940 1912 16992
rect 7840 16940 7892 16992
rect 8484 16983 8536 16992
rect 8484 16949 8493 16983
rect 8493 16949 8527 16983
rect 8527 16949 8536 16983
rect 8484 16940 8536 16949
rect 15292 17008 15344 17060
rect 17960 17008 18012 17060
rect 19524 17187 19576 17196
rect 19524 17153 19533 17187
rect 19533 17153 19567 17187
rect 19567 17153 19576 17187
rect 19524 17144 19576 17153
rect 19708 17187 19760 17196
rect 19708 17153 19717 17187
rect 19717 17153 19751 17187
rect 19751 17153 19760 17187
rect 19708 17144 19760 17153
rect 20168 17144 20220 17196
rect 20352 17144 20404 17196
rect 20536 17187 20588 17196
rect 20536 17153 20545 17187
rect 20545 17153 20579 17187
rect 20579 17153 20588 17187
rect 20536 17144 20588 17153
rect 22744 17212 22796 17264
rect 24676 17255 24728 17264
rect 24676 17221 24685 17255
rect 24685 17221 24719 17255
rect 24719 17221 24728 17255
rect 24676 17212 24728 17221
rect 24860 17212 24912 17264
rect 24308 17144 24360 17196
rect 28172 17144 28224 17196
rect 28448 17144 28500 17196
rect 28724 17280 28776 17332
rect 29920 17280 29972 17332
rect 37464 17280 37516 17332
rect 31024 17187 31076 17196
rect 19432 17076 19484 17128
rect 26332 17076 26384 17128
rect 31024 17153 31033 17187
rect 31033 17153 31067 17187
rect 31067 17153 31076 17187
rect 31024 17144 31076 17153
rect 36452 17212 36504 17264
rect 36544 17255 36596 17264
rect 36544 17221 36553 17255
rect 36553 17221 36587 17255
rect 36587 17221 36596 17255
rect 36544 17212 36596 17221
rect 31300 17076 31352 17128
rect 32404 17144 32456 17196
rect 32956 17144 33008 17196
rect 33508 17187 33560 17196
rect 33508 17153 33517 17187
rect 33517 17153 33551 17187
rect 33551 17153 33560 17187
rect 33508 17144 33560 17153
rect 33692 17144 33744 17196
rect 34428 17144 34480 17196
rect 37372 17144 37424 17196
rect 44272 17280 44324 17332
rect 48320 17280 48372 17332
rect 53104 17280 53156 17332
rect 58072 17323 58124 17332
rect 58072 17289 58081 17323
rect 58081 17289 58115 17323
rect 58115 17289 58124 17323
rect 58072 17280 58124 17289
rect 43904 17212 43956 17264
rect 44088 17212 44140 17264
rect 56324 17212 56376 17264
rect 56784 17212 56836 17264
rect 40500 17144 40552 17196
rect 43996 17144 44048 17196
rect 45376 17187 45428 17196
rect 45376 17153 45385 17187
rect 45385 17153 45419 17187
rect 45419 17153 45428 17187
rect 48136 17187 48188 17196
rect 45376 17144 45428 17153
rect 48136 17153 48145 17187
rect 48145 17153 48179 17187
rect 48179 17153 48188 17187
rect 48136 17144 48188 17153
rect 21640 17008 21692 17060
rect 23296 17008 23348 17060
rect 27620 17008 27672 17060
rect 30840 17008 30892 17060
rect 35348 17008 35400 17060
rect 10140 16940 10192 16992
rect 15016 16940 15068 16992
rect 15476 16940 15528 16992
rect 16304 16940 16356 16992
rect 20076 16940 20128 16992
rect 20168 16940 20220 16992
rect 25228 16940 25280 16992
rect 26792 16940 26844 16992
rect 29184 16940 29236 16992
rect 29828 16940 29880 16992
rect 30012 16983 30064 16992
rect 30012 16949 30021 16983
rect 30021 16949 30055 16983
rect 30055 16949 30064 16983
rect 30012 16940 30064 16949
rect 31392 16940 31444 16992
rect 32680 16983 32732 16992
rect 32680 16949 32689 16983
rect 32689 16949 32723 16983
rect 32723 16949 32732 16983
rect 32680 16940 32732 16949
rect 33784 16983 33836 16992
rect 33784 16949 33793 16983
rect 33793 16949 33827 16983
rect 33827 16949 33836 16983
rect 33784 16940 33836 16949
rect 36360 16940 36412 16992
rect 48504 17119 48556 17128
rect 48504 17085 48513 17119
rect 48513 17085 48547 17119
rect 48547 17085 48556 17119
rect 48504 17076 48556 17085
rect 48136 17008 48188 17060
rect 50804 17187 50856 17196
rect 50804 17153 50813 17187
rect 50813 17153 50847 17187
rect 50847 17153 50856 17187
rect 50804 17144 50856 17153
rect 52552 17144 52604 17196
rect 53196 17144 53248 17196
rect 53656 17187 53708 17196
rect 53656 17153 53665 17187
rect 53665 17153 53699 17187
rect 53699 17153 53708 17187
rect 53656 17144 53708 17153
rect 53748 17144 53800 17196
rect 57152 17144 57204 17196
rect 50252 17119 50304 17128
rect 50252 17085 50261 17119
rect 50261 17085 50295 17119
rect 50295 17085 50304 17119
rect 50252 17076 50304 17085
rect 53472 17119 53524 17128
rect 53472 17085 53481 17119
rect 53481 17085 53515 17119
rect 53515 17085 53524 17119
rect 53472 17076 53524 17085
rect 56140 17076 56192 17128
rect 52736 17051 52788 17060
rect 40040 16983 40092 16992
rect 40040 16949 40049 16983
rect 40049 16949 40083 16983
rect 40083 16949 40092 16983
rect 40040 16940 40092 16949
rect 44180 16940 44232 16992
rect 45284 16983 45336 16992
rect 45284 16949 45293 16983
rect 45293 16949 45327 16983
rect 45327 16949 45336 16983
rect 45284 16940 45336 16949
rect 51172 16940 51224 16992
rect 52736 17017 52745 17051
rect 52745 17017 52779 17051
rect 52779 17017 52788 17051
rect 52736 17008 52788 17017
rect 56324 17008 56376 17060
rect 51632 16983 51684 16992
rect 51632 16949 51641 16983
rect 51641 16949 51675 16983
rect 51675 16949 51684 16983
rect 51632 16940 51684 16949
rect 51816 16940 51868 16992
rect 56140 16940 56192 16992
rect 4214 16838 4266 16890
rect 4278 16838 4330 16890
rect 4342 16838 4394 16890
rect 4406 16838 4458 16890
rect 4470 16838 4522 16890
rect 34934 16838 34986 16890
rect 34998 16838 35050 16890
rect 35062 16838 35114 16890
rect 35126 16838 35178 16890
rect 35190 16838 35242 16890
rect 3332 16736 3384 16788
rect 7012 16736 7064 16788
rect 7840 16779 7892 16788
rect 7840 16745 7849 16779
rect 7849 16745 7883 16779
rect 7883 16745 7892 16779
rect 7840 16736 7892 16745
rect 9036 16736 9088 16788
rect 10048 16736 10100 16788
rect 12900 16779 12952 16788
rect 12900 16745 12909 16779
rect 12909 16745 12943 16779
rect 12943 16745 12952 16779
rect 12900 16736 12952 16745
rect 14464 16736 14516 16788
rect 33048 16736 33100 16788
rect 2872 16711 2924 16720
rect 2872 16677 2881 16711
rect 2881 16677 2915 16711
rect 2915 16677 2924 16711
rect 2872 16668 2924 16677
rect 9128 16668 9180 16720
rect 9956 16668 10008 16720
rect 11888 16668 11940 16720
rect 13544 16668 13596 16720
rect 14096 16668 14148 16720
rect 3424 16600 3476 16652
rect 4160 16575 4212 16584
rect 4160 16541 4169 16575
rect 4169 16541 4203 16575
rect 4203 16541 4212 16575
rect 4160 16532 4212 16541
rect 4620 16575 4672 16584
rect 4620 16541 4629 16575
rect 4629 16541 4663 16575
rect 4663 16541 4672 16575
rect 4620 16532 4672 16541
rect 7472 16532 7524 16584
rect 1860 16507 1912 16516
rect 1860 16473 1869 16507
rect 1869 16473 1903 16507
rect 1903 16473 1912 16507
rect 1860 16464 1912 16473
rect 8484 16532 8536 16584
rect 9036 16532 9088 16584
rect 8208 16464 8260 16516
rect 9220 16507 9272 16516
rect 9220 16473 9229 16507
rect 9229 16473 9263 16507
rect 9263 16473 9272 16507
rect 9220 16464 9272 16473
rect 9312 16464 9364 16516
rect 9680 16532 9732 16584
rect 10140 16464 10192 16516
rect 10416 16507 10468 16516
rect 10416 16473 10425 16507
rect 10425 16473 10459 16507
rect 10459 16473 10468 16507
rect 10416 16464 10468 16473
rect 12440 16507 12492 16516
rect 12440 16473 12449 16507
rect 12449 16473 12483 16507
rect 12483 16473 12492 16507
rect 14832 16600 14884 16652
rect 15292 16668 15344 16720
rect 14556 16575 14608 16584
rect 14556 16541 14565 16575
rect 14565 16541 14599 16575
rect 14599 16541 14608 16575
rect 14556 16532 14608 16541
rect 15476 16575 15528 16584
rect 15476 16541 15485 16575
rect 15485 16541 15519 16575
rect 15519 16541 15528 16575
rect 15476 16532 15528 16541
rect 16120 16600 16172 16652
rect 19524 16668 19576 16720
rect 19708 16643 19760 16652
rect 16672 16532 16724 16584
rect 19708 16609 19717 16643
rect 19717 16609 19751 16643
rect 19751 16609 19760 16643
rect 19708 16600 19760 16609
rect 19800 16532 19852 16584
rect 20168 16575 20220 16584
rect 12440 16464 12492 16473
rect 14464 16507 14516 16516
rect 14464 16473 14473 16507
rect 14473 16473 14507 16507
rect 14507 16473 14516 16507
rect 14464 16464 14516 16473
rect 20168 16541 20177 16575
rect 20177 16541 20211 16575
rect 20211 16541 20220 16575
rect 20168 16532 20220 16541
rect 20352 16532 20404 16584
rect 21272 16575 21324 16584
rect 21272 16541 21281 16575
rect 21281 16541 21315 16575
rect 21315 16541 21324 16575
rect 21272 16532 21324 16541
rect 23296 16532 23348 16584
rect 23848 16575 23900 16584
rect 23848 16541 23857 16575
rect 23857 16541 23891 16575
rect 23891 16541 23900 16575
rect 23848 16532 23900 16541
rect 2780 16439 2832 16448
rect 2780 16405 2789 16439
rect 2789 16405 2823 16439
rect 2823 16405 2832 16439
rect 10600 16439 10652 16448
rect 2780 16396 2832 16405
rect 10600 16405 10609 16439
rect 10609 16405 10643 16439
rect 10643 16405 10652 16439
rect 10600 16396 10652 16405
rect 20444 16464 20496 16516
rect 20720 16464 20772 16516
rect 27712 16600 27764 16652
rect 28356 16643 28408 16652
rect 28356 16609 28365 16643
rect 28365 16609 28399 16643
rect 28399 16609 28408 16643
rect 30840 16643 30892 16652
rect 28356 16600 28408 16609
rect 30840 16609 30849 16643
rect 30849 16609 30883 16643
rect 30883 16609 30892 16643
rect 30840 16600 30892 16609
rect 31392 16643 31444 16652
rect 31392 16609 31401 16643
rect 31401 16609 31435 16643
rect 31435 16609 31444 16643
rect 31392 16600 31444 16609
rect 32496 16600 32548 16652
rect 33784 16600 33836 16652
rect 35256 16643 35308 16652
rect 35256 16609 35265 16643
rect 35265 16609 35299 16643
rect 35299 16609 35308 16643
rect 35256 16600 35308 16609
rect 45928 16736 45980 16788
rect 48136 16736 48188 16788
rect 50160 16779 50212 16788
rect 50160 16745 50169 16779
rect 50169 16745 50203 16779
rect 50203 16745 50212 16779
rect 50160 16736 50212 16745
rect 50804 16736 50856 16788
rect 53472 16736 53524 16788
rect 53656 16779 53708 16788
rect 53656 16745 53665 16779
rect 53665 16745 53699 16779
rect 53699 16745 53708 16779
rect 53656 16736 53708 16745
rect 53748 16736 53800 16788
rect 43996 16711 44048 16720
rect 38752 16643 38804 16652
rect 38752 16609 38761 16643
rect 38761 16609 38795 16643
rect 38795 16609 38804 16643
rect 38752 16600 38804 16609
rect 43996 16677 44005 16711
rect 44005 16677 44039 16711
rect 44039 16677 44048 16711
rect 43996 16668 44048 16677
rect 24124 16532 24176 16584
rect 24492 16575 24544 16584
rect 24492 16541 24501 16575
rect 24501 16541 24535 16575
rect 24535 16541 24544 16575
rect 24492 16532 24544 16541
rect 26424 16575 26476 16584
rect 26424 16541 26433 16575
rect 26433 16541 26467 16575
rect 26467 16541 26476 16575
rect 26424 16532 26476 16541
rect 26516 16575 26568 16584
rect 26516 16541 26526 16575
rect 26526 16541 26560 16575
rect 26560 16541 26568 16575
rect 26792 16575 26844 16584
rect 26516 16532 26568 16541
rect 26792 16541 26801 16575
rect 26801 16541 26835 16575
rect 26835 16541 26844 16575
rect 26792 16532 26844 16541
rect 28080 16575 28132 16584
rect 15844 16396 15896 16448
rect 16304 16439 16356 16448
rect 16304 16405 16313 16439
rect 16313 16405 16347 16439
rect 16347 16405 16356 16439
rect 16304 16396 16356 16405
rect 20076 16396 20128 16448
rect 23388 16396 23440 16448
rect 25136 16396 25188 16448
rect 28080 16541 28089 16575
rect 28089 16541 28123 16575
rect 28123 16541 28132 16575
rect 28080 16532 28132 16541
rect 28632 16532 28684 16584
rect 32956 16575 33008 16584
rect 32956 16541 32965 16575
rect 32965 16541 32999 16575
rect 32999 16541 33008 16575
rect 32956 16532 33008 16541
rect 33968 16532 34020 16584
rect 36084 16532 36136 16584
rect 37188 16532 37240 16584
rect 38660 16575 38712 16584
rect 38660 16541 38669 16575
rect 38669 16541 38703 16575
rect 38703 16541 38712 16575
rect 38660 16532 38712 16541
rect 43260 16532 43312 16584
rect 28448 16464 28500 16516
rect 26884 16396 26936 16448
rect 29828 16396 29880 16448
rect 42524 16464 42576 16516
rect 43904 16532 43956 16584
rect 45928 16575 45980 16584
rect 45928 16541 45937 16575
rect 45937 16541 45971 16575
rect 45971 16541 45980 16575
rect 50252 16668 50304 16720
rect 53104 16668 53156 16720
rect 51172 16600 51224 16652
rect 45928 16532 45980 16541
rect 51632 16600 51684 16652
rect 51816 16575 51868 16584
rect 51816 16541 51825 16575
rect 51825 16541 51859 16575
rect 51859 16541 51868 16575
rect 51816 16532 51868 16541
rect 52552 16600 52604 16652
rect 57152 16643 57204 16652
rect 53196 16575 53248 16584
rect 53196 16541 53205 16575
rect 53205 16541 53239 16575
rect 53239 16541 53248 16575
rect 57152 16609 57161 16643
rect 57161 16609 57195 16643
rect 57195 16609 57204 16643
rect 57152 16600 57204 16609
rect 53196 16532 53248 16541
rect 32496 16396 32548 16448
rect 32680 16396 32732 16448
rect 34520 16396 34572 16448
rect 39212 16396 39264 16448
rect 41972 16396 42024 16448
rect 44456 16464 44508 16516
rect 43812 16439 43864 16448
rect 43812 16405 43821 16439
rect 43821 16405 43855 16439
rect 43855 16405 43864 16439
rect 43812 16396 43864 16405
rect 53104 16396 53156 16448
rect 56232 16575 56284 16584
rect 56232 16541 56241 16575
rect 56241 16541 56275 16575
rect 56275 16541 56284 16575
rect 56232 16532 56284 16541
rect 56324 16532 56376 16584
rect 58164 16575 58216 16584
rect 58164 16541 58173 16575
rect 58173 16541 58207 16575
rect 58207 16541 58216 16575
rect 58164 16532 58216 16541
rect 57704 16396 57756 16448
rect 19574 16294 19626 16346
rect 19638 16294 19690 16346
rect 19702 16294 19754 16346
rect 19766 16294 19818 16346
rect 19830 16294 19882 16346
rect 50294 16294 50346 16346
rect 50358 16294 50410 16346
rect 50422 16294 50474 16346
rect 50486 16294 50538 16346
rect 50550 16294 50602 16346
rect 1768 16235 1820 16244
rect 1768 16201 1777 16235
rect 1777 16201 1811 16235
rect 1811 16201 1820 16235
rect 1768 16192 1820 16201
rect 4160 16192 4212 16244
rect 8208 16235 8260 16244
rect 8208 16201 8217 16235
rect 8217 16201 8251 16235
rect 8251 16201 8260 16235
rect 8208 16192 8260 16201
rect 8668 16192 8720 16244
rect 9312 16192 9364 16244
rect 9588 16192 9640 16244
rect 13544 16235 13596 16244
rect 2688 16124 2740 16176
rect 2780 16056 2832 16108
rect 3516 16099 3568 16108
rect 3516 16065 3525 16099
rect 3525 16065 3559 16099
rect 3559 16065 3568 16099
rect 3516 16056 3568 16065
rect 7196 16099 7248 16108
rect 7196 16065 7205 16099
rect 7205 16065 7239 16099
rect 7239 16065 7248 16099
rect 7196 16056 7248 16065
rect 7564 16099 7616 16108
rect 7564 16065 7573 16099
rect 7573 16065 7607 16099
rect 7607 16065 7616 16099
rect 7564 16056 7616 16065
rect 8116 16056 8168 16108
rect 9036 16099 9088 16108
rect 9036 16065 9045 16099
rect 9045 16065 9079 16099
rect 9079 16065 9088 16099
rect 9036 16056 9088 16065
rect 9220 16056 9272 16108
rect 9956 16099 10008 16108
rect 9956 16065 9965 16099
rect 9965 16065 9999 16099
rect 9999 16065 10008 16099
rect 9956 16056 10008 16065
rect 12440 16124 12492 16176
rect 10968 16056 11020 16108
rect 10048 15988 10100 16040
rect 13544 16201 13553 16235
rect 13553 16201 13587 16235
rect 13587 16201 13596 16235
rect 13544 16192 13596 16201
rect 13636 16124 13688 16176
rect 14188 16056 14240 16108
rect 2872 15920 2924 15972
rect 3792 15920 3844 15972
rect 6920 15920 6972 15972
rect 10508 15920 10560 15972
rect 13360 15988 13412 16040
rect 17316 16124 17368 16176
rect 17960 16124 18012 16176
rect 21272 16192 21324 16244
rect 26240 16192 26292 16244
rect 26424 16192 26476 16244
rect 15844 16056 15896 16108
rect 16120 16099 16172 16108
rect 16120 16065 16129 16099
rect 16129 16065 16163 16099
rect 16163 16065 16172 16099
rect 16120 16056 16172 16065
rect 19340 16056 19392 16108
rect 19616 16099 19668 16108
rect 19616 16065 19625 16099
rect 19625 16065 19659 16099
rect 19659 16065 19668 16099
rect 19616 16056 19668 16065
rect 20444 16124 20496 16176
rect 20996 16124 21048 16176
rect 22376 16124 22428 16176
rect 14924 15988 14976 16040
rect 11336 15920 11388 15972
rect 19432 15920 19484 15972
rect 15292 15852 15344 15904
rect 16396 15852 16448 15904
rect 16856 15852 16908 15904
rect 18880 15852 18932 15904
rect 19064 15895 19116 15904
rect 19064 15861 19073 15895
rect 19073 15861 19107 15895
rect 19107 15861 19116 15895
rect 20168 16056 20220 16108
rect 20628 16056 20680 16108
rect 22836 16056 22888 16108
rect 23296 16099 23348 16108
rect 21732 15988 21784 16040
rect 23296 16065 23305 16099
rect 23305 16065 23339 16099
rect 23339 16065 23348 16099
rect 23296 16056 23348 16065
rect 25044 16124 25096 16176
rect 26516 16124 26568 16176
rect 27252 16124 27304 16176
rect 23204 15988 23256 16040
rect 24124 16056 24176 16108
rect 24952 16056 25004 16108
rect 27620 16192 27672 16244
rect 27712 16192 27764 16244
rect 32496 16235 32548 16244
rect 28080 16124 28132 16176
rect 28448 16167 28500 16176
rect 28448 16133 28457 16167
rect 28457 16133 28491 16167
rect 28491 16133 28500 16167
rect 28448 16124 28500 16133
rect 29184 16167 29236 16176
rect 29184 16133 29193 16167
rect 29193 16133 29227 16167
rect 29227 16133 29236 16167
rect 29184 16124 29236 16133
rect 25044 15988 25096 16040
rect 27436 16099 27488 16108
rect 27436 16065 27445 16099
rect 27445 16065 27479 16099
rect 27479 16065 27488 16099
rect 27436 16056 27488 16065
rect 28172 16056 28224 16108
rect 29092 16056 29144 16108
rect 29644 16056 29696 16108
rect 20352 15920 20404 15972
rect 19064 15852 19116 15861
rect 20628 15852 20680 15904
rect 22376 15920 22428 15972
rect 32496 16201 32505 16235
rect 32505 16201 32539 16235
rect 32539 16201 32548 16235
rect 32496 16192 32548 16201
rect 34428 16192 34480 16244
rect 43996 16192 44048 16244
rect 53196 16192 53248 16244
rect 58164 16235 58216 16244
rect 58164 16201 58173 16235
rect 58173 16201 58207 16235
rect 58207 16201 58216 16235
rect 58164 16192 58216 16201
rect 35256 16124 35308 16176
rect 38568 16124 38620 16176
rect 43812 16124 43864 16176
rect 34520 16056 34572 16108
rect 35808 16056 35860 16108
rect 36360 16099 36412 16108
rect 36360 16065 36369 16099
rect 36369 16065 36403 16099
rect 36403 16065 36412 16099
rect 36360 16056 36412 16065
rect 36544 16056 36596 16108
rect 38660 16099 38712 16108
rect 38660 16065 38669 16099
rect 38669 16065 38703 16099
rect 38703 16065 38712 16099
rect 38660 16056 38712 16065
rect 38936 16056 38988 16108
rect 42800 16099 42852 16108
rect 42800 16065 42809 16099
rect 42809 16065 42843 16099
rect 42843 16065 42852 16099
rect 42800 16056 42852 16065
rect 43260 16056 43312 16108
rect 43904 16056 43956 16108
rect 56140 16124 56192 16176
rect 52920 16056 52972 16108
rect 56324 16056 56376 16108
rect 57152 16056 57204 16108
rect 34060 15988 34112 16040
rect 34336 15988 34388 16040
rect 24492 15852 24544 15904
rect 24768 15895 24820 15904
rect 24768 15861 24777 15895
rect 24777 15861 24811 15895
rect 24811 15861 24820 15895
rect 24768 15852 24820 15861
rect 26240 15852 26292 15904
rect 29828 15852 29880 15904
rect 44088 15988 44140 16040
rect 44456 16031 44508 16040
rect 44456 15997 44465 16031
rect 44465 15997 44499 16031
rect 44499 15997 44508 16031
rect 44456 15988 44508 15997
rect 52828 15988 52880 16040
rect 48688 15920 48740 15972
rect 39212 15852 39264 15904
rect 44180 15852 44232 15904
rect 47308 15852 47360 15904
rect 53012 15852 53064 15904
rect 56324 15895 56376 15904
rect 56324 15861 56333 15895
rect 56333 15861 56367 15895
rect 56367 15861 56376 15895
rect 56324 15852 56376 15861
rect 56784 15895 56836 15904
rect 56784 15861 56793 15895
rect 56793 15861 56827 15895
rect 56827 15861 56836 15895
rect 56784 15852 56836 15861
rect 4214 15750 4266 15802
rect 4278 15750 4330 15802
rect 4342 15750 4394 15802
rect 4406 15750 4458 15802
rect 4470 15750 4522 15802
rect 34934 15750 34986 15802
rect 34998 15750 35050 15802
rect 35062 15750 35114 15802
rect 35126 15750 35178 15802
rect 35190 15750 35242 15802
rect 2688 15648 2740 15700
rect 9036 15648 9088 15700
rect 9680 15580 9732 15632
rect 9220 15512 9272 15564
rect 3792 15487 3844 15496
rect 3792 15453 3801 15487
rect 3801 15453 3835 15487
rect 3835 15453 3844 15487
rect 3792 15444 3844 15453
rect 4620 15444 4672 15496
rect 6920 15487 6972 15496
rect 6920 15453 6929 15487
rect 6929 15453 6963 15487
rect 6963 15453 6972 15487
rect 6920 15444 6972 15453
rect 7748 15487 7800 15496
rect 7748 15453 7757 15487
rect 7757 15453 7791 15487
rect 7791 15453 7800 15487
rect 7748 15444 7800 15453
rect 9680 15444 9732 15496
rect 13728 15648 13780 15700
rect 14556 15648 14608 15700
rect 14648 15648 14700 15700
rect 10600 15580 10652 15632
rect 13360 15580 13412 15632
rect 13544 15623 13596 15632
rect 13544 15589 13553 15623
rect 13553 15589 13587 15623
rect 13587 15589 13596 15623
rect 13544 15580 13596 15589
rect 11336 15555 11388 15564
rect 10048 15444 10100 15496
rect 11336 15521 11345 15555
rect 11345 15521 11379 15555
rect 11379 15521 11388 15555
rect 11336 15512 11388 15521
rect 10784 15487 10836 15496
rect 10784 15453 10793 15487
rect 10793 15453 10827 15487
rect 10827 15453 10836 15487
rect 14648 15512 14700 15564
rect 19616 15648 19668 15700
rect 22836 15691 22888 15700
rect 22836 15657 22845 15691
rect 22845 15657 22879 15691
rect 22879 15657 22888 15691
rect 22836 15648 22888 15657
rect 26884 15648 26936 15700
rect 27436 15648 27488 15700
rect 29092 15648 29144 15700
rect 29644 15648 29696 15700
rect 31024 15691 31076 15700
rect 31024 15657 31033 15691
rect 31033 15657 31067 15691
rect 31067 15657 31076 15691
rect 31024 15648 31076 15657
rect 32036 15648 32088 15700
rect 32404 15648 32456 15700
rect 39856 15691 39908 15700
rect 39856 15657 39865 15691
rect 39865 15657 39899 15691
rect 39899 15657 39908 15691
rect 39856 15648 39908 15657
rect 43812 15648 43864 15700
rect 19432 15580 19484 15632
rect 20076 15580 20128 15632
rect 20444 15580 20496 15632
rect 20904 15580 20956 15632
rect 20352 15512 20404 15564
rect 14188 15487 14240 15496
rect 10784 15444 10836 15453
rect 14188 15453 14197 15487
rect 14197 15453 14231 15487
rect 14231 15453 14240 15487
rect 14188 15444 14240 15453
rect 10416 15376 10468 15428
rect 13544 15376 13596 15428
rect 14464 15444 14516 15496
rect 15108 15487 15160 15496
rect 15108 15453 15117 15487
rect 15117 15453 15151 15487
rect 15151 15453 15160 15487
rect 15108 15444 15160 15453
rect 15476 15444 15528 15496
rect 15752 15444 15804 15496
rect 16396 15487 16448 15496
rect 16396 15453 16405 15487
rect 16405 15453 16439 15487
rect 16439 15453 16448 15487
rect 16396 15444 16448 15453
rect 16580 15487 16632 15496
rect 16580 15453 16587 15487
rect 16587 15453 16632 15487
rect 16580 15444 16632 15453
rect 16948 15444 17000 15496
rect 19340 15444 19392 15496
rect 19432 15487 19484 15496
rect 19432 15453 19441 15487
rect 19441 15453 19475 15487
rect 19475 15453 19484 15487
rect 19432 15444 19484 15453
rect 20260 15444 20312 15496
rect 16764 15419 16816 15428
rect 16764 15385 16773 15419
rect 16773 15385 16807 15419
rect 16807 15385 16816 15419
rect 16764 15376 16816 15385
rect 21732 15444 21784 15496
rect 23756 15580 23808 15632
rect 24308 15580 24360 15632
rect 24768 15580 24820 15632
rect 30840 15580 30892 15632
rect 36360 15580 36412 15632
rect 37372 15580 37424 15632
rect 23112 15419 23164 15428
rect 23112 15385 23121 15419
rect 23121 15385 23155 15419
rect 23155 15385 23164 15419
rect 23112 15376 23164 15385
rect 23480 15512 23532 15564
rect 24676 15512 24728 15564
rect 23388 15487 23440 15496
rect 23388 15453 23397 15487
rect 23397 15453 23431 15487
rect 23431 15453 23440 15487
rect 23388 15444 23440 15453
rect 24400 15444 24452 15496
rect 26240 15512 26292 15564
rect 28540 15512 28592 15564
rect 32680 15512 32732 15564
rect 52552 15648 52604 15700
rect 53104 15691 53156 15700
rect 25228 15444 25280 15496
rect 3792 15308 3844 15360
rect 8944 15351 8996 15360
rect 8944 15317 8953 15351
rect 8953 15317 8987 15351
rect 8987 15317 8996 15351
rect 8944 15308 8996 15317
rect 10692 15351 10744 15360
rect 10692 15317 10701 15351
rect 10701 15317 10735 15351
rect 10735 15317 10744 15351
rect 10692 15308 10744 15317
rect 14280 15308 14332 15360
rect 15844 15308 15896 15360
rect 17592 15308 17644 15360
rect 20260 15308 20312 15360
rect 21916 15308 21968 15360
rect 22284 15308 22336 15360
rect 24860 15376 24912 15428
rect 26884 15376 26936 15428
rect 25872 15351 25924 15360
rect 25872 15317 25881 15351
rect 25881 15317 25915 15351
rect 25915 15317 25924 15351
rect 25872 15308 25924 15317
rect 31392 15308 31444 15360
rect 32312 15444 32364 15496
rect 33140 15444 33192 15496
rect 40592 15487 40644 15496
rect 40592 15453 40601 15487
rect 40601 15453 40635 15487
rect 40635 15453 40644 15487
rect 40592 15444 40644 15453
rect 41972 15487 42024 15496
rect 41972 15453 41981 15487
rect 41981 15453 42015 15487
rect 42015 15453 42024 15487
rect 41972 15444 42024 15453
rect 42524 15487 42576 15496
rect 42524 15453 42533 15487
rect 42533 15453 42567 15487
rect 42567 15453 42576 15487
rect 42524 15444 42576 15453
rect 42800 15487 42852 15496
rect 42800 15453 42809 15487
rect 42809 15453 42843 15487
rect 42843 15453 42852 15487
rect 42800 15444 42852 15453
rect 43904 15419 43956 15428
rect 43904 15385 43913 15419
rect 43913 15385 43947 15419
rect 43947 15385 43956 15419
rect 43904 15376 43956 15385
rect 32128 15351 32180 15360
rect 32128 15317 32137 15351
rect 32137 15317 32171 15351
rect 32171 15317 32180 15351
rect 32128 15308 32180 15317
rect 32220 15308 32272 15360
rect 32404 15351 32456 15360
rect 32404 15317 32413 15351
rect 32413 15317 32447 15351
rect 32447 15317 32456 15351
rect 32404 15308 32456 15317
rect 33324 15308 33376 15360
rect 33508 15351 33560 15360
rect 33508 15317 33517 15351
rect 33517 15317 33551 15351
rect 33551 15317 33560 15351
rect 33508 15308 33560 15317
rect 44456 15376 44508 15428
rect 45284 15308 45336 15360
rect 52276 15580 52328 15632
rect 53104 15657 53113 15691
rect 53113 15657 53147 15691
rect 53147 15657 53156 15691
rect 53104 15648 53156 15657
rect 53012 15580 53064 15632
rect 47308 15555 47360 15564
rect 47308 15521 47317 15555
rect 47317 15521 47351 15555
rect 47351 15521 47360 15555
rect 47308 15512 47360 15521
rect 46848 15444 46900 15496
rect 49976 15444 50028 15496
rect 50068 15444 50120 15496
rect 52828 15512 52880 15564
rect 53564 15555 53616 15564
rect 53564 15521 53573 15555
rect 53573 15521 53607 15555
rect 53607 15521 53616 15555
rect 53564 15512 53616 15521
rect 56784 15555 56836 15564
rect 56784 15521 56793 15555
rect 56793 15521 56827 15555
rect 56827 15521 56836 15555
rect 56784 15512 56836 15521
rect 57888 15512 57940 15564
rect 52920 15487 52972 15496
rect 52920 15453 52929 15487
rect 52929 15453 52963 15487
rect 52963 15453 52972 15487
rect 52920 15444 52972 15453
rect 57060 15487 57112 15496
rect 57060 15453 57069 15487
rect 57069 15453 57103 15487
rect 57103 15453 57112 15487
rect 57060 15444 57112 15453
rect 48688 15308 48740 15360
rect 49700 15308 49752 15360
rect 50160 15308 50212 15360
rect 19574 15206 19626 15258
rect 19638 15206 19690 15258
rect 19702 15206 19754 15258
rect 19766 15206 19818 15258
rect 19830 15206 19882 15258
rect 50294 15206 50346 15258
rect 50358 15206 50410 15258
rect 50422 15206 50474 15258
rect 50486 15206 50538 15258
rect 50550 15206 50602 15258
rect 2688 15036 2740 15088
rect 3516 15036 3568 15088
rect 3792 15079 3844 15088
rect 3792 15045 3801 15079
rect 3801 15045 3835 15079
rect 3835 15045 3844 15079
rect 3792 15036 3844 15045
rect 2780 15011 2832 15020
rect 2780 14977 2789 15011
rect 2789 14977 2823 15011
rect 2823 14977 2832 15011
rect 2780 14968 2832 14977
rect 3424 14968 3476 15020
rect 3884 15011 3936 15020
rect 3884 14977 3893 15011
rect 3893 14977 3927 15011
rect 3927 14977 3936 15011
rect 3884 14968 3936 14977
rect 7748 15104 7800 15156
rect 9220 15147 9272 15156
rect 9220 15113 9229 15147
rect 9229 15113 9263 15147
rect 9263 15113 9272 15147
rect 9220 15104 9272 15113
rect 12348 15104 12400 15156
rect 14188 15104 14240 15156
rect 6644 15036 6696 15088
rect 10048 15079 10100 15088
rect 5816 15011 5868 15020
rect 5816 14977 5825 15011
rect 5825 14977 5859 15011
rect 5859 14977 5868 15011
rect 5816 14968 5868 14977
rect 4988 14832 5040 14884
rect 4712 14807 4764 14816
rect 4712 14773 4721 14807
rect 4721 14773 4755 14807
rect 4755 14773 4764 14807
rect 4712 14764 4764 14773
rect 7196 14968 7248 15020
rect 10048 15045 10057 15079
rect 10057 15045 10091 15079
rect 10091 15045 10100 15079
rect 10048 15036 10100 15045
rect 10140 14968 10192 15020
rect 10692 15011 10744 15020
rect 10692 14977 10701 15011
rect 10701 14977 10735 15011
rect 10735 14977 10744 15011
rect 10692 14968 10744 14977
rect 8944 14832 8996 14884
rect 10416 14832 10468 14884
rect 12072 15036 12124 15088
rect 19340 15104 19392 15156
rect 15016 15036 15068 15088
rect 11888 14968 11940 15020
rect 12440 15011 12492 15020
rect 12440 14977 12449 15011
rect 12449 14977 12483 15011
rect 12483 14977 12492 15011
rect 12440 14968 12492 14977
rect 12624 15011 12676 15020
rect 12624 14977 12633 15011
rect 12633 14977 12667 15011
rect 12667 14977 12676 15011
rect 12624 14968 12676 14977
rect 13452 14968 13504 15020
rect 15200 14968 15252 15020
rect 15568 15011 15620 15020
rect 15568 14977 15577 15011
rect 15577 14977 15611 15011
rect 15611 14977 15620 15011
rect 15568 14968 15620 14977
rect 12532 14832 12584 14884
rect 15476 14900 15528 14952
rect 15844 15079 15896 15088
rect 15844 15045 15853 15079
rect 15853 15045 15887 15079
rect 15887 15045 15896 15079
rect 15844 15036 15896 15045
rect 17960 15036 18012 15088
rect 17592 15011 17644 15020
rect 17592 14977 17601 15011
rect 17601 14977 17635 15011
rect 17635 14977 17644 15011
rect 17592 14968 17644 14977
rect 20076 15011 20128 15020
rect 20076 14977 20085 15011
rect 20085 14977 20119 15011
rect 20119 14977 20128 15011
rect 20076 14968 20128 14977
rect 20536 15104 20588 15156
rect 20720 15147 20772 15156
rect 20720 15113 20729 15147
rect 20729 15113 20763 15147
rect 20763 15113 20772 15147
rect 20720 15104 20772 15113
rect 23572 15104 23624 15156
rect 24216 15104 24268 15156
rect 20996 15036 21048 15088
rect 22100 15036 22152 15088
rect 23112 15036 23164 15088
rect 27620 15104 27672 15156
rect 28816 15104 28868 15156
rect 13360 14875 13412 14884
rect 13360 14841 13369 14875
rect 13369 14841 13403 14875
rect 13403 14841 13412 14875
rect 13360 14832 13412 14841
rect 14464 14875 14516 14884
rect 14464 14841 14473 14875
rect 14473 14841 14507 14875
rect 14507 14841 14516 14875
rect 14464 14832 14516 14841
rect 15844 14832 15896 14884
rect 15936 14832 15988 14884
rect 16856 14900 16908 14952
rect 17408 14900 17460 14952
rect 20536 15011 20588 15020
rect 20536 14977 20569 15011
rect 20569 14977 20588 15011
rect 20536 14968 20588 14977
rect 23296 14968 23348 15020
rect 25044 15036 25096 15088
rect 26240 15036 26292 15088
rect 20352 14900 20404 14952
rect 24768 15011 24820 15020
rect 24768 14977 24777 15011
rect 24777 14977 24811 15011
rect 24811 14977 24820 15011
rect 25872 15011 25924 15020
rect 24768 14968 24820 14977
rect 25872 14977 25881 15011
rect 25881 14977 25915 15011
rect 25915 14977 25924 15011
rect 25872 14968 25924 14977
rect 25596 14900 25648 14952
rect 26884 14968 26936 15020
rect 28080 15036 28132 15088
rect 38384 15147 38436 15156
rect 30932 15079 30984 15088
rect 28632 14968 28684 15020
rect 30012 14968 30064 15020
rect 30932 15045 30941 15079
rect 30941 15045 30975 15079
rect 30975 15045 30984 15079
rect 30932 15036 30984 15045
rect 30840 15011 30892 15020
rect 30840 14977 30849 15011
rect 30849 14977 30883 15011
rect 30883 14977 30892 15011
rect 31116 15011 31168 15020
rect 30840 14968 30892 14977
rect 31116 14977 31125 15011
rect 31125 14977 31159 15011
rect 31159 14977 31168 15011
rect 31116 14968 31168 14977
rect 17684 14875 17736 14884
rect 17684 14841 17693 14875
rect 17693 14841 17727 14875
rect 17727 14841 17736 14875
rect 17684 14832 17736 14841
rect 19524 14875 19576 14884
rect 19524 14841 19533 14875
rect 19533 14841 19567 14875
rect 19567 14841 19576 14875
rect 19524 14832 19576 14841
rect 20720 14832 20772 14884
rect 29000 14900 29052 14952
rect 10600 14764 10652 14816
rect 10968 14764 11020 14816
rect 11796 14764 11848 14816
rect 14648 14807 14700 14816
rect 14648 14773 14657 14807
rect 14657 14773 14691 14807
rect 14691 14773 14700 14807
rect 14648 14764 14700 14773
rect 15292 14764 15344 14816
rect 17224 14764 17276 14816
rect 20168 14764 20220 14816
rect 20536 14764 20588 14816
rect 23572 14807 23624 14816
rect 23572 14773 23581 14807
rect 23581 14773 23615 14807
rect 23615 14773 23624 14807
rect 23572 14764 23624 14773
rect 24124 14807 24176 14816
rect 24124 14773 24133 14807
rect 24133 14773 24167 14807
rect 24167 14773 24176 14807
rect 24124 14764 24176 14773
rect 30104 14943 30156 14952
rect 30104 14909 30113 14943
rect 30113 14909 30147 14943
rect 30147 14909 30156 14943
rect 32220 15036 32272 15088
rect 32036 14968 32088 15020
rect 33140 15036 33192 15088
rect 38384 15113 38393 15147
rect 38393 15113 38427 15147
rect 38427 15113 38436 15147
rect 38384 15104 38436 15113
rect 33508 15011 33560 15020
rect 30104 14900 30156 14909
rect 33508 14977 33517 15011
rect 33517 14977 33551 15011
rect 33551 14977 33560 15011
rect 33508 14968 33560 14977
rect 34336 15011 34388 15020
rect 34336 14977 34345 15011
rect 34345 14977 34379 15011
rect 34379 14977 34388 15011
rect 34336 14968 34388 14977
rect 37464 15011 37516 15020
rect 37464 14977 37473 15011
rect 37473 14977 37507 15011
rect 37507 14977 37516 15011
rect 37464 14968 37516 14977
rect 43260 15036 43312 15088
rect 44088 15036 44140 15088
rect 33324 14943 33376 14952
rect 32312 14832 32364 14884
rect 33324 14909 33333 14943
rect 33333 14909 33367 14943
rect 33367 14909 33376 14943
rect 33324 14900 33376 14909
rect 33876 14943 33928 14952
rect 33876 14909 33885 14943
rect 33885 14909 33919 14943
rect 33919 14909 33928 14943
rect 33876 14900 33928 14909
rect 40592 14968 40644 15020
rect 44180 14968 44232 15020
rect 38016 14900 38068 14952
rect 44364 15011 44416 15020
rect 44364 14977 44373 15011
rect 44373 14977 44407 15011
rect 44407 14977 44416 15011
rect 44364 14968 44416 14977
rect 45376 15011 45428 15020
rect 45376 14977 45385 15011
rect 45385 14977 45419 15011
rect 45419 14977 45428 15011
rect 45376 14968 45428 14977
rect 45928 14900 45980 14952
rect 33784 14875 33836 14884
rect 33784 14841 33793 14875
rect 33793 14841 33827 14875
rect 33827 14841 33836 14875
rect 33784 14832 33836 14841
rect 48688 15011 48740 15020
rect 30840 14764 30892 14816
rect 32036 14764 32088 14816
rect 34520 14764 34572 14816
rect 34612 14764 34664 14816
rect 36360 14764 36412 14816
rect 40776 14807 40828 14816
rect 40776 14773 40785 14807
rect 40785 14773 40819 14807
rect 40819 14773 40828 14807
rect 40776 14764 40828 14773
rect 44364 14764 44416 14816
rect 45376 14764 45428 14816
rect 45836 14764 45888 14816
rect 48688 14977 48697 15011
rect 48697 14977 48731 15011
rect 48731 14977 48740 15011
rect 48688 14968 48740 14977
rect 48780 14968 48832 15020
rect 50160 15104 50212 15156
rect 50252 15036 50304 15088
rect 56692 15104 56744 15156
rect 57428 15104 57480 15156
rect 52920 15036 52972 15088
rect 49700 15011 49752 15020
rect 48780 14832 48832 14884
rect 49700 14977 49709 15011
rect 49709 14977 49743 15011
rect 49743 14977 49752 15011
rect 49700 14968 49752 14977
rect 49976 14968 50028 15020
rect 50436 14968 50488 15020
rect 52552 14968 52604 15020
rect 53564 15036 53616 15088
rect 53380 14968 53432 15020
rect 56784 15011 56836 15020
rect 56784 14977 56793 15011
rect 56793 14977 56827 15011
rect 56827 14977 56836 15011
rect 56784 14968 56836 14977
rect 57060 14968 57112 15020
rect 57888 14968 57940 15020
rect 52276 14900 52328 14952
rect 50068 14832 50120 14884
rect 52828 14832 52880 14884
rect 53012 14875 53064 14884
rect 53012 14841 53021 14875
rect 53021 14841 53055 14875
rect 53055 14841 53064 14875
rect 53012 14832 53064 14841
rect 46848 14764 46900 14816
rect 50160 14764 50212 14816
rect 53196 14764 53248 14816
rect 54484 14764 54536 14816
rect 4214 14662 4266 14714
rect 4278 14662 4330 14714
rect 4342 14662 4394 14714
rect 4406 14662 4458 14714
rect 4470 14662 4522 14714
rect 34934 14662 34986 14714
rect 34998 14662 35050 14714
rect 35062 14662 35114 14714
rect 35126 14662 35178 14714
rect 35190 14662 35242 14714
rect 1492 14560 1544 14612
rect 3884 14560 3936 14612
rect 6920 14603 6972 14612
rect 6920 14569 6929 14603
rect 6929 14569 6963 14603
rect 6963 14569 6972 14603
rect 6920 14560 6972 14569
rect 10048 14560 10100 14612
rect 10784 14560 10836 14612
rect 12348 14560 12400 14612
rect 13452 14560 13504 14612
rect 14556 14560 14608 14612
rect 15844 14560 15896 14612
rect 16212 14560 16264 14612
rect 20076 14560 20128 14612
rect 20536 14560 20588 14612
rect 22284 14560 22336 14612
rect 26884 14560 26936 14612
rect 28448 14560 28500 14612
rect 30104 14560 30156 14612
rect 31024 14603 31076 14612
rect 31024 14569 31033 14603
rect 31033 14569 31067 14603
rect 31067 14569 31076 14603
rect 31024 14560 31076 14569
rect 32220 14560 32272 14612
rect 40040 14603 40092 14612
rect 40040 14569 40049 14603
rect 40049 14569 40083 14603
rect 40083 14569 40092 14603
rect 40040 14560 40092 14569
rect 14372 14492 14424 14544
rect 18420 14492 18472 14544
rect 8944 14424 8996 14476
rect 14096 14424 14148 14476
rect 14648 14424 14700 14476
rect 1400 14399 1452 14408
rect 1400 14365 1409 14399
rect 1409 14365 1443 14399
rect 1443 14365 1452 14399
rect 1400 14356 1452 14365
rect 10324 14356 10376 14408
rect 15568 14356 15620 14408
rect 15936 14399 15988 14408
rect 15936 14365 15945 14399
rect 15945 14365 15979 14399
rect 15979 14365 15988 14399
rect 15936 14356 15988 14365
rect 16672 14356 16724 14408
rect 17224 14399 17276 14408
rect 3516 14288 3568 14340
rect 6644 14288 6696 14340
rect 16028 14331 16080 14340
rect 16028 14297 16037 14331
rect 16037 14297 16071 14331
rect 16071 14297 16080 14331
rect 16028 14288 16080 14297
rect 4160 14220 4212 14272
rect 4712 14263 4764 14272
rect 4712 14229 4721 14263
rect 4721 14229 4755 14263
rect 4755 14229 4764 14263
rect 4712 14220 4764 14229
rect 5356 14220 5408 14272
rect 15016 14263 15068 14272
rect 15016 14229 15025 14263
rect 15025 14229 15059 14263
rect 15059 14229 15068 14263
rect 15016 14220 15068 14229
rect 17224 14365 17233 14399
rect 17233 14365 17267 14399
rect 17267 14365 17276 14399
rect 17224 14356 17276 14365
rect 17776 14356 17828 14408
rect 21824 14492 21876 14544
rect 20536 14424 20588 14476
rect 20812 14424 20864 14476
rect 20260 14399 20312 14408
rect 20260 14365 20269 14399
rect 20269 14365 20303 14399
rect 20303 14365 20312 14399
rect 20996 14399 21048 14408
rect 20260 14356 20312 14365
rect 20996 14365 21005 14399
rect 21005 14365 21039 14399
rect 21039 14365 21048 14399
rect 20996 14356 21048 14365
rect 21180 14399 21232 14408
rect 21180 14365 21189 14399
rect 21189 14365 21223 14399
rect 21223 14365 21232 14399
rect 21180 14356 21232 14365
rect 21640 14356 21692 14408
rect 17500 14331 17552 14340
rect 17500 14297 17509 14331
rect 17509 14297 17543 14331
rect 17543 14297 17552 14331
rect 17500 14288 17552 14297
rect 19432 14288 19484 14340
rect 27988 14424 28040 14476
rect 22008 14356 22060 14408
rect 24952 14399 25004 14408
rect 24952 14365 24961 14399
rect 24961 14365 24995 14399
rect 24995 14365 25004 14399
rect 24952 14356 25004 14365
rect 28080 14356 28132 14408
rect 28540 14399 28592 14408
rect 28540 14365 28549 14399
rect 28549 14365 28583 14399
rect 28583 14365 28592 14399
rect 28540 14356 28592 14365
rect 22376 14331 22428 14340
rect 22376 14297 22385 14331
rect 22385 14297 22419 14331
rect 22419 14297 22428 14331
rect 22376 14288 22428 14297
rect 24492 14288 24544 14340
rect 26332 14288 26384 14340
rect 28264 14331 28316 14340
rect 28264 14297 28273 14331
rect 28273 14297 28307 14331
rect 28307 14297 28316 14331
rect 28264 14288 28316 14297
rect 28356 14331 28408 14340
rect 28356 14297 28365 14331
rect 28365 14297 28399 14331
rect 28399 14297 28408 14331
rect 28816 14356 28868 14408
rect 31116 14492 31168 14544
rect 33876 14492 33928 14544
rect 30564 14356 30616 14408
rect 31484 14356 31536 14408
rect 32036 14399 32088 14408
rect 32036 14365 32045 14399
rect 32045 14365 32079 14399
rect 32079 14365 32088 14399
rect 32036 14356 32088 14365
rect 32128 14399 32180 14408
rect 32128 14365 32137 14399
rect 32137 14365 32171 14399
rect 32171 14365 32180 14399
rect 32128 14356 32180 14365
rect 32312 14399 32364 14408
rect 32312 14365 32321 14399
rect 32321 14365 32355 14399
rect 32355 14365 32364 14399
rect 33416 14424 33468 14476
rect 34612 14424 34664 14476
rect 32312 14356 32364 14365
rect 34980 14399 35032 14408
rect 34980 14365 34989 14399
rect 34989 14365 35023 14399
rect 35023 14365 35032 14399
rect 34980 14356 35032 14365
rect 43904 14492 43956 14544
rect 53012 14560 53064 14612
rect 53380 14603 53432 14612
rect 53380 14569 53389 14603
rect 53389 14569 53423 14603
rect 53423 14569 53432 14603
rect 53380 14560 53432 14569
rect 53564 14492 53616 14544
rect 28356 14288 28408 14297
rect 30932 14288 30984 14340
rect 21824 14263 21876 14272
rect 21824 14229 21833 14263
rect 21833 14229 21867 14263
rect 21867 14229 21876 14263
rect 21824 14220 21876 14229
rect 23664 14263 23716 14272
rect 23664 14229 23673 14263
rect 23673 14229 23707 14263
rect 23707 14229 23716 14263
rect 23664 14220 23716 14229
rect 27988 14263 28040 14272
rect 27988 14229 27997 14263
rect 27997 14229 28031 14263
rect 28031 14229 28040 14263
rect 27988 14220 28040 14229
rect 29644 14263 29696 14272
rect 29644 14229 29653 14263
rect 29653 14229 29687 14263
rect 29687 14229 29696 14263
rect 29644 14220 29696 14229
rect 31392 14220 31444 14272
rect 34520 14288 34572 14340
rect 32956 14220 33008 14272
rect 33324 14220 33376 14272
rect 33784 14220 33836 14272
rect 36360 14399 36412 14408
rect 36360 14365 36369 14399
rect 36369 14365 36403 14399
rect 36403 14365 36412 14399
rect 36360 14356 36412 14365
rect 37464 14356 37516 14408
rect 38016 14399 38068 14408
rect 38016 14365 38025 14399
rect 38025 14365 38059 14399
rect 38059 14365 38068 14399
rect 38016 14356 38068 14365
rect 38752 14288 38804 14340
rect 40040 14424 40092 14476
rect 44088 14467 44140 14476
rect 44088 14433 44097 14467
rect 44097 14433 44131 14467
rect 44131 14433 44140 14467
rect 44088 14424 44140 14433
rect 44272 14424 44324 14476
rect 45284 14424 45336 14476
rect 40776 14399 40828 14408
rect 40776 14365 40785 14399
rect 40785 14365 40819 14399
rect 40819 14365 40828 14399
rect 40776 14356 40828 14365
rect 43996 14399 44048 14408
rect 43996 14365 44005 14399
rect 44005 14365 44039 14399
rect 44039 14365 44048 14399
rect 43996 14356 44048 14365
rect 45836 14399 45888 14408
rect 45836 14365 45845 14399
rect 45845 14365 45879 14399
rect 45879 14365 45888 14399
rect 45836 14356 45888 14365
rect 45928 14399 45980 14408
rect 45928 14365 45937 14399
rect 45937 14365 45971 14399
rect 45971 14365 45980 14399
rect 52276 14424 52328 14476
rect 45928 14356 45980 14365
rect 50160 14399 50212 14408
rect 50160 14365 50169 14399
rect 50169 14365 50203 14399
rect 50203 14365 50212 14399
rect 50160 14356 50212 14365
rect 50252 14399 50304 14408
rect 50252 14365 50261 14399
rect 50261 14365 50295 14399
rect 50295 14365 50304 14399
rect 50252 14356 50304 14365
rect 50436 14399 50488 14408
rect 50436 14365 50445 14399
rect 50445 14365 50479 14399
rect 50479 14365 50488 14399
rect 50436 14356 50488 14365
rect 54484 14399 54536 14408
rect 54484 14365 54493 14399
rect 54493 14365 54527 14399
rect 54527 14365 54536 14399
rect 54484 14356 54536 14365
rect 56324 14424 56376 14476
rect 55496 14356 55548 14408
rect 38384 14220 38436 14272
rect 48780 14288 48832 14340
rect 55128 14288 55180 14340
rect 57336 14356 57388 14408
rect 42340 14220 42392 14272
rect 45008 14220 45060 14272
rect 46940 14220 46992 14272
rect 58072 14263 58124 14272
rect 58072 14229 58081 14263
rect 58081 14229 58115 14263
rect 58115 14229 58124 14263
rect 58072 14220 58124 14229
rect 19574 14118 19626 14170
rect 19638 14118 19690 14170
rect 19702 14118 19754 14170
rect 19766 14118 19818 14170
rect 19830 14118 19882 14170
rect 50294 14118 50346 14170
rect 50358 14118 50410 14170
rect 50422 14118 50474 14170
rect 50486 14118 50538 14170
rect 50550 14118 50602 14170
rect 16488 14016 16540 14068
rect 4160 13948 4212 14000
rect 12532 13991 12584 14000
rect 3516 13880 3568 13932
rect 9680 13880 9732 13932
rect 12532 13957 12541 13991
rect 12541 13957 12575 13991
rect 12575 13957 12584 13991
rect 14372 13991 14424 14000
rect 12532 13948 12584 13957
rect 14372 13957 14381 13991
rect 14381 13957 14415 13991
rect 14415 13957 14424 13991
rect 14372 13948 14424 13957
rect 15752 13991 15804 14000
rect 15752 13957 15761 13991
rect 15761 13957 15795 13991
rect 15795 13957 15804 13991
rect 15752 13948 15804 13957
rect 5356 13855 5408 13864
rect 5356 13821 5365 13855
rect 5365 13821 5399 13855
rect 5399 13821 5408 13855
rect 5356 13812 5408 13821
rect 7380 13812 7432 13864
rect 10968 13812 11020 13864
rect 4620 13787 4672 13796
rect 4620 13753 4629 13787
rect 4629 13753 4663 13787
rect 4663 13753 4672 13787
rect 4620 13744 4672 13753
rect 8852 13744 8904 13796
rect 14280 13880 14332 13932
rect 15568 13923 15620 13932
rect 15568 13889 15577 13923
rect 15577 13889 15611 13923
rect 15611 13889 15620 13923
rect 15568 13880 15620 13889
rect 15844 13923 15896 13932
rect 15844 13889 15853 13923
rect 15853 13889 15887 13923
rect 15887 13889 15896 13923
rect 15844 13880 15896 13889
rect 16212 13948 16264 14000
rect 16304 13948 16356 14000
rect 20812 13948 20864 14000
rect 22100 14016 22152 14068
rect 22376 14016 22428 14068
rect 23388 14016 23440 14068
rect 26240 14016 26292 14068
rect 26332 14016 26384 14068
rect 28632 14016 28684 14068
rect 29920 14016 29972 14068
rect 32312 14016 32364 14068
rect 38016 14016 38068 14068
rect 49792 14016 49844 14068
rect 50712 14016 50764 14068
rect 57888 14059 57940 14068
rect 57888 14025 57897 14059
rect 57897 14025 57931 14059
rect 57931 14025 57940 14059
rect 57888 14016 57940 14025
rect 16672 13923 16724 13932
rect 16672 13889 16681 13923
rect 16681 13889 16715 13923
rect 16715 13889 16724 13923
rect 16672 13880 16724 13889
rect 20168 13923 20220 13932
rect 20168 13889 20177 13923
rect 20177 13889 20211 13923
rect 20211 13889 20220 13923
rect 20168 13880 20220 13889
rect 20352 13880 20404 13932
rect 20904 13923 20956 13932
rect 20904 13889 20913 13923
rect 20913 13889 20947 13923
rect 20947 13889 20956 13923
rect 20904 13880 20956 13889
rect 21640 13948 21692 14000
rect 16948 13855 17000 13864
rect 13360 13719 13412 13728
rect 13360 13685 13369 13719
rect 13369 13685 13403 13719
rect 13403 13685 13412 13719
rect 13360 13676 13412 13685
rect 16948 13821 16957 13855
rect 16957 13821 16991 13855
rect 16991 13821 17000 13855
rect 16948 13812 17000 13821
rect 17868 13812 17920 13864
rect 20260 13812 20312 13864
rect 16120 13719 16172 13728
rect 16120 13685 16129 13719
rect 16129 13685 16163 13719
rect 16163 13685 16172 13719
rect 16120 13676 16172 13685
rect 20168 13744 20220 13796
rect 20996 13744 21048 13796
rect 21916 13923 21968 13932
rect 21916 13889 21926 13923
rect 21926 13889 21960 13923
rect 21960 13889 21968 13923
rect 21916 13880 21968 13889
rect 22836 13880 22888 13932
rect 22928 13880 22980 13932
rect 23664 13948 23716 14000
rect 27344 13948 27396 14000
rect 29000 13948 29052 14000
rect 29736 13948 29788 14000
rect 31116 13948 31168 14000
rect 33232 13948 33284 14000
rect 21364 13744 21416 13796
rect 24400 13880 24452 13932
rect 24768 13880 24820 13932
rect 30104 13880 30156 13932
rect 32496 13923 32548 13932
rect 32496 13889 32505 13923
rect 32505 13889 32539 13923
rect 32539 13889 32548 13923
rect 32496 13880 32548 13889
rect 32588 13923 32640 13932
rect 32588 13889 32597 13923
rect 32597 13889 32631 13923
rect 32631 13889 32640 13923
rect 32588 13880 32640 13889
rect 24952 13812 25004 13864
rect 28264 13812 28316 13864
rect 39120 13948 39172 14000
rect 45100 13948 45152 14000
rect 33784 13880 33836 13932
rect 34980 13923 35032 13932
rect 34980 13889 34989 13923
rect 34989 13889 35023 13923
rect 35023 13889 35032 13923
rect 34980 13880 35032 13889
rect 35808 13880 35860 13932
rect 37188 13880 37240 13932
rect 37372 13880 37424 13932
rect 38752 13880 38804 13932
rect 43904 13923 43956 13932
rect 43904 13889 43913 13923
rect 43913 13889 43947 13923
rect 43947 13889 43956 13923
rect 43904 13880 43956 13889
rect 43996 13923 44048 13932
rect 43996 13889 44005 13923
rect 44005 13889 44039 13923
rect 44039 13889 44048 13923
rect 53196 13923 53248 13932
rect 43996 13880 44048 13889
rect 53196 13889 53205 13923
rect 53205 13889 53239 13923
rect 53239 13889 53248 13923
rect 53196 13880 53248 13889
rect 55128 13880 55180 13932
rect 55496 13923 55548 13932
rect 55496 13889 55505 13923
rect 55505 13889 55539 13923
rect 55539 13889 55548 13923
rect 55496 13880 55548 13889
rect 56600 13923 56652 13932
rect 56600 13889 56609 13923
rect 56609 13889 56643 13923
rect 56643 13889 56652 13923
rect 56600 13880 56652 13889
rect 57888 13923 57940 13932
rect 57888 13889 57897 13923
rect 57897 13889 57931 13923
rect 57931 13889 57940 13923
rect 57888 13880 57940 13889
rect 34520 13812 34572 13864
rect 27804 13744 27856 13796
rect 22284 13676 22336 13728
rect 22468 13719 22520 13728
rect 22468 13685 22477 13719
rect 22477 13685 22511 13719
rect 22511 13685 22520 13719
rect 22468 13676 22520 13685
rect 23112 13719 23164 13728
rect 23112 13685 23121 13719
rect 23121 13685 23155 13719
rect 23155 13685 23164 13719
rect 23112 13676 23164 13685
rect 25136 13719 25188 13728
rect 25136 13685 25145 13719
rect 25145 13685 25179 13719
rect 25179 13685 25188 13719
rect 25136 13676 25188 13685
rect 32680 13719 32732 13728
rect 32680 13685 32689 13719
rect 32689 13685 32723 13719
rect 32723 13685 32732 13719
rect 32680 13676 32732 13685
rect 33232 13676 33284 13728
rect 34060 13676 34112 13728
rect 44088 13812 44140 13864
rect 53012 13855 53064 13864
rect 53012 13821 53021 13855
rect 53021 13821 53055 13855
rect 53055 13821 53064 13855
rect 53012 13812 53064 13821
rect 54484 13812 54536 13864
rect 56876 13855 56928 13864
rect 56876 13821 56885 13855
rect 56885 13821 56919 13855
rect 56919 13821 56928 13855
rect 56876 13812 56928 13821
rect 36176 13719 36228 13728
rect 36176 13685 36185 13719
rect 36185 13685 36219 13719
rect 36219 13685 36228 13719
rect 36176 13676 36228 13685
rect 40776 13676 40828 13728
rect 55404 13719 55456 13728
rect 55404 13685 55413 13719
rect 55413 13685 55447 13719
rect 55447 13685 55456 13719
rect 55404 13676 55456 13685
rect 56784 13676 56836 13728
rect 4214 13574 4266 13626
rect 4278 13574 4330 13626
rect 4342 13574 4394 13626
rect 4406 13574 4458 13626
rect 4470 13574 4522 13626
rect 34934 13574 34986 13626
rect 34998 13574 35050 13626
rect 35062 13574 35114 13626
rect 35126 13574 35178 13626
rect 35190 13574 35242 13626
rect 7932 13515 7984 13524
rect 7932 13481 7941 13515
rect 7941 13481 7975 13515
rect 7975 13481 7984 13515
rect 7932 13472 7984 13481
rect 9680 13515 9732 13524
rect 9680 13481 9689 13515
rect 9689 13481 9723 13515
rect 9723 13481 9732 13515
rect 9680 13472 9732 13481
rect 3240 13404 3292 13456
rect 9864 13404 9916 13456
rect 12348 13447 12400 13456
rect 12348 13413 12357 13447
rect 12357 13413 12391 13447
rect 12391 13413 12400 13447
rect 12348 13404 12400 13413
rect 15660 13472 15712 13524
rect 17500 13472 17552 13524
rect 3148 13311 3200 13320
rect 3148 13277 3157 13311
rect 3157 13277 3191 13311
rect 3191 13277 3200 13311
rect 3148 13268 3200 13277
rect 6368 13268 6420 13320
rect 7380 13311 7432 13320
rect 3056 13200 3108 13252
rect 6276 13200 6328 13252
rect 7380 13277 7389 13311
rect 7389 13277 7423 13311
rect 7423 13277 7432 13311
rect 7380 13268 7432 13277
rect 18236 13404 18288 13456
rect 20168 13404 20220 13456
rect 22836 13404 22888 13456
rect 23756 13447 23808 13456
rect 23756 13413 23765 13447
rect 23765 13413 23799 13447
rect 23799 13413 23808 13447
rect 23756 13404 23808 13413
rect 15384 13336 15436 13388
rect 14556 13311 14608 13320
rect 14556 13277 14565 13311
rect 14565 13277 14599 13311
rect 14599 13277 14608 13311
rect 14556 13268 14608 13277
rect 16028 13311 16080 13320
rect 16028 13277 16037 13311
rect 16037 13277 16071 13311
rect 16071 13277 16080 13311
rect 16028 13268 16080 13277
rect 16948 13268 17000 13320
rect 17408 13268 17460 13320
rect 17868 13311 17920 13320
rect 17868 13277 17877 13311
rect 17877 13277 17911 13311
rect 17911 13277 17920 13311
rect 17868 13268 17920 13277
rect 9680 13132 9732 13184
rect 10876 13132 10928 13184
rect 13084 13200 13136 13252
rect 13176 13200 13228 13252
rect 14832 13132 14884 13184
rect 15936 13200 15988 13252
rect 16304 13243 16356 13252
rect 16304 13209 16313 13243
rect 16313 13209 16347 13243
rect 16347 13209 16356 13243
rect 17776 13243 17828 13252
rect 16304 13200 16356 13209
rect 16672 13132 16724 13184
rect 17776 13209 17785 13243
rect 17785 13209 17819 13243
rect 17819 13209 17828 13243
rect 17776 13200 17828 13209
rect 21364 13336 21416 13388
rect 23112 13336 23164 13388
rect 19340 13268 19392 13320
rect 20536 13268 20588 13320
rect 22100 13311 22152 13320
rect 22100 13277 22109 13311
rect 22109 13277 22143 13311
rect 22143 13277 22152 13311
rect 22100 13268 22152 13277
rect 23020 13268 23072 13320
rect 19984 13243 20036 13252
rect 19984 13209 19993 13243
rect 19993 13209 20027 13243
rect 20027 13209 20036 13243
rect 19984 13200 20036 13209
rect 20352 13200 20404 13252
rect 22652 13200 22704 13252
rect 23296 13243 23348 13252
rect 23296 13209 23305 13243
rect 23305 13209 23339 13243
rect 23339 13209 23348 13243
rect 23296 13200 23348 13209
rect 22100 13132 22152 13184
rect 24124 13472 24176 13524
rect 30932 13472 30984 13524
rect 31116 13515 31168 13524
rect 31116 13481 31125 13515
rect 31125 13481 31159 13515
rect 31159 13481 31168 13515
rect 31116 13472 31168 13481
rect 31208 13472 31260 13524
rect 53196 13515 53248 13524
rect 53196 13481 53205 13515
rect 53205 13481 53239 13515
rect 53239 13481 53248 13515
rect 53196 13472 53248 13481
rect 56600 13472 56652 13524
rect 57888 13472 57940 13524
rect 24860 13311 24912 13320
rect 24860 13277 24869 13311
rect 24869 13277 24903 13311
rect 24903 13277 24912 13311
rect 24860 13268 24912 13277
rect 25044 13268 25096 13320
rect 25228 13311 25280 13320
rect 25228 13277 25237 13311
rect 25237 13277 25271 13311
rect 25271 13277 25280 13311
rect 25228 13268 25280 13277
rect 25596 13268 25648 13320
rect 26240 13311 26292 13320
rect 26240 13277 26249 13311
rect 26249 13277 26283 13311
rect 26283 13277 26292 13311
rect 26240 13268 26292 13277
rect 27804 13311 27856 13320
rect 27804 13277 27813 13311
rect 27813 13277 27847 13311
rect 27847 13277 27856 13311
rect 27804 13268 27856 13277
rect 27988 13268 28040 13320
rect 29644 13268 29696 13320
rect 30012 13268 30064 13320
rect 30196 13268 30248 13320
rect 32036 13268 32088 13320
rect 32588 13268 32640 13320
rect 24124 13200 24176 13252
rect 25136 13243 25188 13252
rect 25136 13209 25145 13243
rect 25145 13209 25179 13243
rect 25179 13209 25188 13243
rect 25136 13200 25188 13209
rect 28724 13200 28776 13252
rect 32128 13200 32180 13252
rect 32312 13243 32364 13252
rect 32312 13209 32321 13243
rect 32321 13209 32355 13243
rect 32355 13209 32364 13243
rect 32312 13200 32364 13209
rect 57796 13404 57848 13456
rect 41144 13336 41196 13388
rect 46756 13379 46808 13388
rect 46756 13345 46765 13379
rect 46765 13345 46799 13379
rect 46799 13345 46808 13379
rect 46756 13336 46808 13345
rect 50712 13379 50764 13388
rect 50712 13345 50721 13379
rect 50721 13345 50755 13379
rect 50755 13345 50764 13379
rect 50712 13336 50764 13345
rect 56876 13379 56928 13388
rect 56876 13345 56885 13379
rect 56885 13345 56919 13379
rect 56919 13345 56928 13379
rect 56876 13336 56928 13345
rect 36176 13268 36228 13320
rect 40776 13311 40828 13320
rect 40776 13277 40785 13311
rect 40785 13277 40819 13311
rect 40819 13277 40828 13311
rect 40776 13268 40828 13277
rect 42340 13311 42392 13320
rect 42340 13277 42349 13311
rect 42349 13277 42383 13311
rect 42383 13277 42392 13311
rect 42340 13268 42392 13277
rect 45008 13311 45060 13320
rect 37740 13200 37792 13252
rect 45008 13277 45017 13311
rect 45017 13277 45051 13311
rect 45051 13277 45060 13311
rect 45008 13268 45060 13277
rect 45100 13311 45152 13320
rect 45100 13277 45109 13311
rect 45109 13277 45143 13311
rect 45143 13277 45152 13311
rect 45100 13268 45152 13277
rect 45284 13311 45336 13320
rect 45284 13277 45293 13311
rect 45293 13277 45327 13311
rect 45327 13277 45336 13311
rect 46940 13311 46992 13320
rect 45284 13268 45336 13277
rect 46940 13277 46949 13311
rect 46949 13277 46983 13311
rect 46983 13277 46992 13311
rect 46940 13268 46992 13277
rect 48320 13311 48372 13320
rect 48320 13277 48329 13311
rect 48329 13277 48363 13311
rect 48363 13277 48372 13311
rect 48320 13268 48372 13277
rect 50804 13311 50856 13320
rect 27068 13175 27120 13184
rect 27068 13141 27077 13175
rect 27077 13141 27111 13175
rect 27111 13141 27120 13175
rect 27068 13132 27120 13141
rect 27252 13132 27304 13184
rect 29368 13132 29420 13184
rect 31760 13175 31812 13184
rect 31760 13141 31769 13175
rect 31769 13141 31803 13175
rect 31803 13141 31812 13175
rect 31760 13132 31812 13141
rect 32496 13132 32548 13184
rect 34796 13132 34848 13184
rect 37556 13132 37608 13184
rect 38476 13175 38528 13184
rect 38476 13141 38485 13175
rect 38485 13141 38519 13175
rect 38519 13141 38528 13175
rect 38476 13132 38528 13141
rect 42892 13200 42944 13252
rect 47952 13200 48004 13252
rect 50804 13277 50813 13311
rect 50813 13277 50847 13311
rect 50847 13277 50856 13311
rect 50804 13268 50856 13277
rect 53012 13311 53064 13320
rect 53012 13277 53021 13311
rect 53021 13277 53055 13311
rect 53055 13277 53064 13311
rect 53012 13268 53064 13277
rect 56784 13311 56836 13320
rect 56784 13277 56793 13311
rect 56793 13277 56827 13311
rect 56827 13277 56836 13311
rect 56784 13268 56836 13277
rect 43352 13175 43404 13184
rect 43352 13141 43361 13175
rect 43361 13141 43395 13175
rect 43395 13141 43404 13175
rect 43352 13132 43404 13141
rect 45468 13175 45520 13184
rect 45468 13141 45477 13175
rect 45477 13141 45511 13175
rect 45511 13141 45520 13175
rect 45468 13132 45520 13141
rect 51172 13175 51224 13184
rect 51172 13141 51181 13175
rect 51181 13141 51215 13175
rect 51215 13141 51224 13175
rect 51172 13132 51224 13141
rect 54484 13132 54536 13184
rect 19574 13030 19626 13082
rect 19638 13030 19690 13082
rect 19702 13030 19754 13082
rect 19766 13030 19818 13082
rect 19830 13030 19882 13082
rect 50294 13030 50346 13082
rect 50358 13030 50410 13082
rect 50422 13030 50474 13082
rect 50486 13030 50538 13082
rect 50550 13030 50602 13082
rect 1584 12971 1636 12980
rect 1584 12937 1593 12971
rect 1593 12937 1627 12971
rect 1627 12937 1636 12971
rect 1584 12928 1636 12937
rect 3056 12860 3108 12912
rect 3240 12860 3292 12912
rect 6368 12903 6420 12912
rect 1400 12835 1452 12844
rect 1400 12801 1409 12835
rect 1409 12801 1443 12835
rect 1443 12801 1452 12835
rect 1400 12792 1452 12801
rect 2872 12792 2924 12844
rect 2596 12767 2648 12776
rect 2596 12733 2605 12767
rect 2605 12733 2639 12767
rect 2639 12733 2648 12767
rect 2596 12724 2648 12733
rect 3056 12588 3108 12640
rect 6368 12869 6377 12903
rect 6377 12869 6411 12903
rect 6411 12869 6420 12903
rect 6368 12860 6420 12869
rect 6552 12835 6604 12844
rect 6552 12801 6561 12835
rect 6561 12801 6595 12835
rect 6595 12801 6604 12835
rect 6552 12792 6604 12801
rect 7288 12792 7340 12844
rect 8668 12792 8720 12844
rect 8852 12835 8904 12844
rect 8852 12801 8861 12835
rect 8861 12801 8895 12835
rect 8895 12801 8904 12835
rect 8852 12792 8904 12801
rect 9680 12860 9732 12912
rect 10968 12928 11020 12980
rect 13084 12971 13136 12980
rect 13084 12937 13093 12971
rect 13093 12937 13127 12971
rect 13127 12937 13136 12971
rect 13084 12928 13136 12937
rect 14924 12971 14976 12980
rect 14924 12937 14933 12971
rect 14933 12937 14967 12971
rect 14967 12937 14976 12971
rect 14924 12928 14976 12937
rect 15108 12928 15160 12980
rect 11980 12792 12032 12844
rect 15660 12860 15712 12912
rect 16120 12860 16172 12912
rect 12716 12792 12768 12844
rect 13176 12835 13228 12844
rect 13176 12801 13185 12835
rect 13185 12801 13219 12835
rect 13219 12801 13228 12835
rect 13176 12792 13228 12801
rect 14740 12792 14792 12844
rect 15844 12792 15896 12844
rect 16672 12835 16724 12844
rect 16672 12801 16681 12835
rect 16681 12801 16715 12835
rect 16715 12801 16724 12835
rect 16672 12792 16724 12801
rect 17776 12860 17828 12912
rect 19340 12928 19392 12980
rect 19432 12928 19484 12980
rect 20076 12928 20128 12980
rect 23296 12928 23348 12980
rect 24032 12860 24084 12912
rect 17960 12792 18012 12844
rect 18880 12835 18932 12844
rect 18880 12801 18889 12835
rect 18889 12801 18923 12835
rect 18923 12801 18932 12835
rect 18880 12792 18932 12801
rect 12440 12724 12492 12776
rect 16028 12724 16080 12776
rect 17040 12724 17092 12776
rect 18512 12724 18564 12776
rect 20076 12792 20128 12844
rect 24676 12903 24728 12912
rect 24676 12869 24685 12903
rect 24685 12869 24719 12903
rect 24719 12869 24728 12903
rect 24676 12860 24728 12869
rect 24860 12928 24912 12980
rect 27068 12928 27120 12980
rect 37188 12928 37240 12980
rect 37556 12928 37608 12980
rect 43352 12928 43404 12980
rect 24492 12835 24544 12844
rect 24492 12801 24501 12835
rect 24501 12801 24535 12835
rect 24535 12801 24544 12835
rect 24768 12835 24820 12844
rect 24492 12792 24544 12801
rect 24768 12801 24777 12835
rect 24777 12801 24811 12835
rect 24811 12801 24820 12835
rect 24768 12792 24820 12801
rect 24952 12792 25004 12844
rect 25596 12835 25648 12844
rect 25596 12801 25605 12835
rect 25605 12801 25639 12835
rect 25639 12801 25648 12835
rect 25596 12792 25648 12801
rect 28540 12792 28592 12844
rect 29184 12792 29236 12844
rect 29368 12835 29420 12844
rect 29368 12801 29377 12835
rect 29377 12801 29411 12835
rect 29411 12801 29420 12835
rect 29368 12792 29420 12801
rect 30564 12835 30616 12844
rect 30564 12801 30573 12835
rect 30573 12801 30607 12835
rect 30607 12801 30616 12835
rect 30564 12792 30616 12801
rect 20352 12724 20404 12776
rect 25044 12724 25096 12776
rect 27436 12724 27488 12776
rect 28172 12724 28224 12776
rect 28816 12724 28868 12776
rect 32036 12792 32088 12844
rect 32312 12835 32364 12844
rect 32312 12801 32321 12835
rect 32321 12801 32355 12835
rect 32355 12801 32364 12835
rect 32312 12792 32364 12801
rect 37740 12835 37792 12844
rect 37740 12801 37749 12835
rect 37749 12801 37783 12835
rect 37783 12801 37792 12835
rect 37740 12792 37792 12801
rect 38752 12860 38804 12912
rect 42892 12903 42944 12912
rect 42892 12869 42901 12903
rect 42901 12869 42935 12903
rect 42935 12869 42944 12903
rect 42892 12860 42944 12869
rect 45100 12860 45152 12912
rect 48320 12928 48372 12980
rect 50712 12928 50764 12980
rect 54484 12971 54536 12980
rect 54484 12937 54493 12971
rect 54493 12937 54527 12971
rect 54527 12937 54536 12971
rect 54484 12928 54536 12937
rect 32496 12724 32548 12776
rect 32680 12724 32732 12776
rect 33140 12724 33192 12776
rect 25780 12699 25832 12708
rect 25780 12665 25789 12699
rect 25789 12665 25823 12699
rect 25823 12665 25832 12699
rect 25780 12656 25832 12665
rect 29460 12656 29512 12708
rect 38476 12656 38528 12708
rect 40776 12792 40828 12844
rect 45008 12835 45060 12844
rect 41144 12767 41196 12776
rect 41144 12733 41153 12767
rect 41153 12733 41187 12767
rect 41187 12733 41196 12767
rect 41144 12724 41196 12733
rect 42340 12656 42392 12708
rect 45008 12801 45017 12835
rect 45017 12801 45051 12835
rect 45051 12801 45060 12835
rect 45008 12792 45060 12801
rect 55036 12928 55088 12980
rect 55404 12928 55456 12980
rect 45284 12792 45336 12844
rect 46756 12835 46808 12844
rect 46756 12801 46765 12835
rect 46765 12801 46799 12835
rect 46799 12801 46808 12835
rect 46756 12792 46808 12801
rect 46848 12792 46900 12844
rect 47952 12835 48004 12844
rect 47952 12801 47961 12835
rect 47961 12801 47995 12835
rect 47995 12801 48004 12835
rect 50804 12835 50856 12844
rect 47952 12792 48004 12801
rect 50804 12801 50813 12835
rect 50813 12801 50847 12835
rect 50847 12801 50856 12835
rect 50804 12792 50856 12801
rect 51172 12792 51224 12844
rect 51448 12792 51500 12844
rect 55036 12835 55088 12844
rect 55036 12801 55045 12835
rect 55045 12801 55079 12835
rect 55079 12801 55088 12835
rect 55036 12792 55088 12801
rect 46112 12724 46164 12776
rect 51632 12767 51684 12776
rect 51632 12733 51641 12767
rect 51641 12733 51675 12767
rect 51675 12733 51684 12767
rect 51632 12724 51684 12733
rect 52552 12656 52604 12708
rect 54484 12724 54536 12776
rect 5908 12588 5960 12640
rect 7840 12631 7892 12640
rect 7840 12597 7849 12631
rect 7849 12597 7883 12631
rect 7883 12597 7892 12631
rect 7840 12588 7892 12597
rect 10876 12631 10928 12640
rect 10876 12597 10885 12631
rect 10885 12597 10919 12631
rect 10919 12597 10928 12631
rect 10876 12588 10928 12597
rect 18880 12588 18932 12640
rect 23020 12631 23072 12640
rect 23020 12597 23029 12631
rect 23029 12597 23063 12631
rect 23063 12597 23072 12631
rect 23020 12588 23072 12597
rect 30656 12588 30708 12640
rect 38292 12588 38344 12640
rect 38752 12631 38804 12640
rect 38752 12597 38761 12631
rect 38761 12597 38795 12631
rect 38795 12597 38804 12631
rect 38752 12588 38804 12597
rect 49056 12588 49108 12640
rect 51724 12631 51776 12640
rect 51724 12597 51733 12631
rect 51733 12597 51767 12631
rect 51767 12597 51776 12631
rect 51724 12588 51776 12597
rect 52460 12588 52512 12640
rect 56600 12792 56652 12844
rect 56784 12860 56836 12912
rect 56876 12792 56928 12844
rect 56140 12724 56192 12776
rect 4214 12486 4266 12538
rect 4278 12486 4330 12538
rect 4342 12486 4394 12538
rect 4406 12486 4458 12538
rect 4470 12486 4522 12538
rect 34934 12486 34986 12538
rect 34998 12486 35050 12538
rect 35062 12486 35114 12538
rect 35126 12486 35178 12538
rect 35190 12486 35242 12538
rect 3148 12384 3200 12436
rect 5908 12427 5960 12436
rect 1400 12359 1452 12368
rect 1400 12325 1409 12359
rect 1409 12325 1443 12359
rect 1443 12325 1452 12359
rect 1400 12316 1452 12325
rect 4252 12223 4304 12232
rect 4252 12189 4261 12223
rect 4261 12189 4295 12223
rect 4295 12189 4304 12223
rect 4252 12180 4304 12189
rect 5908 12393 5917 12427
rect 5917 12393 5951 12427
rect 5951 12393 5960 12427
rect 5908 12384 5960 12393
rect 8668 12384 8720 12436
rect 10416 12316 10468 12368
rect 6552 12248 6604 12300
rect 8852 12248 8904 12300
rect 12440 12248 12492 12300
rect 13544 12316 13596 12368
rect 5724 12112 5776 12164
rect 6184 12155 6236 12164
rect 6184 12121 6193 12155
rect 6193 12121 6227 12155
rect 6227 12121 6236 12155
rect 6184 12112 6236 12121
rect 6460 12223 6512 12232
rect 6460 12189 6469 12223
rect 6469 12189 6503 12223
rect 6503 12189 6512 12223
rect 7104 12223 7156 12232
rect 6460 12180 6512 12189
rect 7104 12189 7113 12223
rect 7113 12189 7147 12223
rect 7147 12189 7156 12223
rect 8024 12223 8076 12232
rect 7104 12180 7156 12189
rect 7288 12155 7340 12164
rect 7288 12121 7297 12155
rect 7297 12121 7331 12155
rect 7331 12121 7340 12155
rect 7288 12112 7340 12121
rect 8024 12189 8033 12223
rect 8033 12189 8067 12223
rect 8067 12189 8076 12223
rect 8024 12180 8076 12189
rect 8944 12180 8996 12232
rect 9864 12180 9916 12232
rect 17132 12384 17184 12436
rect 21180 12384 21232 12436
rect 22652 12384 22704 12436
rect 19340 12316 19392 12368
rect 21088 12316 21140 12368
rect 9680 12112 9732 12164
rect 15108 12180 15160 12232
rect 15568 12180 15620 12232
rect 15752 12112 15804 12164
rect 16212 12112 16264 12164
rect 10232 12044 10284 12096
rect 11888 12044 11940 12096
rect 15660 12044 15712 12096
rect 16488 12087 16540 12096
rect 16488 12053 16497 12087
rect 16497 12053 16531 12087
rect 16531 12053 16540 12087
rect 16488 12044 16540 12053
rect 17040 12223 17092 12232
rect 17040 12189 17049 12223
rect 17049 12189 17083 12223
rect 17083 12189 17092 12223
rect 17040 12180 17092 12189
rect 19432 12223 19484 12232
rect 19432 12189 19441 12223
rect 19441 12189 19475 12223
rect 19475 12189 19484 12223
rect 19432 12180 19484 12189
rect 16764 12155 16816 12164
rect 16764 12121 16773 12155
rect 16773 12121 16807 12155
rect 16807 12121 16816 12155
rect 16764 12112 16816 12121
rect 17132 12112 17184 12164
rect 17776 12112 17828 12164
rect 18788 12112 18840 12164
rect 17592 12044 17644 12096
rect 18512 12087 18564 12096
rect 18512 12053 18521 12087
rect 18521 12053 18555 12087
rect 18555 12053 18564 12087
rect 18512 12044 18564 12053
rect 19248 12087 19300 12096
rect 19248 12053 19257 12087
rect 19257 12053 19291 12087
rect 19291 12053 19300 12087
rect 19248 12044 19300 12053
rect 20168 12223 20220 12232
rect 20168 12189 20177 12223
rect 20177 12189 20211 12223
rect 20211 12189 20220 12223
rect 20352 12223 20404 12232
rect 20168 12180 20220 12189
rect 20352 12189 20361 12223
rect 20361 12189 20395 12223
rect 20395 12189 20404 12223
rect 20352 12180 20404 12189
rect 21180 12180 21232 12232
rect 20628 12155 20680 12164
rect 20628 12121 20637 12155
rect 20637 12121 20671 12155
rect 20671 12121 20680 12155
rect 20628 12112 20680 12121
rect 20996 12112 21048 12164
rect 21456 12155 21508 12164
rect 21456 12121 21465 12155
rect 21465 12121 21499 12155
rect 21499 12121 21508 12155
rect 22100 12180 22152 12232
rect 22376 12223 22428 12232
rect 22376 12189 22385 12223
rect 22385 12189 22419 12223
rect 22419 12189 22428 12223
rect 22376 12180 22428 12189
rect 22468 12180 22520 12232
rect 24216 12180 24268 12232
rect 24676 12180 24728 12232
rect 25688 12180 25740 12232
rect 30196 12384 30248 12436
rect 30288 12384 30340 12436
rect 32496 12427 32548 12436
rect 28816 12316 28868 12368
rect 28632 12248 28684 12300
rect 30656 12316 30708 12368
rect 32496 12393 32505 12427
rect 32505 12393 32539 12427
rect 32539 12393 32548 12427
rect 32496 12384 32548 12393
rect 34796 12384 34848 12436
rect 37556 12427 37608 12436
rect 37556 12393 37565 12427
rect 37565 12393 37599 12427
rect 37599 12393 37608 12427
rect 37556 12384 37608 12393
rect 21456 12112 21508 12121
rect 21916 12112 21968 12164
rect 21272 12044 21324 12096
rect 29644 12180 29696 12232
rect 30012 12248 30064 12300
rect 30104 12223 30156 12232
rect 30104 12189 30113 12223
rect 30113 12189 30147 12223
rect 30147 12189 30156 12223
rect 30104 12180 30156 12189
rect 34520 12248 34572 12300
rect 30840 12223 30892 12232
rect 30840 12189 30849 12223
rect 30849 12189 30883 12223
rect 30883 12189 30892 12223
rect 30840 12180 30892 12189
rect 31760 12180 31812 12232
rect 29920 12155 29972 12164
rect 25780 12044 25832 12096
rect 29920 12121 29929 12155
rect 29929 12121 29963 12155
rect 29963 12121 29972 12155
rect 29920 12112 29972 12121
rect 34704 12155 34756 12164
rect 34704 12121 34713 12155
rect 34713 12121 34747 12155
rect 34747 12121 34756 12155
rect 34704 12112 34756 12121
rect 38752 12248 38804 12300
rect 38292 12223 38344 12232
rect 38292 12189 38301 12223
rect 38301 12189 38335 12223
rect 38335 12189 38344 12223
rect 38292 12180 38344 12189
rect 37188 12112 37240 12164
rect 38384 12112 38436 12164
rect 40684 12180 40736 12232
rect 41144 12223 41196 12232
rect 41144 12189 41153 12223
rect 41153 12189 41187 12223
rect 41187 12189 41196 12223
rect 41144 12180 41196 12189
rect 45744 12223 45796 12232
rect 45744 12189 45753 12223
rect 45753 12189 45787 12223
rect 45787 12189 45796 12223
rect 45744 12180 45796 12189
rect 48596 12223 48648 12232
rect 48596 12189 48605 12223
rect 48605 12189 48639 12223
rect 48639 12189 48648 12223
rect 48596 12180 48648 12189
rect 51724 12248 51776 12300
rect 49056 12223 49108 12232
rect 43812 12112 43864 12164
rect 45376 12112 45428 12164
rect 49056 12189 49065 12223
rect 49065 12189 49099 12223
rect 49099 12189 49108 12223
rect 49056 12180 49108 12189
rect 51448 12223 51500 12232
rect 51448 12189 51457 12223
rect 51457 12189 51491 12223
rect 51491 12189 51500 12223
rect 51448 12180 51500 12189
rect 51632 12180 51684 12232
rect 52460 12180 52512 12232
rect 56508 12180 56560 12232
rect 57152 12180 57204 12232
rect 57796 12248 57848 12300
rect 58164 12223 58216 12232
rect 58164 12189 58173 12223
rect 58173 12189 58207 12223
rect 58207 12189 58216 12223
rect 58164 12180 58216 12189
rect 48964 12112 49016 12164
rect 51172 12155 51224 12164
rect 51172 12121 51181 12155
rect 51181 12121 51215 12155
rect 51215 12121 51224 12155
rect 51908 12155 51960 12164
rect 51172 12112 51224 12121
rect 51908 12121 51917 12155
rect 51917 12121 51951 12155
rect 51951 12121 51960 12155
rect 51908 12112 51960 12121
rect 56232 12155 56284 12164
rect 56232 12121 56241 12155
rect 56241 12121 56275 12155
rect 56275 12121 56284 12155
rect 56232 12112 56284 12121
rect 30748 12044 30800 12096
rect 31944 12087 31996 12096
rect 31944 12053 31953 12087
rect 31953 12053 31987 12087
rect 31987 12053 31996 12087
rect 31944 12044 31996 12053
rect 33784 12044 33836 12096
rect 35348 12044 35400 12096
rect 43168 12044 43220 12096
rect 43720 12044 43772 12096
rect 45836 12087 45888 12096
rect 45836 12053 45845 12087
rect 45845 12053 45879 12087
rect 45879 12053 45888 12087
rect 45836 12044 45888 12053
rect 56600 12087 56652 12096
rect 56600 12053 56609 12087
rect 56609 12053 56643 12087
rect 56643 12053 56652 12087
rect 56600 12044 56652 12053
rect 57060 12087 57112 12096
rect 57060 12053 57069 12087
rect 57069 12053 57103 12087
rect 57103 12053 57112 12087
rect 57060 12044 57112 12053
rect 19574 11942 19626 11994
rect 19638 11942 19690 11994
rect 19702 11942 19754 11994
rect 19766 11942 19818 11994
rect 19830 11942 19882 11994
rect 50294 11942 50346 11994
rect 50358 11942 50410 11994
rect 50422 11942 50474 11994
rect 50486 11942 50538 11994
rect 50550 11942 50602 11994
rect 4252 11840 4304 11892
rect 5724 11840 5776 11892
rect 7288 11840 7340 11892
rect 8944 11883 8996 11892
rect 8944 11849 8953 11883
rect 8953 11849 8987 11883
rect 8987 11849 8996 11883
rect 8944 11840 8996 11849
rect 17316 11840 17368 11892
rect 18788 11883 18840 11892
rect 18788 11849 18797 11883
rect 18797 11849 18831 11883
rect 18831 11849 18840 11883
rect 18788 11840 18840 11849
rect 19340 11883 19392 11892
rect 19340 11849 19349 11883
rect 19349 11849 19383 11883
rect 19383 11849 19392 11883
rect 19340 11840 19392 11849
rect 20168 11840 20220 11892
rect 3240 11704 3292 11756
rect 3608 11772 3660 11824
rect 3792 11704 3844 11756
rect 3884 11747 3936 11756
rect 3884 11713 3893 11747
rect 3893 11713 3927 11747
rect 3927 11713 3936 11747
rect 3884 11704 3936 11713
rect 6184 11704 6236 11756
rect 6368 11747 6420 11756
rect 6368 11713 6377 11747
rect 6377 11713 6411 11747
rect 6411 11713 6420 11747
rect 6368 11704 6420 11713
rect 7104 11704 7156 11756
rect 9680 11772 9732 11824
rect 10048 11772 10100 11824
rect 12624 11772 12676 11824
rect 9312 11747 9364 11756
rect 8024 11636 8076 11688
rect 9312 11713 9321 11747
rect 9321 11713 9355 11747
rect 9355 11713 9364 11747
rect 9312 11704 9364 11713
rect 11888 11747 11940 11756
rect 11888 11713 11897 11747
rect 11897 11713 11931 11747
rect 11931 11713 11940 11747
rect 11888 11704 11940 11713
rect 12348 11747 12400 11756
rect 12348 11713 12357 11747
rect 12357 11713 12391 11747
rect 12391 11713 12400 11747
rect 12348 11704 12400 11713
rect 15384 11747 15436 11756
rect 15384 11713 15393 11747
rect 15393 11713 15427 11747
rect 15427 11713 15436 11747
rect 15384 11704 15436 11713
rect 16304 11772 16356 11824
rect 21272 11840 21324 11892
rect 15660 11747 15712 11756
rect 15660 11713 15669 11747
rect 15669 11713 15703 11747
rect 15703 11713 15712 11747
rect 15660 11704 15712 11713
rect 16488 11704 16540 11756
rect 10232 11636 10284 11688
rect 16120 11636 16172 11688
rect 21456 11772 21508 11824
rect 23572 11772 23624 11824
rect 16672 11704 16724 11756
rect 16948 11747 17000 11756
rect 16948 11713 16957 11747
rect 16957 11713 16991 11747
rect 16991 11713 17000 11747
rect 16948 11704 17000 11713
rect 17132 11704 17184 11756
rect 19340 11704 19392 11756
rect 20444 11704 20496 11756
rect 22284 11704 22336 11756
rect 22652 11747 22704 11756
rect 22100 11636 22152 11688
rect 22652 11713 22661 11747
rect 22661 11713 22695 11747
rect 22695 11713 22704 11747
rect 22652 11704 22704 11713
rect 22836 11747 22888 11756
rect 22836 11713 22850 11747
rect 22850 11713 22884 11747
rect 22884 11713 22888 11747
rect 22836 11704 22888 11713
rect 23664 11704 23716 11756
rect 24492 11704 24544 11756
rect 24952 11704 25004 11756
rect 25780 11815 25832 11824
rect 25780 11781 25789 11815
rect 25789 11781 25823 11815
rect 25823 11781 25832 11815
rect 25780 11772 25832 11781
rect 27804 11772 27856 11824
rect 28264 11772 28316 11824
rect 23940 11636 23992 11688
rect 25228 11636 25280 11688
rect 25964 11747 26016 11756
rect 25964 11713 25973 11747
rect 25973 11713 26007 11747
rect 26007 11713 26016 11747
rect 25964 11704 26016 11713
rect 27620 11704 27672 11756
rect 28172 11747 28224 11756
rect 28172 11713 28181 11747
rect 28181 11713 28215 11747
rect 28215 11713 28224 11747
rect 28172 11704 28224 11713
rect 29644 11840 29696 11892
rect 30104 11840 30156 11892
rect 32496 11840 32548 11892
rect 29184 11747 29236 11756
rect 6460 11568 6512 11620
rect 7104 11611 7156 11620
rect 7104 11577 7113 11611
rect 7113 11577 7147 11611
rect 7147 11577 7156 11611
rect 7104 11568 7156 11577
rect 14832 11568 14884 11620
rect 15108 11568 15160 11620
rect 18512 11568 18564 11620
rect 3700 11500 3752 11552
rect 9864 11543 9916 11552
rect 9864 11509 9873 11543
rect 9873 11509 9907 11543
rect 9907 11509 9916 11543
rect 9864 11500 9916 11509
rect 13176 11500 13228 11552
rect 15844 11500 15896 11552
rect 21088 11543 21140 11552
rect 21088 11509 21097 11543
rect 21097 11509 21131 11543
rect 21131 11509 21140 11543
rect 21088 11500 21140 11509
rect 23020 11543 23072 11552
rect 23020 11509 23029 11543
rect 23029 11509 23063 11543
rect 23063 11509 23072 11543
rect 23020 11500 23072 11509
rect 23296 11568 23348 11620
rect 25596 11568 25648 11620
rect 25320 11500 25372 11552
rect 27988 11636 28040 11688
rect 29184 11713 29193 11747
rect 29193 11713 29227 11747
rect 29227 11713 29236 11747
rect 29184 11704 29236 11713
rect 29644 11704 29696 11756
rect 30656 11772 30708 11824
rect 33692 11840 33744 11892
rect 34796 11840 34848 11892
rect 45376 11883 45428 11892
rect 33600 11815 33652 11824
rect 33600 11781 33609 11815
rect 33609 11781 33643 11815
rect 33643 11781 33652 11815
rect 33600 11772 33652 11781
rect 36268 11772 36320 11824
rect 38292 11772 38344 11824
rect 38752 11772 38804 11824
rect 45376 11849 45385 11883
rect 45385 11849 45419 11883
rect 45419 11849 45428 11883
rect 45376 11840 45428 11849
rect 51172 11840 51224 11892
rect 58164 11883 58216 11892
rect 58164 11849 58173 11883
rect 58173 11849 58207 11883
rect 58207 11849 58216 11883
rect 58164 11840 58216 11849
rect 43076 11772 43128 11824
rect 43720 11815 43772 11824
rect 29920 11704 29972 11756
rect 30196 11747 30248 11756
rect 30196 11713 30205 11747
rect 30205 11713 30239 11747
rect 30239 11713 30248 11747
rect 30196 11704 30248 11713
rect 34520 11747 34572 11756
rect 34520 11713 34529 11747
rect 34529 11713 34563 11747
rect 34563 11713 34572 11747
rect 34520 11704 34572 11713
rect 34704 11704 34756 11756
rect 36084 11704 36136 11756
rect 38384 11747 38436 11756
rect 38384 11713 38393 11747
rect 38393 11713 38427 11747
rect 38427 11713 38436 11747
rect 38384 11704 38436 11713
rect 39120 11747 39172 11756
rect 39120 11713 39129 11747
rect 39129 11713 39163 11747
rect 39163 11713 39172 11747
rect 39120 11704 39172 11713
rect 43168 11747 43220 11756
rect 43168 11713 43177 11747
rect 43177 11713 43211 11747
rect 43211 11713 43220 11747
rect 43168 11704 43220 11713
rect 43720 11781 43729 11815
rect 43729 11781 43763 11815
rect 43763 11781 43772 11815
rect 43720 11772 43772 11781
rect 43812 11747 43864 11756
rect 43812 11713 43821 11747
rect 43821 11713 43855 11747
rect 43855 11713 43864 11747
rect 43812 11704 43864 11713
rect 45468 11704 45520 11756
rect 46112 11747 46164 11756
rect 46112 11713 46121 11747
rect 46121 11713 46155 11747
rect 46155 11713 46164 11747
rect 46112 11704 46164 11713
rect 54668 11772 54720 11824
rect 56232 11772 56284 11824
rect 49056 11704 49108 11756
rect 53840 11704 53892 11756
rect 56048 11747 56100 11756
rect 56048 11713 56057 11747
rect 56057 11713 56091 11747
rect 56091 11713 56100 11747
rect 56048 11704 56100 11713
rect 56692 11747 56744 11756
rect 56692 11713 56701 11747
rect 56701 11713 56735 11747
rect 56735 11713 56744 11747
rect 56692 11704 56744 11713
rect 57152 11704 57204 11756
rect 30564 11636 30616 11688
rect 44916 11679 44968 11688
rect 44916 11645 44925 11679
rect 44925 11645 44959 11679
rect 44959 11645 44968 11679
rect 44916 11636 44968 11645
rect 45928 11679 45980 11688
rect 45928 11645 45937 11679
rect 45937 11645 45971 11679
rect 45971 11645 45980 11679
rect 45928 11636 45980 11645
rect 38476 11568 38528 11620
rect 27620 11500 27672 11552
rect 29368 11500 29420 11552
rect 31484 11500 31536 11552
rect 33784 11543 33836 11552
rect 33784 11509 33793 11543
rect 33793 11509 33827 11543
rect 33827 11509 33836 11543
rect 33784 11500 33836 11509
rect 34704 11500 34756 11552
rect 35440 11500 35492 11552
rect 39304 11543 39356 11552
rect 39304 11509 39313 11543
rect 39313 11509 39347 11543
rect 39347 11509 39356 11543
rect 39304 11500 39356 11509
rect 39856 11500 39908 11552
rect 48596 11636 48648 11688
rect 48964 11636 49016 11688
rect 56600 11679 56652 11688
rect 56600 11645 56609 11679
rect 56609 11645 56643 11679
rect 56643 11645 56652 11679
rect 56600 11636 56652 11645
rect 47952 11500 48004 11552
rect 53288 11543 53340 11552
rect 53288 11509 53297 11543
rect 53297 11509 53331 11543
rect 53331 11509 53340 11543
rect 53288 11500 53340 11509
rect 4214 11398 4266 11450
rect 4278 11398 4330 11450
rect 4342 11398 4394 11450
rect 4406 11398 4458 11450
rect 4470 11398 4522 11450
rect 34934 11398 34986 11450
rect 34998 11398 35050 11450
rect 35062 11398 35114 11450
rect 35126 11398 35178 11450
rect 35190 11398 35242 11450
rect 2872 11339 2924 11348
rect 2872 11305 2881 11339
rect 2881 11305 2915 11339
rect 2915 11305 2924 11339
rect 2872 11296 2924 11305
rect 3608 11296 3660 11348
rect 22284 11339 22336 11348
rect 22284 11305 22293 11339
rect 22293 11305 22327 11339
rect 22327 11305 22336 11339
rect 22284 11296 22336 11305
rect 22376 11296 22428 11348
rect 25596 11296 25648 11348
rect 30380 11296 30432 11348
rect 2872 11092 2924 11144
rect 3884 11160 3936 11212
rect 11888 11160 11940 11212
rect 4068 11092 4120 11144
rect 12348 11092 12400 11144
rect 15108 11092 15160 11144
rect 15844 11135 15896 11144
rect 15844 11101 15853 11135
rect 15853 11101 15887 11135
rect 15887 11101 15896 11135
rect 15844 11092 15896 11101
rect 14280 11024 14332 11076
rect 15200 11024 15252 11076
rect 16396 11160 16448 11212
rect 16120 11135 16172 11144
rect 16120 11101 16129 11135
rect 16129 11101 16163 11135
rect 16163 11101 16172 11135
rect 16120 11092 16172 11101
rect 16764 11228 16816 11280
rect 17592 11203 17644 11212
rect 17592 11169 17601 11203
rect 17601 11169 17635 11203
rect 17635 11169 17644 11203
rect 17592 11160 17644 11169
rect 19340 11160 19392 11212
rect 24216 11228 24268 11280
rect 20996 11160 21048 11212
rect 16672 11092 16724 11144
rect 17868 11092 17920 11144
rect 19984 11092 20036 11144
rect 21088 11092 21140 11144
rect 25320 11135 25372 11144
rect 25320 11101 25329 11135
rect 25329 11101 25363 11135
rect 25363 11101 25372 11135
rect 25320 11092 25372 11101
rect 26516 11160 26568 11212
rect 29184 11160 29236 11212
rect 29828 11160 29880 11212
rect 31944 11160 31996 11212
rect 25688 11092 25740 11144
rect 16304 11024 16356 11076
rect 20536 11024 20588 11076
rect 21916 11067 21968 11076
rect 21916 11033 21925 11067
rect 21925 11033 21959 11067
rect 21959 11033 21968 11067
rect 21916 11024 21968 11033
rect 23664 11024 23716 11076
rect 27620 11092 27672 11144
rect 27804 11135 27856 11144
rect 27804 11101 27813 11135
rect 27813 11101 27847 11135
rect 27847 11101 27856 11135
rect 27804 11092 27856 11101
rect 27988 11092 28040 11144
rect 41052 11296 41104 11348
rect 44916 11296 44968 11348
rect 45836 11296 45888 11348
rect 46664 11296 46716 11348
rect 47676 11339 47728 11348
rect 47676 11305 47685 11339
rect 47685 11305 47719 11339
rect 47719 11305 47728 11339
rect 47676 11296 47728 11305
rect 35808 11228 35860 11280
rect 36176 11228 36228 11280
rect 30288 11092 30340 11144
rect 31484 11135 31536 11144
rect 31484 11101 31493 11135
rect 31493 11101 31527 11135
rect 31527 11101 31536 11135
rect 31484 11092 31536 11101
rect 33692 11135 33744 11144
rect 33692 11101 33701 11135
rect 33701 11101 33735 11135
rect 33735 11101 33744 11135
rect 33692 11092 33744 11101
rect 33784 11135 33836 11144
rect 33784 11101 33793 11135
rect 33793 11101 33827 11135
rect 33827 11101 33836 11135
rect 34796 11135 34848 11144
rect 33784 11092 33836 11101
rect 34796 11101 34805 11135
rect 34805 11101 34839 11135
rect 34839 11101 34848 11135
rect 34796 11092 34848 11101
rect 35348 11160 35400 11212
rect 35440 11135 35492 11144
rect 32680 11024 32732 11076
rect 33600 11024 33652 11076
rect 3792 10956 3844 11008
rect 4068 10956 4120 11008
rect 10140 10956 10192 11008
rect 12348 10999 12400 11008
rect 12348 10965 12357 10999
rect 12357 10965 12391 10999
rect 12391 10965 12400 10999
rect 12348 10956 12400 10965
rect 16948 10956 17000 11008
rect 22928 10999 22980 11008
rect 22928 10965 22937 10999
rect 22937 10965 22971 10999
rect 22971 10965 22980 10999
rect 22928 10956 22980 10965
rect 28080 10999 28132 11008
rect 28080 10965 28089 10999
rect 28089 10965 28123 10999
rect 28123 10965 28132 10999
rect 28080 10956 28132 10965
rect 34704 11024 34756 11076
rect 35440 11101 35449 11135
rect 35449 11101 35483 11135
rect 35483 11101 35492 11135
rect 35440 11092 35492 11101
rect 36084 11092 36136 11144
rect 38568 11135 38620 11144
rect 38568 11101 38577 11135
rect 38577 11101 38611 11135
rect 38611 11101 38620 11135
rect 38568 11092 38620 11101
rect 39028 11160 39080 11212
rect 40316 11203 40368 11212
rect 40316 11169 40325 11203
rect 40325 11169 40359 11203
rect 40359 11169 40368 11203
rect 40316 11160 40368 11169
rect 38936 11135 38988 11144
rect 38936 11101 38945 11135
rect 38945 11101 38979 11135
rect 38979 11101 38988 11135
rect 38936 11092 38988 11101
rect 43168 11228 43220 11280
rect 45928 11228 45980 11280
rect 48596 11228 48648 11280
rect 52736 11271 52788 11280
rect 52736 11237 52745 11271
rect 52745 11237 52779 11271
rect 52779 11237 52788 11271
rect 52736 11228 52788 11237
rect 56968 11228 57020 11280
rect 42340 11135 42392 11144
rect 42340 11101 42349 11135
rect 42349 11101 42383 11135
rect 42383 11101 42392 11135
rect 42340 11092 42392 11101
rect 43076 11092 43128 11144
rect 45744 11092 45796 11144
rect 47676 11160 47728 11212
rect 53288 11203 53340 11212
rect 53288 11169 53297 11203
rect 53297 11169 53331 11203
rect 53331 11169 53340 11203
rect 53288 11160 53340 11169
rect 54024 11203 54076 11212
rect 54024 11169 54033 11203
rect 54033 11169 54067 11203
rect 54067 11169 54076 11203
rect 54024 11160 54076 11169
rect 38476 11024 38528 11076
rect 39856 11024 39908 11076
rect 43812 11024 43864 11076
rect 35532 10956 35584 11008
rect 41420 10956 41472 11008
rect 45376 11024 45428 11076
rect 48596 11092 48648 11144
rect 48688 11067 48740 11076
rect 48412 10956 48464 11008
rect 48688 11033 48697 11067
rect 48697 11033 48731 11067
rect 48731 11033 48740 11067
rect 48688 11024 48740 11033
rect 51540 11092 51592 11144
rect 53012 11135 53064 11144
rect 53012 11101 53021 11135
rect 53021 11101 53055 11135
rect 53055 11101 53064 11135
rect 53012 11092 53064 11101
rect 53840 11092 53892 11144
rect 54668 11092 54720 11144
rect 56508 11092 56560 11144
rect 57612 11160 57664 11212
rect 57428 11092 57480 11144
rect 48964 10956 49016 11008
rect 51816 10999 51868 11008
rect 51816 10965 51825 10999
rect 51825 10965 51859 10999
rect 51859 10965 51868 10999
rect 51816 10956 51868 10965
rect 56968 10956 57020 11008
rect 19574 10854 19626 10906
rect 19638 10854 19690 10906
rect 19702 10854 19754 10906
rect 19766 10854 19818 10906
rect 19830 10854 19882 10906
rect 50294 10854 50346 10906
rect 50358 10854 50410 10906
rect 50422 10854 50474 10906
rect 50486 10854 50538 10906
rect 50550 10854 50602 10906
rect 2780 10752 2832 10804
rect 3884 10752 3936 10804
rect 6368 10795 6420 10804
rect 6368 10761 6377 10795
rect 6377 10761 6411 10795
rect 6411 10761 6420 10795
rect 6368 10752 6420 10761
rect 9312 10752 9364 10804
rect 10048 10795 10100 10804
rect 10048 10761 10057 10795
rect 10057 10761 10091 10795
rect 10091 10761 10100 10795
rect 10048 10752 10100 10761
rect 15200 10752 15252 10804
rect 16120 10752 16172 10804
rect 17040 10752 17092 10804
rect 1400 10659 1452 10668
rect 1400 10625 1409 10659
rect 1409 10625 1443 10659
rect 1443 10625 1452 10659
rect 1400 10616 1452 10625
rect 3700 10616 3752 10668
rect 4068 10616 4120 10668
rect 6828 10616 6880 10668
rect 15108 10727 15160 10736
rect 15108 10693 15117 10727
rect 15117 10693 15151 10727
rect 15151 10693 15160 10727
rect 15108 10684 15160 10693
rect 20076 10684 20128 10736
rect 24768 10752 24820 10804
rect 24308 10684 24360 10736
rect 24400 10727 24452 10736
rect 24400 10693 24409 10727
rect 24409 10693 24443 10727
rect 24443 10693 24452 10727
rect 27436 10752 27488 10804
rect 24400 10684 24452 10693
rect 10140 10659 10192 10668
rect 10140 10625 10149 10659
rect 10149 10625 10183 10659
rect 10183 10625 10192 10659
rect 12164 10659 12216 10668
rect 10140 10616 10192 10625
rect 12164 10625 12173 10659
rect 12173 10625 12207 10659
rect 12207 10625 12216 10659
rect 12164 10616 12216 10625
rect 12348 10659 12400 10668
rect 12348 10625 12357 10659
rect 12357 10625 12391 10659
rect 12391 10625 12400 10659
rect 12348 10616 12400 10625
rect 13176 10659 13228 10668
rect 13176 10625 13185 10659
rect 13185 10625 13219 10659
rect 13219 10625 13228 10659
rect 13176 10616 13228 10625
rect 3240 10591 3292 10600
rect 3240 10557 3249 10591
rect 3249 10557 3283 10591
rect 3283 10557 3292 10591
rect 3240 10548 3292 10557
rect 6000 10548 6052 10600
rect 9496 10591 9548 10600
rect 9496 10557 9505 10591
rect 9505 10557 9539 10591
rect 9539 10557 9548 10591
rect 9496 10548 9548 10557
rect 10692 10591 10744 10600
rect 10692 10557 10701 10591
rect 10701 10557 10735 10591
rect 10735 10557 10744 10591
rect 10692 10548 10744 10557
rect 6644 10480 6696 10532
rect 11520 10412 11572 10464
rect 12440 10412 12492 10464
rect 15752 10412 15804 10464
rect 19708 10659 19760 10668
rect 18696 10412 18748 10464
rect 19708 10625 19716 10659
rect 19716 10625 19750 10659
rect 19750 10625 19760 10659
rect 19708 10616 19760 10625
rect 22928 10659 22980 10668
rect 20352 10548 20404 10600
rect 22928 10625 22937 10659
rect 22937 10625 22971 10659
rect 22971 10625 22980 10659
rect 22928 10616 22980 10625
rect 23296 10659 23348 10668
rect 23296 10625 23305 10659
rect 23305 10625 23339 10659
rect 23339 10625 23348 10659
rect 23296 10616 23348 10625
rect 23664 10548 23716 10600
rect 25228 10659 25280 10668
rect 25228 10625 25237 10659
rect 25237 10625 25271 10659
rect 25271 10625 25280 10659
rect 25228 10616 25280 10625
rect 25964 10616 26016 10668
rect 29460 10752 29512 10804
rect 28080 10616 28132 10668
rect 29368 10659 29420 10668
rect 29368 10625 29377 10659
rect 29377 10625 29411 10659
rect 29411 10625 29420 10659
rect 29368 10616 29420 10625
rect 29736 10659 29788 10668
rect 29736 10625 29745 10659
rect 29745 10625 29779 10659
rect 29779 10625 29788 10659
rect 29736 10616 29788 10625
rect 29920 10616 29972 10668
rect 25412 10548 25464 10600
rect 27712 10548 27764 10600
rect 28724 10548 28776 10600
rect 43168 10752 43220 10804
rect 47676 10752 47728 10804
rect 31484 10684 31536 10736
rect 23940 10480 23992 10532
rect 27804 10523 27856 10532
rect 24124 10412 24176 10464
rect 24308 10455 24360 10464
rect 24308 10421 24317 10455
rect 24317 10421 24351 10455
rect 24351 10421 24360 10455
rect 24308 10412 24360 10421
rect 24952 10455 25004 10464
rect 24952 10421 24961 10455
rect 24961 10421 24995 10455
rect 24995 10421 25004 10455
rect 24952 10412 25004 10421
rect 26056 10455 26108 10464
rect 26056 10421 26065 10455
rect 26065 10421 26099 10455
rect 26099 10421 26108 10455
rect 26056 10412 26108 10421
rect 27804 10489 27813 10523
rect 27813 10489 27847 10523
rect 27847 10489 27856 10523
rect 27804 10480 27856 10489
rect 33600 10659 33652 10668
rect 33600 10625 33609 10659
rect 33609 10625 33643 10659
rect 33643 10625 33652 10659
rect 33600 10616 33652 10625
rect 34704 10684 34756 10736
rect 35440 10616 35492 10668
rect 37372 10659 37424 10668
rect 37372 10625 37381 10659
rect 37381 10625 37415 10659
rect 37415 10625 37424 10659
rect 37372 10616 37424 10625
rect 39856 10727 39908 10736
rect 39856 10693 39865 10727
rect 39865 10693 39899 10727
rect 39899 10693 39908 10727
rect 39856 10684 39908 10693
rect 38936 10659 38988 10668
rect 34796 10548 34848 10600
rect 38292 10591 38344 10600
rect 38292 10557 38301 10591
rect 38301 10557 38335 10591
rect 38335 10557 38344 10591
rect 38292 10548 38344 10557
rect 38936 10625 38945 10659
rect 38945 10625 38979 10659
rect 38979 10625 38988 10659
rect 38936 10616 38988 10625
rect 40316 10616 40368 10668
rect 41144 10684 41196 10736
rect 53012 10752 53064 10804
rect 53840 10752 53892 10804
rect 56232 10752 56284 10804
rect 51816 10684 51868 10736
rect 48964 10659 49016 10668
rect 48964 10625 48973 10659
rect 48973 10625 49007 10659
rect 49007 10625 49016 10659
rect 48964 10616 49016 10625
rect 51724 10659 51776 10668
rect 51724 10625 51733 10659
rect 51733 10625 51767 10659
rect 51767 10625 51776 10659
rect 51724 10616 51776 10625
rect 52092 10659 52144 10668
rect 52092 10625 52101 10659
rect 52101 10625 52135 10659
rect 52135 10625 52144 10659
rect 52092 10616 52144 10625
rect 53656 10659 53708 10668
rect 49516 10591 49568 10600
rect 49516 10557 49525 10591
rect 49525 10557 49559 10591
rect 49559 10557 49568 10591
rect 49516 10548 49568 10557
rect 51540 10548 51592 10600
rect 53656 10625 53665 10659
rect 53665 10625 53699 10659
rect 53699 10625 53708 10659
rect 53656 10616 53708 10625
rect 55128 10684 55180 10736
rect 56876 10684 56928 10736
rect 54116 10616 54168 10668
rect 54668 10659 54720 10668
rect 54668 10625 54677 10659
rect 54677 10625 54711 10659
rect 54711 10625 54720 10659
rect 54668 10616 54720 10625
rect 56784 10616 56836 10668
rect 57428 10616 57480 10668
rect 57612 10616 57664 10668
rect 54024 10548 54076 10600
rect 29828 10412 29880 10464
rect 30288 10412 30340 10464
rect 31024 10412 31076 10464
rect 35256 10480 35308 10532
rect 38936 10523 38988 10532
rect 38936 10489 38945 10523
rect 38945 10489 38979 10523
rect 38979 10489 38988 10523
rect 38936 10480 38988 10489
rect 35532 10412 35584 10464
rect 39856 10412 39908 10464
rect 40960 10455 41012 10464
rect 40960 10421 40969 10455
rect 40969 10421 41003 10455
rect 41003 10421 41012 10455
rect 40960 10412 41012 10421
rect 54576 10455 54628 10464
rect 54576 10421 54585 10455
rect 54585 10421 54619 10455
rect 54619 10421 54628 10455
rect 54576 10412 54628 10421
rect 56508 10412 56560 10464
rect 58072 10455 58124 10464
rect 58072 10421 58081 10455
rect 58081 10421 58115 10455
rect 58115 10421 58124 10455
rect 58072 10412 58124 10421
rect 4214 10310 4266 10362
rect 4278 10310 4330 10362
rect 4342 10310 4394 10362
rect 4406 10310 4458 10362
rect 4470 10310 4522 10362
rect 34934 10310 34986 10362
rect 34998 10310 35050 10362
rect 35062 10310 35114 10362
rect 35126 10310 35178 10362
rect 35190 10310 35242 10362
rect 1400 10251 1452 10260
rect 1400 10217 1409 10251
rect 1409 10217 1443 10251
rect 1443 10217 1452 10251
rect 1400 10208 1452 10217
rect 6000 10208 6052 10260
rect 6828 10251 6880 10260
rect 2872 10004 2924 10056
rect 3148 10047 3200 10056
rect 3148 10013 3157 10047
rect 3157 10013 3191 10047
rect 3191 10013 3200 10047
rect 3148 10004 3200 10013
rect 6828 10217 6837 10251
rect 6837 10217 6871 10251
rect 6871 10217 6880 10251
rect 6828 10208 6880 10217
rect 9496 10208 9548 10260
rect 12164 10208 12216 10260
rect 21824 10208 21876 10260
rect 22468 10208 22520 10260
rect 25320 10208 25372 10260
rect 31576 10208 31628 10260
rect 36360 10251 36412 10260
rect 6920 10140 6972 10192
rect 19156 10140 19208 10192
rect 20352 10140 20404 10192
rect 27436 10140 27488 10192
rect 29736 10140 29788 10192
rect 6368 10072 6420 10124
rect 8852 10072 8904 10124
rect 12624 10115 12676 10124
rect 12624 10081 12633 10115
rect 12633 10081 12667 10115
rect 12667 10081 12676 10115
rect 12624 10072 12676 10081
rect 18696 10072 18748 10124
rect 4068 9936 4120 9988
rect 8208 10004 8260 10056
rect 14924 10047 14976 10056
rect 14924 10013 14933 10047
rect 14933 10013 14967 10047
rect 14967 10013 14976 10047
rect 14924 10004 14976 10013
rect 15108 10004 15160 10056
rect 16948 10004 17000 10056
rect 17040 10047 17092 10056
rect 17040 10013 17049 10047
rect 17049 10013 17083 10047
rect 17083 10013 17092 10047
rect 19248 10047 19300 10056
rect 17040 10004 17092 10013
rect 19248 10013 19257 10047
rect 19257 10013 19291 10047
rect 19291 10013 19300 10047
rect 19248 10004 19300 10013
rect 20260 10004 20312 10056
rect 20444 10004 20496 10056
rect 21824 10047 21876 10056
rect 21824 10013 21833 10047
rect 21833 10013 21867 10047
rect 21867 10013 21876 10047
rect 21824 10004 21876 10013
rect 27528 10072 27580 10124
rect 27620 10072 27672 10124
rect 29368 10072 29420 10124
rect 24952 10004 25004 10056
rect 26516 10047 26568 10056
rect 26516 10013 26525 10047
rect 26525 10013 26559 10047
rect 26559 10013 26568 10047
rect 26516 10004 26568 10013
rect 28448 10047 28500 10056
rect 28448 10013 28457 10047
rect 28457 10013 28491 10047
rect 28491 10013 28500 10047
rect 28448 10004 28500 10013
rect 23388 9936 23440 9988
rect 23664 9936 23716 9988
rect 25504 9936 25556 9988
rect 25596 9936 25648 9988
rect 25964 9936 26016 9988
rect 30748 10004 30800 10056
rect 3424 9868 3476 9920
rect 3792 9868 3844 9920
rect 9588 9868 9640 9920
rect 13084 9868 13136 9920
rect 15752 9911 15804 9920
rect 15752 9877 15761 9911
rect 15761 9877 15795 9911
rect 15795 9877 15804 9911
rect 15752 9868 15804 9877
rect 16580 9868 16632 9920
rect 16856 9868 16908 9920
rect 22376 9911 22428 9920
rect 22376 9877 22385 9911
rect 22385 9877 22419 9911
rect 22419 9877 22428 9911
rect 22376 9868 22428 9877
rect 22652 9868 22704 9920
rect 24768 9868 24820 9920
rect 27712 9868 27764 9920
rect 30840 9868 30892 9920
rect 36360 10217 36369 10251
rect 36369 10217 36403 10251
rect 36403 10217 36412 10251
rect 36360 10208 36412 10217
rect 39304 10208 39356 10260
rect 41052 10208 41104 10260
rect 32680 10047 32732 10056
rect 32680 10013 32689 10047
rect 32689 10013 32723 10047
rect 32723 10013 32732 10047
rect 32680 10004 32732 10013
rect 33416 10004 33468 10056
rect 41880 10140 41932 10192
rect 33692 9911 33744 9920
rect 33692 9877 33701 9911
rect 33701 9877 33735 9911
rect 33735 9877 33744 9911
rect 33692 9868 33744 9877
rect 35348 9868 35400 9920
rect 36544 10047 36596 10056
rect 36544 10013 36553 10047
rect 36553 10013 36587 10047
rect 36587 10013 36596 10047
rect 36544 10004 36596 10013
rect 40960 10047 41012 10056
rect 40960 10013 40969 10047
rect 40969 10013 41003 10047
rect 41003 10013 41012 10047
rect 40960 10004 41012 10013
rect 41052 10004 41104 10056
rect 41420 10004 41472 10056
rect 41788 10004 41840 10056
rect 51724 10208 51776 10260
rect 53656 10208 53708 10260
rect 56692 10208 56744 10260
rect 43168 10115 43220 10124
rect 43168 10081 43177 10115
rect 43177 10081 43211 10115
rect 43211 10081 43220 10115
rect 43168 10072 43220 10081
rect 45560 10115 45612 10124
rect 45560 10081 45569 10115
rect 45569 10081 45603 10115
rect 45603 10081 45612 10115
rect 45560 10072 45612 10081
rect 38476 9936 38528 9988
rect 38660 9936 38712 9988
rect 42892 9936 42944 9988
rect 36728 9911 36780 9920
rect 36728 9877 36737 9911
rect 36737 9877 36771 9911
rect 36771 9877 36780 9911
rect 36728 9868 36780 9877
rect 41512 9868 41564 9920
rect 41696 9911 41748 9920
rect 41696 9877 41705 9911
rect 41705 9877 41739 9911
rect 41739 9877 41748 9911
rect 41696 9868 41748 9877
rect 41788 9868 41840 9920
rect 42708 9868 42760 9920
rect 47768 10047 47820 10056
rect 47768 10013 47777 10047
rect 47777 10013 47811 10047
rect 47811 10013 47820 10047
rect 47768 10004 47820 10013
rect 48412 10004 48464 10056
rect 55588 10115 55640 10124
rect 55588 10081 55597 10115
rect 55597 10081 55631 10115
rect 55631 10081 55640 10115
rect 55588 10072 55640 10081
rect 56508 10072 56560 10124
rect 51172 9979 51224 9988
rect 51172 9945 51181 9979
rect 51181 9945 51215 9979
rect 51215 9945 51224 9979
rect 51172 9936 51224 9945
rect 51816 10004 51868 10056
rect 55956 10004 56008 10056
rect 56968 10047 57020 10056
rect 56968 10013 56977 10047
rect 56977 10013 57011 10047
rect 57011 10013 57020 10047
rect 56968 10004 57020 10013
rect 52092 9936 52144 9988
rect 44180 9868 44232 9920
rect 57152 9911 57204 9920
rect 57152 9877 57161 9911
rect 57161 9877 57195 9911
rect 57195 9877 57204 9911
rect 57152 9868 57204 9877
rect 57612 9868 57664 9920
rect 19574 9766 19626 9818
rect 19638 9766 19690 9818
rect 19702 9766 19754 9818
rect 19766 9766 19818 9818
rect 19830 9766 19882 9818
rect 50294 9766 50346 9818
rect 50358 9766 50410 9818
rect 50422 9766 50474 9818
rect 50486 9766 50538 9818
rect 50550 9766 50602 9818
rect 6368 9707 6420 9716
rect 6368 9673 6377 9707
rect 6377 9673 6411 9707
rect 6411 9673 6420 9707
rect 6368 9664 6420 9673
rect 14004 9664 14056 9716
rect 15752 9664 15804 9716
rect 6920 9596 6972 9648
rect 9588 9639 9640 9648
rect 3056 9528 3108 9580
rect 3424 9571 3476 9580
rect 3424 9537 3433 9571
rect 3433 9537 3467 9571
rect 3467 9537 3476 9571
rect 3424 9528 3476 9537
rect 3792 9571 3844 9580
rect 3792 9537 3801 9571
rect 3801 9537 3835 9571
rect 3835 9537 3844 9571
rect 3792 9528 3844 9537
rect 4620 9528 4672 9580
rect 8852 9571 8904 9580
rect 6552 9460 6604 9512
rect 8852 9537 8861 9571
rect 8861 9537 8895 9571
rect 8895 9537 8904 9571
rect 8852 9528 8904 9537
rect 9588 9605 9597 9639
rect 9597 9605 9631 9639
rect 9631 9605 9640 9639
rect 9588 9596 9640 9605
rect 13728 9596 13780 9648
rect 17040 9596 17092 9648
rect 11520 9571 11572 9580
rect 11520 9537 11529 9571
rect 11529 9537 11563 9571
rect 11563 9537 11572 9571
rect 11520 9528 11572 9537
rect 12440 9528 12492 9580
rect 12624 9571 12676 9580
rect 12624 9537 12633 9571
rect 12633 9537 12667 9571
rect 12667 9537 12676 9571
rect 12624 9528 12676 9537
rect 13084 9571 13136 9580
rect 13084 9537 13093 9571
rect 13093 9537 13127 9571
rect 13127 9537 13136 9571
rect 13084 9528 13136 9537
rect 16948 9528 17000 9580
rect 7012 9460 7064 9512
rect 19156 9571 19208 9580
rect 19156 9537 19165 9571
rect 19165 9537 19199 9571
rect 19199 9537 19208 9571
rect 19156 9528 19208 9537
rect 20352 9571 20404 9580
rect 20352 9537 20361 9571
rect 20361 9537 20395 9571
rect 20395 9537 20404 9571
rect 20352 9528 20404 9537
rect 20536 9596 20588 9648
rect 23296 9664 23348 9716
rect 22928 9639 22980 9648
rect 22928 9605 22937 9639
rect 22937 9605 22971 9639
rect 22971 9605 22980 9639
rect 22928 9596 22980 9605
rect 20628 9571 20680 9580
rect 20628 9537 20637 9571
rect 20637 9537 20671 9571
rect 20671 9537 20680 9571
rect 20628 9528 20680 9537
rect 20720 9571 20772 9580
rect 20720 9537 20729 9571
rect 20729 9537 20763 9571
rect 20763 9537 20772 9571
rect 20720 9528 20772 9537
rect 22652 9528 22704 9580
rect 23388 9596 23440 9648
rect 23296 9528 23348 9580
rect 23664 9528 23716 9580
rect 3056 9392 3108 9444
rect 22284 9392 22336 9444
rect 24032 9596 24084 9648
rect 29092 9664 29144 9716
rect 29736 9664 29788 9716
rect 35348 9707 35400 9716
rect 25596 9639 25648 9648
rect 25596 9605 25605 9639
rect 25605 9605 25639 9639
rect 25639 9605 25648 9639
rect 25596 9596 25648 9605
rect 24676 9571 24728 9580
rect 24676 9537 24685 9571
rect 24685 9537 24719 9571
rect 24719 9537 24728 9571
rect 24676 9528 24728 9537
rect 24768 9528 24820 9580
rect 25504 9571 25556 9580
rect 25504 9537 25513 9571
rect 25513 9537 25547 9571
rect 25547 9537 25556 9571
rect 25504 9528 25556 9537
rect 25688 9571 25740 9580
rect 25688 9537 25697 9571
rect 25697 9537 25731 9571
rect 25731 9537 25740 9571
rect 25688 9528 25740 9537
rect 26516 9528 26568 9580
rect 27344 9596 27396 9648
rect 28724 9596 28776 9648
rect 28632 9528 28684 9580
rect 29368 9596 29420 9648
rect 29460 9596 29512 9648
rect 29920 9639 29972 9648
rect 29920 9605 29929 9639
rect 29929 9605 29963 9639
rect 29963 9605 29972 9639
rect 29920 9596 29972 9605
rect 35348 9673 35357 9707
rect 35357 9673 35391 9707
rect 35391 9673 35400 9707
rect 35348 9664 35400 9673
rect 29000 9528 29052 9580
rect 29828 9571 29880 9580
rect 29828 9537 29835 9571
rect 29835 9537 29880 9571
rect 29828 9528 29880 9537
rect 35900 9596 35952 9648
rect 41512 9596 41564 9648
rect 42708 9639 42760 9648
rect 36360 9571 36412 9580
rect 24216 9460 24268 9512
rect 26056 9460 26108 9512
rect 27436 9460 27488 9512
rect 29460 9460 29512 9512
rect 36360 9537 36369 9571
rect 36369 9537 36403 9571
rect 36403 9537 36412 9571
rect 36360 9528 36412 9537
rect 41696 9571 41748 9580
rect 41696 9537 41705 9571
rect 41705 9537 41739 9571
rect 41739 9537 41748 9571
rect 41696 9528 41748 9537
rect 42708 9605 42717 9639
rect 42717 9605 42751 9639
rect 42751 9605 42760 9639
rect 42708 9596 42760 9605
rect 55128 9664 55180 9716
rect 44180 9639 44232 9648
rect 44180 9605 44189 9639
rect 44189 9605 44223 9639
rect 44223 9605 44232 9639
rect 44180 9596 44232 9605
rect 43168 9528 43220 9580
rect 45560 9528 45612 9580
rect 45836 9571 45888 9580
rect 45836 9537 45845 9571
rect 45845 9537 45879 9571
rect 45879 9537 45888 9571
rect 45836 9528 45888 9537
rect 46020 9571 46072 9580
rect 46020 9537 46029 9571
rect 46029 9537 46063 9571
rect 46063 9537 46072 9571
rect 46020 9528 46072 9537
rect 54024 9571 54076 9580
rect 54024 9537 54033 9571
rect 54033 9537 54067 9571
rect 54067 9537 54076 9571
rect 54024 9528 54076 9537
rect 55312 9571 55364 9580
rect 36544 9503 36596 9512
rect 36544 9469 36553 9503
rect 36553 9469 36587 9503
rect 36587 9469 36596 9503
rect 36544 9460 36596 9469
rect 55312 9537 55321 9571
rect 55321 9537 55355 9571
rect 55355 9537 55364 9571
rect 55312 9528 55364 9537
rect 55588 9460 55640 9512
rect 55956 9528 56008 9580
rect 56232 9460 56284 9512
rect 24308 9392 24360 9444
rect 25688 9392 25740 9444
rect 4712 9324 4764 9376
rect 10876 9324 10928 9376
rect 15844 9367 15896 9376
rect 15844 9333 15853 9367
rect 15853 9333 15887 9367
rect 15887 9333 15896 9367
rect 15844 9324 15896 9333
rect 15936 9324 15988 9376
rect 20168 9367 20220 9376
rect 20168 9333 20177 9367
rect 20177 9333 20211 9367
rect 20211 9333 20220 9367
rect 20168 9324 20220 9333
rect 22468 9324 22520 9376
rect 24860 9367 24912 9376
rect 24860 9333 24869 9367
rect 24869 9333 24903 9367
rect 24903 9333 24912 9367
rect 24860 9324 24912 9333
rect 26884 9324 26936 9376
rect 30564 9324 30616 9376
rect 42524 9324 42576 9376
rect 42892 9367 42944 9376
rect 42892 9333 42901 9367
rect 42901 9333 42935 9367
rect 42935 9333 42944 9367
rect 42892 9324 42944 9333
rect 45928 9324 45980 9376
rect 56140 9392 56192 9444
rect 54484 9367 54536 9376
rect 54484 9333 54493 9367
rect 54493 9333 54527 9367
rect 54527 9333 54536 9367
rect 54484 9324 54536 9333
rect 4214 9222 4266 9274
rect 4278 9222 4330 9274
rect 4342 9222 4394 9274
rect 4406 9222 4458 9274
rect 4470 9222 4522 9274
rect 34934 9222 34986 9274
rect 34998 9222 35050 9274
rect 35062 9222 35114 9274
rect 35126 9222 35178 9274
rect 35190 9222 35242 9274
rect 3240 9163 3292 9172
rect 3240 9129 3249 9163
rect 3249 9129 3283 9163
rect 3283 9129 3292 9163
rect 3240 9120 3292 9129
rect 4068 9120 4120 9172
rect 6552 9163 6604 9172
rect 6552 9129 6561 9163
rect 6561 9129 6595 9163
rect 6595 9129 6604 9163
rect 6552 9120 6604 9129
rect 8208 9163 8260 9172
rect 8208 9129 8217 9163
rect 8217 9129 8251 9163
rect 8251 9129 8260 9163
rect 8208 9120 8260 9129
rect 8852 9120 8904 9172
rect 20628 9120 20680 9172
rect 25504 9120 25556 9172
rect 29000 9163 29052 9172
rect 3148 8916 3200 8968
rect 3608 8916 3660 8968
rect 6460 8916 6512 8968
rect 6920 8916 6972 8968
rect 8576 8984 8628 9036
rect 10048 8984 10100 9036
rect 10600 9052 10652 9104
rect 10968 9027 11020 9036
rect 10968 8993 10977 9027
rect 10977 8993 11011 9027
rect 11011 8993 11020 9027
rect 10968 8984 11020 8993
rect 15936 8984 15988 9036
rect 17500 9027 17552 9036
rect 17500 8993 17509 9027
rect 17509 8993 17543 9027
rect 17543 8993 17552 9027
rect 17500 8984 17552 8993
rect 10876 8959 10928 8968
rect 10876 8925 10885 8959
rect 10885 8925 10919 8959
rect 10919 8925 10928 8959
rect 10876 8916 10928 8925
rect 14924 8916 14976 8968
rect 3056 8891 3108 8900
rect 3056 8857 3065 8891
rect 3065 8857 3099 8891
rect 3099 8857 3108 8891
rect 3056 8848 3108 8857
rect 3792 8891 3844 8900
rect 3792 8857 3801 8891
rect 3801 8857 3835 8891
rect 3835 8857 3844 8891
rect 3792 8848 3844 8857
rect 3884 8848 3936 8900
rect 10048 8891 10100 8900
rect 10048 8857 10057 8891
rect 10057 8857 10091 8891
rect 10091 8857 10100 8891
rect 10048 8848 10100 8857
rect 17224 8916 17276 8968
rect 19248 8916 19300 8968
rect 19524 8959 19576 8968
rect 19524 8925 19533 8959
rect 19533 8925 19567 8959
rect 19567 8925 19576 8959
rect 19524 8916 19576 8925
rect 20260 8916 20312 8968
rect 24676 9052 24728 9104
rect 25596 9052 25648 9104
rect 20904 8984 20956 9036
rect 22468 8959 22520 8968
rect 22468 8925 22477 8959
rect 22477 8925 22511 8959
rect 22511 8925 22520 8959
rect 22468 8916 22520 8925
rect 24216 8984 24268 9036
rect 24860 8984 24912 9036
rect 15844 8891 15896 8900
rect 15844 8857 15853 8891
rect 15853 8857 15887 8891
rect 15887 8857 15896 8891
rect 15844 8848 15896 8857
rect 14464 8780 14516 8832
rect 17684 8780 17736 8832
rect 23020 8916 23072 8968
rect 25044 8916 25096 8968
rect 26056 8916 26108 8968
rect 26332 8916 26384 8968
rect 27252 8959 27304 8968
rect 27252 8925 27261 8959
rect 27261 8925 27295 8959
rect 27295 8925 27304 8959
rect 27252 8916 27304 8925
rect 27528 8959 27580 8968
rect 27528 8925 27537 8959
rect 27537 8925 27571 8959
rect 27571 8925 27580 8959
rect 27528 8916 27580 8925
rect 20260 8780 20312 8832
rect 22284 8780 22336 8832
rect 23020 8823 23072 8832
rect 23020 8789 23029 8823
rect 23029 8789 23063 8823
rect 23063 8789 23072 8823
rect 26516 8891 26568 8900
rect 26516 8857 26525 8891
rect 26525 8857 26559 8891
rect 26559 8857 26568 8891
rect 26516 8848 26568 8857
rect 23020 8780 23072 8789
rect 27252 8780 27304 8832
rect 27344 8780 27396 8832
rect 29000 9129 29009 9163
rect 29009 9129 29043 9163
rect 29043 9129 29052 9163
rect 29000 9120 29052 9129
rect 29092 9120 29144 9172
rect 29644 9052 29696 9104
rect 33232 9120 33284 9172
rect 36360 9120 36412 9172
rect 43168 9120 43220 9172
rect 54024 9120 54076 9172
rect 28632 8959 28684 8968
rect 28632 8925 28641 8959
rect 28641 8925 28675 8959
rect 28675 8925 28684 8959
rect 28632 8916 28684 8925
rect 30932 8984 30984 9036
rect 33140 9052 33192 9104
rect 36728 9095 36780 9104
rect 36728 9061 36737 9095
rect 36737 9061 36771 9095
rect 36771 9061 36780 9095
rect 36728 9052 36780 9061
rect 40132 9052 40184 9104
rect 34612 8984 34664 9036
rect 28540 8848 28592 8900
rect 28724 8894 28776 8946
rect 30840 8959 30892 8968
rect 28908 8848 28960 8900
rect 29460 8848 29512 8900
rect 30840 8925 30849 8959
rect 30849 8925 30883 8959
rect 30883 8925 30892 8959
rect 30840 8916 30892 8925
rect 32128 8916 32180 8968
rect 33140 8916 33192 8968
rect 33692 8916 33744 8968
rect 34428 8916 34480 8968
rect 35900 8984 35952 9036
rect 36268 8984 36320 9036
rect 37924 8984 37976 9036
rect 38292 8984 38344 9036
rect 37556 8916 37608 8968
rect 45560 9052 45612 9104
rect 46020 9052 46072 9104
rect 45836 9027 45888 9036
rect 41052 8959 41104 8968
rect 41052 8925 41061 8959
rect 41061 8925 41095 8959
rect 41095 8925 41104 8959
rect 41052 8916 41104 8925
rect 45836 8993 45845 9027
rect 45845 8993 45879 9027
rect 45879 8993 45888 9027
rect 45836 8984 45888 8993
rect 49148 9027 49200 9036
rect 49148 8993 49157 9027
rect 49157 8993 49191 9027
rect 49191 8993 49200 9027
rect 49148 8984 49200 8993
rect 51816 9027 51868 9036
rect 51816 8993 51825 9027
rect 51825 8993 51859 9027
rect 51859 8993 51868 9027
rect 51816 8984 51868 8993
rect 30748 8891 30800 8900
rect 30748 8857 30757 8891
rect 30757 8857 30791 8891
rect 30791 8857 30800 8891
rect 30748 8848 30800 8857
rect 48688 8916 48740 8968
rect 48964 8916 49016 8968
rect 39672 8780 39724 8832
rect 51448 8916 51500 8968
rect 55588 8984 55640 9036
rect 56140 8984 56192 9036
rect 55312 8916 55364 8968
rect 56232 8959 56284 8968
rect 56232 8925 56241 8959
rect 56241 8925 56275 8959
rect 56275 8925 56284 8959
rect 56232 8916 56284 8925
rect 56784 8984 56836 9036
rect 19574 8678 19626 8730
rect 19638 8678 19690 8730
rect 19702 8678 19754 8730
rect 19766 8678 19818 8730
rect 19830 8678 19882 8730
rect 50294 8678 50346 8730
rect 50358 8678 50410 8730
rect 50422 8678 50474 8730
rect 50486 8678 50538 8730
rect 50550 8678 50602 8730
rect 2964 8576 3016 8628
rect 4620 8576 4672 8628
rect 8576 8619 8628 8628
rect 8576 8585 8585 8619
rect 8585 8585 8619 8619
rect 8619 8585 8628 8619
rect 8576 8576 8628 8585
rect 17776 8576 17828 8628
rect 18236 8576 18288 8628
rect 21180 8576 21232 8628
rect 22008 8576 22060 8628
rect 28264 8576 28316 8628
rect 3884 8440 3936 8492
rect 4528 8440 4580 8492
rect 17132 8508 17184 8560
rect 22928 8508 22980 8560
rect 25044 8551 25096 8560
rect 25044 8517 25053 8551
rect 25053 8517 25087 8551
rect 25087 8517 25096 8551
rect 25044 8508 25096 8517
rect 28172 8508 28224 8560
rect 29000 8508 29052 8560
rect 29368 8576 29420 8628
rect 30380 8576 30432 8628
rect 36544 8576 36596 8628
rect 39120 8619 39172 8628
rect 39120 8585 39129 8619
rect 39129 8585 39163 8619
rect 39163 8585 39172 8619
rect 39120 8576 39172 8585
rect 48320 8576 48372 8628
rect 51540 8619 51592 8628
rect 51540 8585 51549 8619
rect 51549 8585 51583 8619
rect 51583 8585 51592 8619
rect 51540 8576 51592 8585
rect 56232 8576 56284 8628
rect 29736 8508 29788 8560
rect 36268 8551 36320 8560
rect 36268 8517 36277 8551
rect 36277 8517 36311 8551
rect 36311 8517 36320 8551
rect 36268 8508 36320 8517
rect 6552 8483 6604 8492
rect 6552 8449 6561 8483
rect 6561 8449 6595 8483
rect 6595 8449 6604 8483
rect 6552 8440 6604 8449
rect 7012 8483 7064 8492
rect 3976 8415 4028 8424
rect 3976 8381 3985 8415
rect 3985 8381 4019 8415
rect 4019 8381 4028 8415
rect 3976 8372 4028 8381
rect 7012 8449 7021 8483
rect 7021 8449 7055 8483
rect 7055 8449 7064 8483
rect 7012 8440 7064 8449
rect 15568 8440 15620 8492
rect 19432 8440 19484 8492
rect 6920 8372 6972 8424
rect 7656 8372 7708 8424
rect 24768 8440 24820 8492
rect 25320 8440 25372 8492
rect 28540 8440 28592 8492
rect 28816 8483 28868 8492
rect 28816 8449 28825 8483
rect 28825 8449 28859 8483
rect 28859 8449 28868 8483
rect 28816 8440 28868 8449
rect 1492 8347 1544 8356
rect 1492 8313 1501 8347
rect 1501 8313 1535 8347
rect 1535 8313 1544 8347
rect 1492 8304 1544 8313
rect 3056 8347 3108 8356
rect 3056 8313 3065 8347
rect 3065 8313 3099 8347
rect 3099 8313 3108 8347
rect 3056 8304 3108 8313
rect 4068 8304 4120 8356
rect 3608 8236 3660 8288
rect 3884 8236 3936 8288
rect 23388 8304 23440 8356
rect 25596 8372 25648 8424
rect 30288 8440 30340 8492
rect 34428 8483 34480 8492
rect 34428 8449 34437 8483
rect 34437 8449 34471 8483
rect 34471 8449 34480 8483
rect 34428 8440 34480 8449
rect 34612 8483 34664 8492
rect 34612 8449 34621 8483
rect 34621 8449 34655 8483
rect 34655 8449 34664 8483
rect 34612 8440 34664 8449
rect 37556 8483 37608 8492
rect 37556 8449 37565 8483
rect 37565 8449 37599 8483
rect 37599 8449 37608 8483
rect 37556 8440 37608 8449
rect 37924 8483 37976 8492
rect 37924 8449 37933 8483
rect 37933 8449 37967 8483
rect 37967 8449 37976 8483
rect 37924 8440 37976 8449
rect 38108 8440 38160 8492
rect 52552 8508 52604 8560
rect 40132 8483 40184 8492
rect 39120 8372 39172 8424
rect 40132 8449 40141 8483
rect 40141 8449 40175 8483
rect 40175 8449 40184 8483
rect 40132 8440 40184 8449
rect 41052 8440 41104 8492
rect 42340 8440 42392 8492
rect 46020 8483 46072 8492
rect 46020 8449 46029 8483
rect 46029 8449 46063 8483
rect 46063 8449 46072 8483
rect 46020 8440 46072 8449
rect 48688 8440 48740 8492
rect 48964 8483 49016 8492
rect 48964 8449 48973 8483
rect 48973 8449 49007 8483
rect 49007 8449 49016 8483
rect 48964 8440 49016 8449
rect 49148 8440 49200 8492
rect 51448 8483 51500 8492
rect 51448 8449 51457 8483
rect 51457 8449 51491 8483
rect 51491 8449 51500 8483
rect 51448 8440 51500 8449
rect 51816 8440 51868 8492
rect 52092 8440 52144 8492
rect 52828 8483 52880 8492
rect 52828 8449 52837 8483
rect 52837 8449 52871 8483
rect 52871 8449 52880 8483
rect 52828 8440 52880 8449
rect 54484 8483 54536 8492
rect 54484 8449 54493 8483
rect 54493 8449 54527 8483
rect 54527 8449 54536 8483
rect 54484 8440 54536 8449
rect 57060 8483 57112 8492
rect 57060 8449 57069 8483
rect 57069 8449 57103 8483
rect 57103 8449 57112 8483
rect 57060 8440 57112 8449
rect 45928 8415 45980 8424
rect 45928 8381 45937 8415
rect 45937 8381 45971 8415
rect 45971 8381 45980 8415
rect 45928 8372 45980 8381
rect 54576 8415 54628 8424
rect 54576 8381 54585 8415
rect 54585 8381 54619 8415
rect 54619 8381 54628 8415
rect 54576 8372 54628 8381
rect 56140 8372 56192 8424
rect 57152 8415 57204 8424
rect 57152 8381 57161 8415
rect 57161 8381 57195 8415
rect 57195 8381 57204 8415
rect 57152 8372 57204 8381
rect 27528 8304 27580 8356
rect 31576 8304 31628 8356
rect 39672 8304 39724 8356
rect 45008 8304 45060 8356
rect 48320 8304 48372 8356
rect 48412 8347 48464 8356
rect 48412 8313 48421 8347
rect 48421 8313 48455 8347
rect 48455 8313 48464 8347
rect 48412 8304 48464 8313
rect 54668 8304 54720 8356
rect 12440 8236 12492 8288
rect 15016 8236 15068 8288
rect 21364 8236 21416 8288
rect 31668 8236 31720 8288
rect 4214 8134 4266 8186
rect 4278 8134 4330 8186
rect 4342 8134 4394 8186
rect 4406 8134 4458 8186
rect 4470 8134 4522 8186
rect 34934 8134 34986 8186
rect 34998 8134 35050 8186
rect 35062 8134 35114 8186
rect 35126 8134 35178 8186
rect 35190 8134 35242 8186
rect 3792 8075 3844 8084
rect 3792 8041 3801 8075
rect 3801 8041 3835 8075
rect 3835 8041 3844 8075
rect 3792 8032 3844 8041
rect 6552 8032 6604 8084
rect 7656 8075 7708 8084
rect 7656 8041 7665 8075
rect 7665 8041 7699 8075
rect 7699 8041 7708 8075
rect 7656 8032 7708 8041
rect 10876 8075 10928 8084
rect 10876 8041 10885 8075
rect 10885 8041 10919 8075
rect 10919 8041 10928 8075
rect 10876 8032 10928 8041
rect 26516 8032 26568 8084
rect 28264 8032 28316 8084
rect 35624 8032 35676 8084
rect 3976 8007 4028 8016
rect 3976 7973 3985 8007
rect 3985 7973 4019 8007
rect 4019 7973 4028 8007
rect 3976 7964 4028 7973
rect 10968 7939 11020 7948
rect 10968 7905 10977 7939
rect 10977 7905 11011 7939
rect 11011 7905 11020 7939
rect 10968 7896 11020 7905
rect 4252 7803 4304 7812
rect 4252 7769 4261 7803
rect 4261 7769 4295 7803
rect 4295 7769 4304 7803
rect 4252 7760 4304 7769
rect 11428 7871 11480 7880
rect 11428 7837 11437 7871
rect 11437 7837 11471 7871
rect 11471 7837 11480 7871
rect 11428 7828 11480 7837
rect 11612 7871 11664 7880
rect 11612 7837 11621 7871
rect 11621 7837 11655 7871
rect 11655 7837 11664 7871
rect 11612 7828 11664 7837
rect 9588 7760 9640 7812
rect 10416 7760 10468 7812
rect 17408 7896 17460 7948
rect 17776 7896 17828 7948
rect 20168 7939 20220 7948
rect 20168 7905 20177 7939
rect 20177 7905 20211 7939
rect 20211 7905 20220 7939
rect 20168 7896 20220 7905
rect 21364 7939 21416 7948
rect 21364 7905 21373 7939
rect 21373 7905 21407 7939
rect 21407 7905 21416 7939
rect 21364 7896 21416 7905
rect 22376 7939 22428 7948
rect 22376 7905 22385 7939
rect 22385 7905 22419 7939
rect 22419 7905 22428 7939
rect 22376 7896 22428 7905
rect 14464 7871 14516 7880
rect 14464 7837 14473 7871
rect 14473 7837 14507 7871
rect 14507 7837 14516 7871
rect 14464 7828 14516 7837
rect 14924 7871 14976 7880
rect 14924 7837 14933 7871
rect 14933 7837 14967 7871
rect 14967 7837 14976 7871
rect 14924 7828 14976 7837
rect 18236 7828 18288 7880
rect 20260 7871 20312 7880
rect 20260 7837 20269 7871
rect 20269 7837 20303 7871
rect 20303 7837 20312 7871
rect 21180 7871 21232 7880
rect 20260 7828 20312 7837
rect 21180 7837 21189 7871
rect 21189 7837 21223 7871
rect 21223 7837 21232 7871
rect 21180 7828 21232 7837
rect 23848 7896 23900 7948
rect 10508 7735 10560 7744
rect 10508 7701 10517 7735
rect 10517 7701 10551 7735
rect 10551 7701 10560 7735
rect 10508 7692 10560 7701
rect 11520 7735 11572 7744
rect 11520 7701 11529 7735
rect 11529 7701 11563 7735
rect 11563 7701 11572 7735
rect 11520 7692 11572 7701
rect 18052 7735 18104 7744
rect 18052 7701 18061 7735
rect 18061 7701 18095 7735
rect 18095 7701 18104 7735
rect 18052 7692 18104 7701
rect 19984 7692 20036 7744
rect 20628 7760 20680 7812
rect 27344 7871 27396 7880
rect 27344 7837 27353 7871
rect 27353 7837 27387 7871
rect 27387 7837 27396 7871
rect 27344 7828 27396 7837
rect 27804 7828 27856 7880
rect 28264 7871 28316 7880
rect 28264 7837 28273 7871
rect 28273 7837 28307 7871
rect 28307 7837 28316 7871
rect 28264 7828 28316 7837
rect 28816 7896 28868 7948
rect 30380 7896 30432 7948
rect 24216 7760 24268 7812
rect 28540 7803 28592 7812
rect 28540 7769 28549 7803
rect 28549 7769 28583 7803
rect 28583 7769 28592 7803
rect 28540 7760 28592 7769
rect 23572 7692 23624 7744
rect 23848 7735 23900 7744
rect 23848 7701 23857 7735
rect 23857 7701 23891 7735
rect 23891 7701 23900 7735
rect 23848 7692 23900 7701
rect 27344 7692 27396 7744
rect 27988 7692 28040 7744
rect 29920 7828 29972 7880
rect 45836 7964 45888 8016
rect 49148 7964 49200 8016
rect 52092 8007 52144 8016
rect 52092 7973 52101 8007
rect 52101 7973 52135 8007
rect 52135 7973 52144 8007
rect 52092 7964 52144 7973
rect 31576 7939 31628 7948
rect 31576 7905 31585 7939
rect 31585 7905 31619 7939
rect 31619 7905 31628 7939
rect 31576 7896 31628 7905
rect 32128 7939 32180 7948
rect 32128 7905 32137 7939
rect 32137 7905 32171 7939
rect 32171 7905 32180 7939
rect 32128 7896 32180 7905
rect 33140 7896 33192 7948
rect 33416 7871 33468 7880
rect 33416 7837 33425 7871
rect 33425 7837 33459 7871
rect 33459 7837 33468 7871
rect 38660 7896 38712 7948
rect 33416 7828 33468 7837
rect 35716 7871 35768 7880
rect 35716 7837 35725 7871
rect 35725 7837 35759 7871
rect 35759 7837 35768 7871
rect 35716 7828 35768 7837
rect 35900 7871 35952 7880
rect 35900 7837 35909 7871
rect 35909 7837 35943 7871
rect 35943 7837 35952 7871
rect 35900 7828 35952 7837
rect 39120 7871 39172 7880
rect 39120 7837 39129 7871
rect 39129 7837 39163 7871
rect 39163 7837 39172 7871
rect 39120 7828 39172 7837
rect 39856 7896 39908 7948
rect 41052 7896 41104 7948
rect 39672 7828 39724 7880
rect 41880 7871 41932 7880
rect 37740 7760 37792 7812
rect 41880 7837 41889 7871
rect 41889 7837 41923 7871
rect 41923 7837 41932 7871
rect 41880 7828 41932 7837
rect 42340 7871 42392 7880
rect 42340 7837 42349 7871
rect 42349 7837 42383 7871
rect 42383 7837 42392 7871
rect 42340 7828 42392 7837
rect 42524 7871 42576 7880
rect 42524 7837 42533 7871
rect 42533 7837 42567 7871
rect 42567 7837 42576 7871
rect 42524 7828 42576 7837
rect 48320 7896 48372 7948
rect 45560 7871 45612 7880
rect 45560 7837 45569 7871
rect 45569 7837 45603 7871
rect 45603 7837 45612 7871
rect 45560 7828 45612 7837
rect 45928 7871 45980 7880
rect 45928 7837 45937 7871
rect 45937 7837 45971 7871
rect 45971 7837 45980 7871
rect 45928 7828 45980 7837
rect 46020 7828 46072 7880
rect 48688 7828 48740 7880
rect 51632 7871 51684 7880
rect 51632 7837 51641 7871
rect 51641 7837 51675 7871
rect 51675 7837 51684 7871
rect 51632 7828 51684 7837
rect 51908 7871 51960 7880
rect 51908 7837 51917 7871
rect 51917 7837 51951 7871
rect 51951 7837 51960 7871
rect 51908 7828 51960 7837
rect 52828 7896 52880 7948
rect 52552 7828 52604 7880
rect 58072 7871 58124 7880
rect 58072 7837 58081 7871
rect 58081 7837 58115 7871
rect 58115 7837 58124 7871
rect 58072 7828 58124 7837
rect 57520 7803 57572 7812
rect 31944 7735 31996 7744
rect 31944 7701 31953 7735
rect 31953 7701 31987 7735
rect 31987 7701 31996 7735
rect 31944 7692 31996 7701
rect 33968 7735 34020 7744
rect 33968 7701 33977 7735
rect 33977 7701 34011 7735
rect 34011 7701 34020 7735
rect 33968 7692 34020 7701
rect 34888 7692 34940 7744
rect 35808 7692 35860 7744
rect 36452 7692 36504 7744
rect 38936 7692 38988 7744
rect 57520 7769 57529 7803
rect 57529 7769 57563 7803
rect 57563 7769 57572 7803
rect 57520 7760 57572 7769
rect 42616 7692 42668 7744
rect 45192 7692 45244 7744
rect 19574 7590 19626 7642
rect 19638 7590 19690 7642
rect 19702 7590 19754 7642
rect 19766 7590 19818 7642
rect 19830 7590 19882 7642
rect 50294 7590 50346 7642
rect 50358 7590 50410 7642
rect 50422 7590 50474 7642
rect 50486 7590 50538 7642
rect 50550 7590 50602 7642
rect 10968 7488 11020 7540
rect 11428 7488 11480 7540
rect 12440 7488 12492 7540
rect 13728 7488 13780 7540
rect 20628 7531 20680 7540
rect 20628 7497 20637 7531
rect 20637 7497 20671 7531
rect 20671 7497 20680 7531
rect 20628 7488 20680 7497
rect 27804 7531 27856 7540
rect 27804 7497 27813 7531
rect 27813 7497 27847 7531
rect 27847 7497 27856 7531
rect 27804 7488 27856 7497
rect 28172 7488 28224 7540
rect 31484 7531 31536 7540
rect 14924 7420 14976 7472
rect 6736 7395 6788 7404
rect 6736 7361 6745 7395
rect 6745 7361 6779 7395
rect 6779 7361 6788 7395
rect 6736 7352 6788 7361
rect 10416 7395 10468 7404
rect 10416 7361 10425 7395
rect 10425 7361 10459 7395
rect 10459 7361 10468 7395
rect 10416 7352 10468 7361
rect 14188 7352 14240 7404
rect 17408 7352 17460 7404
rect 17684 7395 17736 7404
rect 17684 7361 17693 7395
rect 17693 7361 17727 7395
rect 17727 7361 17736 7395
rect 17684 7352 17736 7361
rect 4252 7284 4304 7336
rect 6828 7327 6880 7336
rect 6828 7293 6837 7327
rect 6837 7293 6871 7327
rect 6871 7293 6880 7327
rect 6828 7284 6880 7293
rect 11520 7284 11572 7336
rect 14372 7284 14424 7336
rect 23572 7420 23624 7472
rect 14464 7216 14516 7268
rect 18052 7216 18104 7268
rect 23664 7352 23716 7404
rect 23756 7395 23808 7404
rect 23756 7361 23765 7395
rect 23765 7361 23799 7395
rect 23799 7361 23808 7395
rect 26332 7420 26384 7472
rect 23756 7352 23808 7361
rect 27160 7395 27212 7404
rect 20260 7216 20312 7268
rect 27160 7361 27169 7395
rect 27169 7361 27203 7395
rect 27203 7361 27212 7395
rect 27160 7352 27212 7361
rect 28264 7420 28316 7472
rect 27988 7395 28040 7404
rect 27988 7361 27997 7395
rect 27997 7361 28031 7395
rect 28031 7361 28040 7395
rect 27988 7352 28040 7361
rect 28172 7395 28224 7404
rect 28172 7361 28181 7395
rect 28181 7361 28215 7395
rect 28215 7361 28224 7395
rect 31484 7497 31493 7531
rect 31493 7497 31527 7531
rect 31527 7497 31536 7531
rect 31484 7488 31536 7497
rect 31668 7488 31720 7540
rect 28172 7352 28224 7361
rect 29000 7395 29052 7404
rect 29000 7361 29009 7395
rect 29009 7361 29043 7395
rect 29043 7361 29052 7395
rect 29000 7352 29052 7361
rect 30564 7327 30616 7336
rect 30564 7293 30573 7327
rect 30573 7293 30607 7327
rect 30607 7293 30616 7327
rect 30564 7284 30616 7293
rect 27344 7216 27396 7268
rect 27436 7216 27488 7268
rect 31484 7352 31536 7404
rect 31024 7259 31076 7268
rect 31024 7225 31033 7259
rect 31033 7225 31067 7259
rect 31067 7225 31076 7259
rect 31024 7216 31076 7225
rect 35532 7488 35584 7540
rect 31944 7420 31996 7472
rect 43536 7488 43588 7540
rect 46020 7531 46072 7540
rect 46020 7497 46029 7531
rect 46029 7497 46063 7531
rect 46063 7497 46072 7531
rect 46020 7488 46072 7497
rect 58072 7531 58124 7540
rect 58072 7497 58081 7531
rect 58081 7497 58115 7531
rect 58115 7497 58124 7531
rect 58072 7488 58124 7497
rect 35900 7420 35952 7472
rect 42524 7420 42576 7472
rect 32312 7352 32364 7404
rect 33968 7352 34020 7404
rect 34888 7395 34940 7404
rect 34888 7361 34897 7395
rect 34897 7361 34931 7395
rect 34931 7361 34940 7395
rect 34888 7352 34940 7361
rect 35716 7395 35768 7404
rect 33232 7327 33284 7336
rect 33232 7293 33241 7327
rect 33241 7293 33275 7327
rect 33275 7293 33284 7327
rect 33232 7284 33284 7293
rect 35716 7361 35725 7395
rect 35725 7361 35759 7395
rect 35759 7361 35768 7395
rect 35716 7352 35768 7361
rect 38936 7352 38988 7404
rect 42616 7395 42668 7404
rect 42616 7361 42625 7395
rect 42625 7361 42659 7395
rect 42659 7361 42668 7395
rect 42616 7352 42668 7361
rect 52828 7420 52880 7472
rect 45008 7395 45060 7404
rect 45008 7361 45017 7395
rect 45017 7361 45051 7395
rect 45051 7361 45060 7395
rect 45008 7352 45060 7361
rect 45192 7395 45244 7404
rect 45192 7361 45201 7395
rect 45201 7361 45235 7395
rect 45235 7361 45244 7395
rect 45192 7352 45244 7361
rect 51632 7352 51684 7404
rect 56232 7352 56284 7404
rect 35624 7327 35676 7336
rect 35624 7293 35633 7327
rect 35633 7293 35667 7327
rect 35667 7293 35676 7327
rect 35624 7284 35676 7293
rect 39672 7327 39724 7336
rect 39672 7293 39681 7327
rect 39681 7293 39715 7327
rect 39715 7293 39724 7327
rect 39672 7284 39724 7293
rect 45468 7284 45520 7336
rect 51908 7284 51960 7336
rect 57060 7327 57112 7336
rect 57060 7293 57069 7327
rect 57069 7293 57103 7327
rect 57103 7293 57112 7327
rect 57060 7284 57112 7293
rect 57336 7327 57388 7336
rect 57336 7293 57345 7327
rect 57345 7293 57379 7327
rect 57379 7293 57388 7327
rect 57336 7284 57388 7293
rect 34704 7259 34756 7268
rect 34704 7225 34713 7259
rect 34713 7225 34747 7259
rect 34747 7225 34756 7259
rect 34704 7216 34756 7225
rect 12900 7191 12952 7200
rect 12900 7157 12909 7191
rect 12909 7157 12943 7191
rect 12943 7157 12952 7191
rect 12900 7148 12952 7157
rect 14188 7148 14240 7200
rect 14372 7148 14424 7200
rect 16856 7148 16908 7200
rect 23296 7148 23348 7200
rect 25228 7191 25280 7200
rect 25228 7157 25237 7191
rect 25237 7157 25271 7191
rect 25271 7157 25280 7191
rect 25228 7148 25280 7157
rect 27620 7148 27672 7200
rect 28908 7191 28960 7200
rect 28908 7157 28917 7191
rect 28917 7157 28951 7191
rect 28951 7157 28960 7191
rect 28908 7148 28960 7157
rect 32312 7191 32364 7200
rect 32312 7157 32321 7191
rect 32321 7157 32355 7191
rect 32355 7157 32364 7191
rect 32312 7148 32364 7157
rect 35624 7148 35676 7200
rect 38476 7191 38528 7200
rect 38476 7157 38485 7191
rect 38485 7157 38519 7191
rect 38519 7157 38528 7191
rect 38476 7148 38528 7157
rect 55772 7191 55824 7200
rect 55772 7157 55781 7191
rect 55781 7157 55815 7191
rect 55815 7157 55824 7191
rect 55772 7148 55824 7157
rect 4214 7046 4266 7098
rect 4278 7046 4330 7098
rect 4342 7046 4394 7098
rect 4406 7046 4458 7098
rect 4470 7046 4522 7098
rect 34934 7046 34986 7098
rect 34998 7046 35050 7098
rect 35062 7046 35114 7098
rect 35126 7046 35178 7098
rect 35190 7046 35242 7098
rect 9588 6987 9640 6996
rect 9588 6953 9597 6987
rect 9597 6953 9631 6987
rect 9631 6953 9640 6987
rect 9588 6944 9640 6953
rect 10508 6944 10560 6996
rect 11612 6944 11664 6996
rect 17408 6987 17460 6996
rect 17408 6953 17417 6987
rect 17417 6953 17451 6987
rect 17451 6953 17460 6987
rect 17408 6944 17460 6953
rect 18328 6944 18380 6996
rect 27160 6944 27212 6996
rect 27344 6944 27396 6996
rect 33140 6944 33192 6996
rect 35900 6944 35952 6996
rect 45560 6987 45612 6996
rect 45560 6953 45569 6987
rect 45569 6953 45603 6987
rect 45603 6953 45612 6987
rect 45560 6944 45612 6953
rect 48688 6987 48740 6996
rect 48688 6953 48697 6987
rect 48697 6953 48731 6987
rect 48731 6953 48740 6987
rect 48688 6944 48740 6953
rect 51264 6944 51316 6996
rect 51632 6944 51684 6996
rect 6736 6876 6788 6928
rect 12900 6876 12952 6928
rect 14188 6919 14240 6928
rect 14188 6885 14197 6919
rect 14197 6885 14231 6919
rect 14231 6885 14240 6919
rect 14188 6876 14240 6885
rect 19984 6919 20036 6928
rect 19984 6885 19993 6919
rect 19993 6885 20027 6919
rect 20027 6885 20036 6919
rect 19984 6876 20036 6885
rect 38844 6876 38896 6928
rect 40132 6919 40184 6928
rect 10048 6851 10100 6860
rect 10048 6817 10057 6851
rect 10057 6817 10091 6851
rect 10091 6817 10100 6851
rect 10048 6808 10100 6817
rect 12808 6808 12860 6860
rect 14372 6851 14424 6860
rect 10416 6740 10468 6792
rect 11612 6740 11664 6792
rect 12900 6740 12952 6792
rect 10140 6672 10192 6724
rect 14372 6817 14381 6851
rect 14381 6817 14415 6851
rect 14415 6817 14424 6851
rect 14372 6808 14424 6817
rect 16580 6851 16632 6860
rect 16580 6817 16589 6851
rect 16589 6817 16623 6851
rect 16623 6817 16632 6851
rect 16580 6808 16632 6817
rect 16764 6851 16816 6860
rect 16764 6817 16773 6851
rect 16773 6817 16807 6851
rect 16807 6817 16816 6851
rect 16764 6808 16816 6817
rect 20260 6851 20312 6860
rect 20260 6817 20269 6851
rect 20269 6817 20303 6851
rect 20303 6817 20312 6851
rect 20260 6808 20312 6817
rect 14280 6740 14332 6792
rect 16856 6783 16908 6792
rect 16856 6749 16865 6783
rect 16865 6749 16899 6783
rect 16899 6749 16908 6783
rect 16856 6740 16908 6749
rect 24216 6740 24268 6792
rect 25228 6783 25280 6792
rect 25228 6749 25237 6783
rect 25237 6749 25271 6783
rect 25271 6749 25280 6783
rect 25228 6740 25280 6749
rect 20444 6672 20496 6724
rect 21088 6672 21140 6724
rect 27344 6672 27396 6724
rect 32312 6808 32364 6860
rect 40132 6885 40141 6919
rect 40141 6885 40175 6919
rect 40175 6885 40184 6919
rect 40132 6876 40184 6885
rect 31024 6740 31076 6792
rect 31484 6740 31536 6792
rect 34704 6740 34756 6792
rect 35532 6783 35584 6792
rect 35532 6749 35541 6783
rect 35541 6749 35575 6783
rect 35575 6749 35584 6783
rect 35532 6740 35584 6749
rect 35808 6783 35860 6792
rect 35808 6749 35817 6783
rect 35817 6749 35851 6783
rect 35851 6749 35860 6783
rect 35808 6740 35860 6749
rect 27988 6672 28040 6724
rect 38476 6672 38528 6724
rect 17224 6604 17276 6656
rect 21364 6604 21416 6656
rect 27804 6604 27856 6656
rect 31208 6647 31260 6656
rect 31208 6613 31217 6647
rect 31217 6613 31251 6647
rect 31251 6613 31260 6647
rect 31208 6604 31260 6613
rect 37004 6604 37056 6656
rect 38108 6647 38160 6656
rect 38108 6613 38117 6647
rect 38117 6613 38151 6647
rect 38151 6613 38160 6647
rect 38108 6604 38160 6613
rect 45192 6808 45244 6860
rect 39948 6740 40000 6792
rect 45468 6808 45520 6860
rect 47676 6808 47728 6860
rect 47952 6808 48004 6860
rect 49516 6740 49568 6792
rect 54576 6783 54628 6792
rect 54576 6749 54585 6783
rect 54585 6749 54619 6783
rect 54619 6749 54628 6783
rect 54576 6740 54628 6749
rect 54944 6740 54996 6792
rect 55496 6783 55548 6792
rect 55496 6749 55505 6783
rect 55505 6749 55539 6783
rect 55539 6749 55548 6783
rect 55496 6740 55548 6749
rect 40040 6672 40092 6724
rect 45008 6672 45060 6724
rect 55404 6672 55456 6724
rect 56692 6808 56744 6860
rect 56232 6783 56284 6792
rect 56232 6749 56241 6783
rect 56241 6749 56275 6783
rect 56275 6749 56284 6783
rect 56232 6740 56284 6749
rect 56784 6783 56836 6792
rect 56784 6749 56793 6783
rect 56793 6749 56827 6783
rect 56827 6749 56836 6783
rect 56784 6740 56836 6749
rect 56876 6672 56928 6724
rect 49056 6647 49108 6656
rect 49056 6613 49065 6647
rect 49065 6613 49099 6647
rect 49099 6613 49108 6647
rect 49056 6604 49108 6613
rect 19574 6502 19626 6554
rect 19638 6502 19690 6554
rect 19702 6502 19754 6554
rect 19766 6502 19818 6554
rect 19830 6502 19882 6554
rect 50294 6502 50346 6554
rect 50358 6502 50410 6554
rect 50422 6502 50474 6554
rect 50486 6502 50538 6554
rect 50550 6502 50602 6554
rect 6828 6443 6880 6452
rect 6828 6409 6837 6443
rect 6837 6409 6871 6443
rect 6871 6409 6880 6443
rect 6828 6400 6880 6409
rect 12808 6443 12860 6452
rect 12808 6409 12817 6443
rect 12817 6409 12851 6443
rect 12851 6409 12860 6443
rect 12808 6400 12860 6409
rect 3516 6332 3568 6384
rect 1584 6264 1636 6316
rect 3424 6307 3476 6316
rect 3424 6273 3433 6307
rect 3433 6273 3467 6307
rect 3467 6273 3476 6307
rect 3424 6264 3476 6273
rect 4712 6332 4764 6384
rect 10232 6332 10284 6384
rect 10416 6332 10468 6384
rect 11612 6332 11664 6384
rect 20996 6400 21048 6452
rect 23664 6400 23716 6452
rect 10048 6307 10100 6316
rect 2044 6171 2096 6180
rect 2044 6137 2053 6171
rect 2053 6137 2087 6171
rect 2087 6137 2096 6171
rect 2044 6128 2096 6137
rect 10048 6273 10057 6307
rect 10057 6273 10091 6307
rect 10091 6273 10100 6307
rect 10048 6264 10100 6273
rect 10140 6307 10192 6316
rect 10140 6273 10149 6307
rect 10149 6273 10183 6307
rect 10183 6273 10192 6307
rect 10140 6264 10192 6273
rect 14004 6332 14056 6384
rect 21088 6332 21140 6384
rect 25228 6332 25280 6384
rect 10416 6196 10468 6248
rect 13544 6264 13596 6316
rect 13636 6307 13688 6316
rect 13636 6273 13645 6307
rect 13645 6273 13679 6307
rect 13679 6273 13688 6307
rect 13636 6264 13688 6273
rect 16580 6264 16632 6316
rect 16856 6307 16908 6316
rect 16856 6273 16865 6307
rect 16865 6273 16899 6307
rect 16899 6273 16908 6307
rect 16856 6264 16908 6273
rect 17224 6264 17276 6316
rect 17960 6264 18012 6316
rect 20260 6307 20312 6316
rect 20260 6273 20269 6307
rect 20269 6273 20303 6307
rect 20303 6273 20312 6307
rect 20260 6264 20312 6273
rect 20444 6264 20496 6316
rect 26240 6264 26292 6316
rect 33600 6400 33652 6452
rect 38660 6400 38712 6452
rect 38844 6443 38896 6452
rect 38844 6409 38853 6443
rect 38853 6409 38887 6443
rect 38887 6409 38896 6443
rect 38844 6400 38896 6409
rect 55496 6400 55548 6452
rect 56876 6443 56928 6452
rect 56876 6409 56885 6443
rect 56885 6409 56919 6443
rect 56919 6409 56928 6443
rect 56876 6400 56928 6409
rect 57060 6400 57112 6452
rect 27620 6332 27672 6384
rect 35808 6332 35860 6384
rect 43536 6375 43588 6384
rect 19984 6239 20036 6248
rect 19984 6205 19993 6239
rect 19993 6205 20027 6239
rect 20027 6205 20036 6239
rect 19984 6196 20036 6205
rect 20352 6196 20404 6248
rect 31024 6264 31076 6316
rect 31484 6307 31536 6316
rect 31484 6273 31493 6307
rect 31493 6273 31527 6307
rect 31527 6273 31536 6307
rect 31484 6264 31536 6273
rect 34704 6264 34756 6316
rect 35716 6264 35768 6316
rect 37004 6264 37056 6316
rect 43536 6341 43545 6375
rect 43545 6341 43579 6375
rect 43579 6341 43588 6375
rect 43536 6332 43588 6341
rect 44640 6332 44692 6384
rect 37464 6307 37516 6316
rect 37464 6273 37473 6307
rect 37473 6273 37507 6307
rect 37507 6273 37516 6307
rect 37464 6264 37516 6273
rect 38844 6264 38896 6316
rect 39948 6307 40000 6316
rect 39948 6273 39957 6307
rect 39957 6273 39991 6307
rect 39991 6273 40000 6307
rect 39948 6264 40000 6273
rect 47676 6307 47728 6316
rect 47676 6273 47685 6307
rect 47685 6273 47719 6307
rect 47719 6273 47728 6307
rect 47676 6264 47728 6273
rect 47952 6307 48004 6316
rect 47952 6273 47961 6307
rect 47961 6273 47995 6307
rect 47995 6273 48004 6307
rect 47952 6264 48004 6273
rect 49056 6264 49108 6316
rect 49516 6264 49568 6316
rect 51264 6264 51316 6316
rect 53564 6264 53616 6316
rect 27804 6196 27856 6248
rect 37740 6196 37792 6248
rect 40224 6196 40276 6248
rect 40408 6239 40460 6248
rect 40408 6205 40417 6239
rect 40417 6205 40451 6239
rect 40451 6205 40460 6239
rect 40408 6196 40460 6205
rect 54576 6264 54628 6316
rect 56140 6307 56192 6316
rect 56140 6273 56149 6307
rect 56149 6273 56183 6307
rect 56183 6273 56192 6307
rect 56140 6264 56192 6273
rect 56692 6264 56744 6316
rect 54944 6239 54996 6248
rect 54944 6205 54953 6239
rect 54953 6205 54987 6239
rect 54987 6205 54996 6239
rect 54944 6196 54996 6205
rect 55772 6196 55824 6248
rect 57796 6264 57848 6316
rect 24216 6171 24268 6180
rect 7196 6060 7248 6112
rect 24216 6137 24225 6171
rect 24225 6137 24259 6171
rect 24259 6137 24268 6171
rect 24216 6128 24268 6137
rect 37464 6128 37516 6180
rect 40132 6128 40184 6180
rect 56232 6128 56284 6180
rect 58072 6171 58124 6180
rect 58072 6137 58081 6171
rect 58081 6137 58115 6171
rect 58115 6137 58124 6171
rect 58072 6128 58124 6137
rect 9680 6060 9732 6112
rect 13452 6060 13504 6112
rect 16764 6103 16816 6112
rect 16764 6069 16773 6103
rect 16773 6069 16807 6103
rect 16807 6069 16816 6103
rect 16764 6060 16816 6069
rect 17592 6060 17644 6112
rect 17684 6103 17736 6112
rect 17684 6069 17693 6103
rect 17693 6069 17727 6103
rect 17727 6069 17736 6103
rect 17684 6060 17736 6069
rect 31392 6060 31444 6112
rect 32036 6060 32088 6112
rect 35440 6103 35492 6112
rect 35440 6069 35449 6103
rect 35449 6069 35483 6103
rect 35483 6069 35492 6103
rect 35440 6060 35492 6069
rect 37832 6060 37884 6112
rect 43536 6060 43588 6112
rect 44456 6060 44508 6112
rect 53564 6060 53616 6112
rect 4214 5958 4266 6010
rect 4278 5958 4330 6010
rect 4342 5958 4394 6010
rect 4406 5958 4458 6010
rect 4470 5958 4522 6010
rect 34934 5958 34986 6010
rect 34998 5958 35050 6010
rect 35062 5958 35114 6010
rect 35126 5958 35178 6010
rect 35190 5958 35242 6010
rect 1584 5899 1636 5908
rect 1584 5865 1593 5899
rect 1593 5865 1627 5899
rect 1627 5865 1636 5899
rect 1584 5856 1636 5865
rect 10048 5856 10100 5908
rect 4620 5720 4672 5772
rect 6828 5788 6880 5840
rect 6736 5720 6788 5772
rect 7196 5763 7248 5772
rect 7196 5729 7205 5763
rect 7205 5729 7239 5763
rect 7239 5729 7248 5763
rect 7196 5720 7248 5729
rect 10508 5763 10560 5772
rect 10508 5729 10517 5763
rect 10517 5729 10551 5763
rect 10551 5729 10560 5763
rect 10508 5720 10560 5729
rect 10416 5695 10468 5704
rect 10416 5661 10425 5695
rect 10425 5661 10459 5695
rect 10459 5661 10468 5695
rect 10416 5652 10468 5661
rect 6736 5584 6788 5636
rect 6828 5516 6880 5568
rect 12808 5763 12860 5772
rect 12808 5729 12817 5763
rect 12817 5729 12851 5763
rect 12851 5729 12860 5763
rect 12808 5720 12860 5729
rect 13636 5720 13688 5772
rect 20996 5856 21048 5908
rect 27988 5856 28040 5908
rect 31392 5856 31444 5908
rect 32036 5899 32088 5908
rect 32036 5865 32045 5899
rect 32045 5865 32079 5899
rect 32079 5865 32088 5899
rect 32036 5856 32088 5865
rect 14004 5652 14056 5704
rect 13544 5584 13596 5636
rect 16580 5652 16632 5704
rect 17960 5788 18012 5840
rect 20168 5788 20220 5840
rect 17224 5720 17276 5772
rect 17592 5695 17644 5704
rect 17592 5661 17601 5695
rect 17601 5661 17635 5695
rect 17635 5661 17644 5695
rect 17592 5652 17644 5661
rect 19984 5720 20036 5772
rect 27620 5788 27672 5840
rect 20352 5695 20404 5704
rect 20352 5661 20361 5695
rect 20361 5661 20395 5695
rect 20395 5661 20404 5695
rect 20352 5652 20404 5661
rect 23020 5720 23072 5772
rect 20996 5695 21048 5704
rect 20996 5661 21005 5695
rect 21005 5661 21039 5695
rect 21039 5661 21048 5695
rect 20996 5652 21048 5661
rect 21088 5652 21140 5704
rect 23296 5695 23348 5704
rect 23296 5661 23305 5695
rect 23305 5661 23339 5695
rect 23339 5661 23348 5695
rect 23296 5652 23348 5661
rect 29644 5720 29696 5772
rect 31944 5788 31996 5840
rect 24032 5652 24084 5704
rect 26976 5695 27028 5704
rect 26976 5661 26985 5695
rect 26985 5661 27019 5695
rect 27019 5661 27028 5695
rect 26976 5652 27028 5661
rect 27344 5695 27396 5704
rect 27344 5661 27353 5695
rect 27353 5661 27387 5695
rect 27387 5661 27396 5695
rect 27344 5652 27396 5661
rect 35440 5720 35492 5772
rect 35716 5720 35768 5772
rect 31208 5695 31260 5704
rect 31208 5661 31217 5695
rect 31217 5661 31251 5695
rect 31251 5661 31260 5695
rect 31208 5652 31260 5661
rect 31392 5695 31444 5704
rect 31392 5661 31401 5695
rect 31401 5661 31435 5695
rect 31435 5661 31444 5695
rect 31392 5652 31444 5661
rect 31944 5652 31996 5704
rect 33140 5652 33192 5704
rect 33600 5695 33652 5704
rect 33600 5661 33609 5695
rect 33609 5661 33643 5695
rect 33643 5661 33652 5695
rect 33600 5652 33652 5661
rect 35532 5652 35584 5704
rect 14464 5559 14516 5568
rect 14464 5525 14473 5559
rect 14473 5525 14507 5559
rect 14507 5525 14516 5559
rect 19432 5584 19484 5636
rect 24584 5627 24636 5636
rect 24584 5593 24593 5627
rect 24593 5593 24627 5627
rect 24627 5593 24636 5627
rect 24584 5584 24636 5593
rect 26884 5584 26936 5636
rect 14464 5516 14516 5525
rect 19340 5516 19392 5568
rect 23388 5559 23440 5568
rect 23388 5525 23397 5559
rect 23397 5525 23431 5559
rect 23431 5525 23440 5559
rect 23388 5516 23440 5525
rect 24768 5559 24820 5568
rect 24768 5525 24777 5559
rect 24777 5525 24811 5559
rect 24811 5525 24820 5559
rect 24768 5516 24820 5525
rect 25320 5516 25372 5568
rect 30472 5559 30524 5568
rect 30472 5525 30481 5559
rect 30481 5525 30515 5559
rect 30515 5525 30524 5559
rect 30472 5516 30524 5525
rect 54944 5856 54996 5908
rect 55772 5856 55824 5908
rect 57796 5899 57848 5908
rect 57796 5865 57805 5899
rect 57805 5865 57839 5899
rect 57839 5865 57848 5899
rect 57796 5856 57848 5865
rect 37004 5695 37056 5704
rect 37004 5661 37013 5695
rect 37013 5661 37047 5695
rect 37047 5661 37056 5695
rect 37004 5652 37056 5661
rect 37464 5652 37516 5704
rect 43444 5763 43496 5772
rect 43444 5729 43453 5763
rect 43453 5729 43487 5763
rect 43487 5729 43496 5763
rect 43444 5720 43496 5729
rect 56876 5720 56928 5772
rect 37832 5695 37884 5704
rect 37832 5661 37841 5695
rect 37841 5661 37875 5695
rect 37875 5661 37884 5695
rect 37832 5652 37884 5661
rect 40040 5695 40092 5704
rect 40040 5661 40049 5695
rect 40049 5661 40083 5695
rect 40083 5661 40092 5695
rect 40040 5652 40092 5661
rect 40224 5652 40276 5704
rect 43536 5695 43588 5704
rect 43536 5661 43545 5695
rect 43545 5661 43579 5695
rect 43579 5661 43588 5695
rect 43536 5652 43588 5661
rect 53564 5652 53616 5704
rect 55772 5652 55824 5704
rect 56140 5652 56192 5704
rect 31576 5559 31628 5568
rect 31576 5525 31585 5559
rect 31585 5525 31619 5559
rect 31619 5525 31628 5559
rect 32404 5559 32456 5568
rect 31576 5516 31628 5525
rect 32404 5525 32413 5559
rect 32413 5525 32447 5559
rect 32447 5525 32456 5559
rect 32404 5516 32456 5525
rect 33232 5559 33284 5568
rect 33232 5525 33241 5559
rect 33241 5525 33275 5559
rect 33275 5525 33284 5559
rect 33232 5516 33284 5525
rect 35900 5516 35952 5568
rect 37096 5516 37148 5568
rect 37832 5516 37884 5568
rect 40500 5559 40552 5568
rect 40500 5525 40509 5559
rect 40509 5525 40543 5559
rect 40543 5525 40552 5559
rect 40500 5516 40552 5525
rect 40868 5516 40920 5568
rect 44180 5516 44232 5568
rect 53564 5559 53616 5568
rect 53564 5525 53573 5559
rect 53573 5525 53607 5559
rect 53607 5525 53616 5559
rect 53564 5516 53616 5525
rect 19574 5414 19626 5466
rect 19638 5414 19690 5466
rect 19702 5414 19754 5466
rect 19766 5414 19818 5466
rect 19830 5414 19882 5466
rect 50294 5414 50346 5466
rect 50358 5414 50410 5466
rect 50422 5414 50474 5466
rect 50486 5414 50538 5466
rect 50550 5414 50602 5466
rect 3424 5312 3476 5364
rect 9680 5312 9732 5364
rect 3056 5244 3108 5296
rect 6736 5244 6788 5296
rect 19340 5244 19392 5296
rect 19984 5244 20036 5296
rect 3240 5219 3292 5228
rect 3240 5185 3249 5219
rect 3249 5185 3283 5219
rect 3283 5185 3292 5219
rect 3240 5176 3292 5185
rect 3792 5219 3844 5228
rect 3792 5185 3802 5219
rect 3802 5185 3836 5219
rect 3836 5185 3844 5219
rect 3976 5219 4028 5228
rect 3792 5176 3844 5185
rect 3976 5185 3985 5219
rect 3985 5185 4019 5219
rect 4019 5185 4028 5219
rect 3976 5176 4028 5185
rect 6460 5176 6512 5228
rect 7288 5176 7340 5228
rect 10048 5176 10100 5228
rect 13452 5219 13504 5228
rect 13452 5185 13461 5219
rect 13461 5185 13495 5219
rect 13495 5185 13504 5219
rect 13452 5176 13504 5185
rect 14464 5176 14516 5228
rect 26976 5312 27028 5364
rect 23480 5244 23532 5296
rect 24584 5244 24636 5296
rect 26148 5244 26200 5296
rect 23388 5176 23440 5228
rect 6644 5108 6696 5160
rect 20168 5108 20220 5160
rect 24032 5219 24084 5228
rect 24032 5185 24041 5219
rect 24041 5185 24075 5219
rect 24075 5185 24084 5219
rect 24032 5176 24084 5185
rect 6276 4972 6328 5024
rect 6828 5040 6880 5092
rect 9680 5040 9732 5092
rect 16580 5040 16632 5092
rect 17684 5083 17736 5092
rect 17684 5049 17693 5083
rect 17693 5049 17727 5083
rect 17727 5049 17736 5083
rect 17684 5040 17736 5049
rect 25320 5151 25372 5160
rect 25320 5117 25329 5151
rect 25329 5117 25363 5151
rect 25363 5117 25372 5151
rect 25320 5108 25372 5117
rect 27436 5176 27488 5228
rect 31576 5244 31628 5296
rect 33140 5244 33192 5296
rect 56692 5312 56744 5364
rect 57704 5244 57756 5296
rect 30472 5176 30524 5228
rect 27620 5151 27672 5160
rect 27620 5117 27629 5151
rect 27629 5117 27663 5151
rect 27663 5117 27672 5151
rect 27620 5108 27672 5117
rect 32404 5176 32456 5228
rect 33232 5176 33284 5228
rect 35900 5176 35952 5228
rect 40500 5176 40552 5228
rect 40868 5219 40920 5228
rect 32220 5108 32272 5160
rect 32864 5151 32916 5160
rect 32864 5117 32873 5151
rect 32873 5117 32907 5151
rect 32907 5117 32916 5151
rect 32864 5108 32916 5117
rect 40868 5185 40877 5219
rect 40877 5185 40911 5219
rect 40911 5185 40920 5219
rect 40868 5176 40920 5185
rect 44180 5219 44232 5228
rect 44180 5185 44189 5219
rect 44189 5185 44223 5219
rect 44223 5185 44232 5219
rect 44180 5176 44232 5185
rect 44272 5219 44324 5228
rect 44272 5185 44281 5219
rect 44281 5185 44315 5219
rect 44315 5185 44324 5219
rect 44456 5219 44508 5228
rect 44272 5176 44324 5185
rect 44456 5185 44465 5219
rect 44465 5185 44499 5219
rect 44499 5185 44508 5219
rect 44456 5176 44508 5185
rect 45192 5219 45244 5228
rect 45192 5185 45201 5219
rect 45201 5185 45235 5219
rect 45235 5185 45244 5219
rect 45192 5176 45244 5185
rect 56876 5176 56928 5228
rect 41236 5108 41288 5160
rect 38660 5040 38712 5092
rect 40500 5040 40552 5092
rect 44364 5151 44416 5160
rect 44364 5117 44373 5151
rect 44373 5117 44407 5151
rect 44407 5117 44416 5151
rect 44364 5108 44416 5117
rect 56692 5108 56744 5160
rect 45560 5083 45612 5092
rect 45560 5049 45569 5083
rect 45569 5049 45603 5083
rect 45603 5049 45612 5083
rect 45560 5040 45612 5049
rect 10324 4972 10376 5024
rect 16672 5015 16724 5024
rect 16672 4981 16681 5015
rect 16681 4981 16715 5015
rect 16715 4981 16724 5015
rect 16672 4972 16724 4981
rect 17592 5015 17644 5024
rect 17592 4981 17601 5015
rect 17601 4981 17635 5015
rect 17635 4981 17644 5015
rect 17592 4972 17644 4981
rect 19432 4972 19484 5024
rect 19892 5015 19944 5024
rect 19892 4981 19901 5015
rect 19901 4981 19935 5015
rect 19935 4981 19944 5015
rect 19892 4972 19944 4981
rect 20076 5015 20128 5024
rect 20076 4981 20085 5015
rect 20085 4981 20119 5015
rect 20119 4981 20128 5015
rect 20076 4972 20128 4981
rect 23756 5015 23808 5024
rect 23756 4981 23765 5015
rect 23765 4981 23799 5015
rect 23799 4981 23808 5015
rect 23756 4972 23808 4981
rect 31576 5015 31628 5024
rect 31576 4981 31585 5015
rect 31585 4981 31619 5015
rect 31619 4981 31628 5015
rect 31576 4972 31628 4981
rect 41512 4972 41564 5024
rect 43812 4972 43864 5024
rect 54576 5015 54628 5024
rect 54576 4981 54585 5015
rect 54585 4981 54619 5015
rect 54619 4981 54628 5015
rect 54576 4972 54628 4981
rect 55772 4972 55824 5024
rect 57888 4972 57940 5024
rect 4214 4870 4266 4922
rect 4278 4870 4330 4922
rect 4342 4870 4394 4922
rect 4406 4870 4458 4922
rect 4470 4870 4522 4922
rect 34934 4870 34986 4922
rect 34998 4870 35050 4922
rect 35062 4870 35114 4922
rect 35126 4870 35178 4922
rect 35190 4870 35242 4922
rect 3976 4811 4028 4820
rect 3976 4777 3985 4811
rect 3985 4777 4019 4811
rect 4019 4777 4028 4811
rect 3976 4768 4028 4777
rect 6644 4811 6696 4820
rect 6644 4777 6653 4811
rect 6653 4777 6687 4811
rect 6687 4777 6696 4811
rect 6644 4768 6696 4777
rect 7104 4768 7156 4820
rect 7288 4811 7340 4820
rect 7288 4777 7297 4811
rect 7297 4777 7331 4811
rect 7331 4777 7340 4811
rect 7288 4768 7340 4777
rect 3240 4700 3292 4752
rect 3884 4564 3936 4616
rect 6276 4675 6328 4684
rect 6276 4641 6285 4675
rect 6285 4641 6319 4675
rect 6319 4641 6328 4675
rect 6276 4632 6328 4641
rect 7380 4632 7432 4684
rect 15844 4768 15896 4820
rect 16028 4768 16080 4820
rect 17960 4768 18012 4820
rect 19892 4768 19944 4820
rect 33140 4768 33192 4820
rect 37648 4768 37700 4820
rect 38108 4768 38160 4820
rect 44364 4768 44416 4820
rect 45192 4768 45244 4820
rect 6460 4607 6512 4616
rect 6460 4573 6469 4607
rect 6469 4573 6503 4607
rect 6503 4573 6512 4607
rect 6460 4564 6512 4573
rect 6736 4564 6788 4616
rect 7288 4564 7340 4616
rect 53564 4700 53616 4752
rect 10232 4675 10284 4684
rect 10232 4641 10241 4675
rect 10241 4641 10275 4675
rect 10275 4641 10284 4675
rect 10232 4632 10284 4641
rect 10324 4607 10376 4616
rect 10324 4573 10333 4607
rect 10333 4573 10367 4607
rect 10367 4573 10376 4607
rect 10324 4564 10376 4573
rect 11060 4607 11112 4616
rect 11060 4573 11069 4607
rect 11069 4573 11103 4607
rect 11103 4573 11112 4607
rect 11060 4564 11112 4573
rect 1492 4471 1544 4480
rect 1492 4437 1501 4471
rect 1501 4437 1535 4471
rect 1535 4437 1544 4471
rect 1492 4428 1544 4437
rect 17592 4564 17644 4616
rect 20076 4564 20128 4616
rect 23388 4632 23440 4684
rect 26700 4632 26752 4684
rect 26976 4632 27028 4684
rect 27436 4632 27488 4684
rect 37280 4632 37332 4684
rect 44272 4632 44324 4684
rect 24768 4564 24820 4616
rect 16672 4496 16724 4548
rect 20168 4496 20220 4548
rect 11152 4471 11204 4480
rect 11152 4437 11161 4471
rect 11161 4437 11195 4471
rect 11195 4437 11204 4471
rect 11152 4428 11204 4437
rect 12716 4428 12768 4480
rect 16948 4428 17000 4480
rect 26884 4496 26936 4548
rect 31576 4564 31628 4616
rect 37556 4564 37608 4616
rect 37648 4607 37700 4616
rect 37648 4573 37657 4607
rect 37657 4573 37691 4607
rect 37691 4573 37700 4607
rect 37648 4564 37700 4573
rect 37832 4607 37884 4616
rect 37832 4573 37841 4607
rect 37841 4573 37875 4607
rect 37875 4573 37884 4607
rect 40408 4607 40460 4616
rect 37832 4564 37884 4573
rect 40408 4573 40417 4607
rect 40417 4573 40451 4607
rect 40451 4573 40460 4607
rect 40408 4564 40460 4573
rect 40684 4564 40736 4616
rect 32864 4496 32916 4548
rect 33140 4428 33192 4480
rect 37096 4539 37148 4548
rect 37096 4505 37105 4539
rect 37105 4505 37139 4539
rect 37139 4505 37148 4539
rect 37096 4496 37148 4505
rect 41328 4564 41380 4616
rect 41512 4607 41564 4616
rect 41512 4573 41521 4607
rect 41521 4573 41555 4607
rect 41555 4573 41564 4607
rect 46296 4632 46348 4684
rect 46388 4632 46440 4684
rect 41512 4564 41564 4573
rect 44364 4496 44416 4548
rect 45560 4564 45612 4616
rect 46204 4496 46256 4548
rect 40868 4428 40920 4480
rect 19574 4326 19626 4378
rect 19638 4326 19690 4378
rect 19702 4326 19754 4378
rect 19766 4326 19818 4378
rect 19830 4326 19882 4378
rect 50294 4326 50346 4378
rect 50358 4326 50410 4378
rect 50422 4326 50474 4378
rect 50486 4326 50538 4378
rect 50550 4326 50602 4378
rect 6460 4224 6512 4276
rect 6276 4156 6328 4208
rect 16028 4224 16080 4276
rect 16212 4224 16264 4276
rect 20536 4224 20588 4276
rect 6736 4199 6788 4208
rect 6736 4165 6745 4199
rect 6745 4165 6779 4199
rect 6779 4165 6788 4199
rect 6736 4156 6788 4165
rect 11152 4156 11204 4208
rect 12716 4156 12768 4208
rect 15752 4156 15804 4208
rect 15844 4156 15896 4208
rect 9680 4131 9732 4140
rect 9680 4097 9689 4131
rect 9689 4097 9723 4131
rect 9723 4097 9732 4131
rect 9680 4088 9732 4097
rect 11796 4088 11848 4140
rect 9772 4063 9824 4072
rect 9772 4029 9781 4063
rect 9781 4029 9815 4063
rect 9815 4029 9824 4063
rect 9772 4020 9824 4029
rect 10324 4020 10376 4072
rect 11336 4020 11388 4072
rect 11888 4020 11940 4072
rect 11980 4020 12032 4072
rect 11060 3952 11112 4004
rect 12900 4063 12952 4072
rect 12900 4029 12909 4063
rect 12909 4029 12943 4063
rect 12943 4029 12952 4063
rect 12900 4020 12952 4029
rect 16672 4131 16724 4140
rect 16672 4097 16681 4131
rect 16681 4097 16715 4131
rect 16715 4097 16724 4131
rect 16672 4088 16724 4097
rect 23756 4156 23808 4208
rect 17684 4020 17736 4072
rect 11796 3927 11848 3936
rect 11796 3893 11805 3927
rect 11805 3893 11839 3927
rect 11839 3893 11848 3927
rect 11796 3884 11848 3893
rect 12440 3884 12492 3936
rect 16672 3952 16724 4004
rect 20260 4088 20312 4140
rect 20628 4088 20680 4140
rect 24768 4088 24820 4140
rect 33140 4088 33192 4140
rect 33600 4088 33652 4140
rect 33692 4131 33744 4140
rect 33692 4097 33701 4131
rect 33701 4097 33735 4131
rect 33735 4097 33744 4131
rect 33692 4088 33744 4097
rect 35808 4088 35860 4140
rect 36452 4131 36504 4140
rect 36452 4097 36461 4131
rect 36461 4097 36495 4131
rect 36495 4097 36504 4131
rect 36452 4088 36504 4097
rect 40868 4156 40920 4208
rect 42248 4156 42300 4208
rect 46296 4199 46348 4208
rect 46296 4165 46305 4199
rect 46305 4165 46339 4199
rect 46339 4165 46348 4199
rect 46296 4156 46348 4165
rect 21640 4020 21692 4072
rect 22192 4020 22244 4072
rect 23388 3952 23440 4004
rect 13452 3927 13504 3936
rect 13452 3893 13461 3927
rect 13461 3893 13495 3927
rect 13495 3893 13504 3927
rect 13452 3884 13504 3893
rect 14924 3884 14976 3936
rect 16948 3884 17000 3936
rect 25872 3952 25924 4004
rect 26424 4020 26476 4072
rect 27528 3952 27580 4004
rect 29276 3952 29328 4004
rect 37372 4020 37424 4072
rect 37556 4063 37608 4072
rect 37556 4029 37565 4063
rect 37565 4029 37599 4063
rect 37599 4029 37608 4063
rect 37556 4020 37608 4029
rect 40500 4131 40552 4140
rect 40500 4097 40509 4131
rect 40509 4097 40543 4131
rect 40543 4097 40552 4131
rect 41328 4131 41380 4140
rect 40500 4088 40552 4097
rect 41328 4097 41337 4131
rect 41337 4097 41371 4131
rect 41371 4097 41380 4131
rect 41328 4088 41380 4097
rect 41512 4131 41564 4140
rect 41512 4097 41521 4131
rect 41521 4097 41555 4131
rect 41555 4097 41564 4131
rect 41512 4088 41564 4097
rect 37832 4020 37884 4072
rect 40684 4063 40736 4072
rect 40684 4029 40693 4063
rect 40693 4029 40727 4063
rect 40727 4029 40736 4063
rect 40684 4020 40736 4029
rect 46204 4131 46256 4140
rect 46204 4097 46213 4131
rect 46213 4097 46247 4131
rect 46247 4097 46256 4131
rect 46204 4088 46256 4097
rect 46388 4020 46440 4072
rect 23572 3884 23624 3936
rect 33232 3884 33284 3936
rect 42064 3952 42116 4004
rect 36544 3884 36596 3936
rect 37464 3884 37516 3936
rect 41052 3884 41104 3936
rect 41420 3884 41472 3936
rect 46112 3952 46164 4004
rect 45192 3884 45244 3936
rect 58072 3927 58124 3936
rect 58072 3893 58081 3927
rect 58081 3893 58115 3927
rect 58115 3893 58124 3927
rect 58072 3884 58124 3893
rect 4214 3782 4266 3834
rect 4278 3782 4330 3834
rect 4342 3782 4394 3834
rect 4406 3782 4458 3834
rect 4470 3782 4522 3834
rect 34934 3782 34986 3834
rect 34998 3782 35050 3834
rect 35062 3782 35114 3834
rect 35126 3782 35178 3834
rect 35190 3782 35242 3834
rect 9772 3680 9824 3732
rect 10048 3680 10100 3732
rect 12440 3680 12492 3732
rect 12900 3680 12952 3732
rect 14924 3680 14976 3732
rect 26148 3680 26200 3732
rect 2044 3544 2096 3596
rect 14280 3612 14332 3664
rect 15016 3612 15068 3664
rect 20904 3612 20956 3664
rect 11888 3544 11940 3596
rect 10600 3519 10652 3528
rect 10600 3485 10609 3519
rect 10609 3485 10643 3519
rect 10643 3485 10652 3519
rect 10600 3476 10652 3485
rect 11336 3476 11388 3528
rect 11428 3519 11480 3528
rect 11428 3485 11437 3519
rect 11437 3485 11471 3519
rect 11471 3485 11480 3519
rect 11428 3476 11480 3485
rect 10048 3451 10100 3460
rect 1400 3383 1452 3392
rect 1400 3349 1409 3383
rect 1409 3349 1443 3383
rect 1443 3349 1452 3383
rect 1400 3340 1452 3349
rect 10048 3417 10057 3451
rect 10057 3417 10091 3451
rect 10091 3417 10100 3451
rect 10048 3408 10100 3417
rect 11060 3340 11112 3392
rect 11980 3408 12032 3460
rect 13452 3476 13504 3528
rect 14924 3519 14976 3528
rect 14924 3485 14933 3519
rect 14933 3485 14967 3519
rect 14967 3485 14976 3519
rect 14924 3476 14976 3485
rect 15108 3519 15160 3528
rect 15108 3485 15117 3519
rect 15117 3485 15151 3519
rect 15151 3485 15160 3519
rect 15108 3476 15160 3485
rect 16672 3519 16724 3528
rect 16672 3485 16681 3519
rect 16681 3485 16715 3519
rect 16715 3485 16724 3519
rect 16672 3476 16724 3485
rect 18052 3544 18104 3596
rect 17316 3519 17368 3528
rect 17316 3485 17325 3519
rect 17325 3485 17359 3519
rect 17359 3485 17368 3519
rect 17316 3476 17368 3485
rect 17408 3519 17460 3528
rect 17408 3485 17418 3519
rect 17418 3485 17452 3519
rect 17452 3485 17460 3519
rect 17684 3519 17736 3528
rect 17408 3476 17460 3485
rect 17684 3485 17693 3519
rect 17693 3485 17727 3519
rect 17727 3485 17736 3519
rect 17684 3476 17736 3485
rect 19248 3519 19300 3528
rect 19248 3485 19257 3519
rect 19257 3485 19291 3519
rect 19291 3485 19300 3519
rect 19248 3476 19300 3485
rect 11520 3340 11572 3392
rect 14096 3383 14148 3392
rect 14096 3349 14105 3383
rect 14105 3349 14139 3383
rect 14139 3349 14148 3383
rect 14096 3340 14148 3349
rect 14280 3340 14332 3392
rect 19432 3519 19484 3528
rect 19432 3485 19441 3519
rect 19441 3485 19475 3519
rect 19475 3485 19484 3519
rect 19432 3476 19484 3485
rect 20260 3519 20312 3528
rect 20260 3485 20269 3519
rect 20269 3485 20303 3519
rect 20303 3485 20312 3519
rect 20260 3476 20312 3485
rect 17960 3383 18012 3392
rect 17960 3349 17969 3383
rect 17969 3349 18003 3383
rect 18003 3349 18012 3383
rect 17960 3340 18012 3349
rect 19340 3340 19392 3392
rect 20628 3340 20680 3392
rect 23940 3544 23992 3596
rect 21088 3476 21140 3528
rect 21640 3519 21692 3528
rect 21640 3485 21649 3519
rect 21649 3485 21683 3519
rect 21683 3485 21692 3519
rect 21640 3476 21692 3485
rect 23756 3476 23808 3528
rect 24768 3587 24820 3596
rect 24768 3553 24777 3587
rect 24777 3553 24811 3587
rect 24811 3553 24820 3587
rect 24768 3544 24820 3553
rect 28540 3544 28592 3596
rect 28908 3587 28960 3596
rect 28908 3553 28917 3587
rect 28917 3553 28951 3587
rect 28951 3553 28960 3587
rect 28908 3544 28960 3553
rect 26424 3519 26476 3528
rect 26424 3485 26433 3519
rect 26433 3485 26467 3519
rect 26467 3485 26476 3519
rect 26424 3476 26476 3485
rect 33692 3612 33744 3664
rect 36544 3680 36596 3732
rect 33048 3544 33100 3596
rect 36360 3544 36412 3596
rect 32220 3519 32272 3528
rect 32220 3485 32229 3519
rect 32229 3485 32263 3519
rect 32263 3485 32272 3519
rect 32220 3476 32272 3485
rect 33600 3476 33652 3528
rect 33876 3519 33928 3528
rect 33876 3485 33885 3519
rect 33885 3485 33919 3519
rect 33919 3485 33928 3519
rect 33876 3476 33928 3485
rect 37096 3519 37148 3528
rect 37096 3485 37105 3519
rect 37105 3485 37139 3519
rect 37139 3485 37148 3519
rect 37096 3476 37148 3485
rect 37280 3519 37332 3528
rect 37280 3485 37289 3519
rect 37289 3485 37323 3519
rect 37323 3485 37332 3519
rect 37280 3476 37332 3485
rect 37464 3519 37516 3528
rect 37464 3485 37473 3519
rect 37473 3485 37507 3519
rect 37507 3485 37516 3519
rect 37464 3476 37516 3485
rect 23756 3340 23808 3392
rect 24216 3340 24268 3392
rect 24400 3383 24452 3392
rect 24400 3349 24409 3383
rect 24409 3349 24443 3383
rect 24443 3349 24452 3383
rect 24400 3340 24452 3349
rect 25964 3383 26016 3392
rect 25964 3349 25973 3383
rect 25973 3349 26007 3383
rect 26007 3349 26016 3383
rect 25964 3340 26016 3349
rect 26332 3383 26384 3392
rect 26332 3349 26341 3383
rect 26341 3349 26375 3383
rect 26375 3349 26384 3383
rect 26332 3340 26384 3349
rect 26976 3383 27028 3392
rect 26976 3349 26985 3383
rect 26985 3349 27019 3383
rect 27019 3349 27028 3383
rect 26976 3340 27028 3349
rect 27712 3383 27764 3392
rect 27712 3349 27721 3383
rect 27721 3349 27755 3383
rect 27755 3349 27764 3383
rect 27712 3340 27764 3349
rect 28356 3340 28408 3392
rect 28540 3340 28592 3392
rect 34244 3408 34296 3460
rect 37372 3451 37424 3460
rect 37372 3417 37381 3451
rect 37381 3417 37415 3451
rect 37415 3417 37424 3451
rect 37740 3612 37792 3664
rect 41604 3655 41656 3664
rect 41604 3621 41613 3655
rect 41613 3621 41647 3655
rect 41647 3621 41656 3655
rect 41604 3612 41656 3621
rect 42064 3655 42116 3664
rect 42064 3621 42073 3655
rect 42073 3621 42107 3655
rect 42107 3621 42116 3655
rect 42064 3612 42116 3621
rect 40040 3519 40092 3528
rect 40040 3485 40049 3519
rect 40049 3485 40083 3519
rect 40083 3485 40092 3519
rect 40040 3476 40092 3485
rect 40868 3519 40920 3528
rect 40868 3485 40877 3519
rect 40877 3485 40911 3519
rect 40911 3485 40920 3519
rect 40868 3476 40920 3485
rect 41052 3519 41104 3528
rect 41052 3485 41061 3519
rect 41061 3485 41095 3519
rect 41095 3485 41104 3519
rect 41052 3476 41104 3485
rect 43076 3476 43128 3528
rect 43260 3476 43312 3528
rect 37372 3408 37424 3417
rect 42248 3451 42300 3460
rect 42248 3417 42257 3451
rect 42257 3417 42291 3451
rect 42291 3417 42300 3451
rect 42248 3408 42300 3417
rect 42432 3451 42484 3460
rect 42432 3417 42441 3451
rect 42441 3417 42475 3451
rect 42475 3417 42484 3451
rect 42432 3408 42484 3417
rect 42616 3408 42668 3460
rect 46296 3544 46348 3596
rect 46112 3519 46164 3528
rect 46112 3485 46121 3519
rect 46121 3485 46155 3519
rect 46155 3485 46164 3519
rect 46112 3476 46164 3485
rect 58072 3519 58124 3528
rect 58072 3485 58081 3519
rect 58081 3485 58115 3519
rect 58115 3485 58124 3519
rect 58072 3476 58124 3485
rect 37740 3340 37792 3392
rect 40224 3383 40276 3392
rect 40224 3349 40233 3383
rect 40233 3349 40267 3383
rect 40267 3349 40276 3383
rect 40224 3340 40276 3349
rect 40868 3340 40920 3392
rect 41328 3340 41380 3392
rect 43168 3340 43220 3392
rect 43352 3383 43404 3392
rect 43352 3349 43361 3383
rect 43361 3349 43395 3383
rect 43395 3349 43404 3383
rect 43352 3340 43404 3349
rect 57612 3408 57664 3460
rect 57152 3383 57204 3392
rect 57152 3349 57161 3383
rect 57161 3349 57195 3383
rect 57195 3349 57204 3383
rect 57152 3340 57204 3349
rect 19574 3238 19626 3290
rect 19638 3238 19690 3290
rect 19702 3238 19754 3290
rect 19766 3238 19818 3290
rect 19830 3238 19882 3290
rect 50294 3238 50346 3290
rect 50358 3238 50410 3290
rect 50422 3238 50474 3290
rect 50486 3238 50538 3290
rect 50550 3238 50602 3290
rect 4988 3136 5040 3188
rect 10140 3136 10192 3188
rect 11336 3136 11388 3188
rect 11520 3179 11572 3188
rect 11520 3145 11529 3179
rect 11529 3145 11563 3179
rect 11563 3145 11572 3179
rect 11520 3136 11572 3145
rect 15108 3136 15160 3188
rect 19248 3179 19300 3188
rect 19248 3145 19257 3179
rect 19257 3145 19291 3179
rect 19291 3145 19300 3179
rect 19248 3136 19300 3145
rect 19340 3136 19392 3188
rect 23388 3179 23440 3188
rect 1400 3043 1452 3052
rect 1400 3009 1409 3043
rect 1409 3009 1443 3043
rect 1443 3009 1452 3043
rect 1400 3000 1452 3009
rect 14096 3111 14148 3120
rect 10140 3043 10192 3052
rect 10140 3009 10149 3043
rect 10149 3009 10183 3043
rect 10183 3009 10192 3043
rect 10140 3000 10192 3009
rect 10324 3043 10376 3052
rect 10324 3009 10333 3043
rect 10333 3009 10367 3043
rect 10367 3009 10376 3043
rect 10324 3000 10376 3009
rect 5080 2907 5132 2916
rect 5080 2873 5089 2907
rect 5089 2873 5123 2907
rect 5123 2873 5132 2907
rect 5080 2864 5132 2873
rect 10600 2932 10652 2984
rect 14096 3077 14105 3111
rect 14105 3077 14139 3111
rect 14139 3077 14148 3111
rect 14096 3068 14148 3077
rect 15016 3068 15068 3120
rect 11980 3043 12032 3052
rect 11980 3009 11989 3043
rect 11989 3009 12023 3043
rect 12023 3009 12032 3043
rect 11980 3000 12032 3009
rect 17316 3000 17368 3052
rect 11796 2932 11848 2984
rect 16948 2975 17000 2984
rect 16948 2941 16957 2975
rect 16957 2941 16991 2975
rect 16991 2941 17000 2975
rect 16948 2932 17000 2941
rect 7380 2864 7432 2916
rect 9680 2864 9732 2916
rect 13452 2907 13504 2916
rect 20 2796 72 2848
rect 1492 2796 1544 2848
rect 2596 2796 2648 2848
rect 8484 2839 8536 2848
rect 8484 2805 8493 2839
rect 8493 2805 8527 2839
rect 8527 2805 8536 2839
rect 8484 2796 8536 2805
rect 13452 2873 13461 2907
rect 13461 2873 13495 2907
rect 13495 2873 13504 2907
rect 13452 2864 13504 2873
rect 17408 2796 17460 2848
rect 18052 3000 18104 3052
rect 20628 3000 20680 3052
rect 21640 3068 21692 3120
rect 23388 3145 23397 3179
rect 23397 3145 23431 3179
rect 23431 3145 23440 3179
rect 23388 3136 23440 3145
rect 24216 3068 24268 3120
rect 21732 3000 21784 3052
rect 24308 3043 24360 3052
rect 24308 3009 24317 3043
rect 24317 3009 24351 3043
rect 24351 3009 24360 3043
rect 24308 3000 24360 3009
rect 26884 3068 26936 3120
rect 27344 3068 27396 3120
rect 17960 2932 18012 2984
rect 20904 2932 20956 2984
rect 23664 2932 23716 2984
rect 24400 2932 24452 2984
rect 26148 2975 26200 2984
rect 26148 2941 26157 2975
rect 26157 2941 26191 2975
rect 26191 2941 26200 2975
rect 26148 2932 26200 2941
rect 27252 3000 27304 3052
rect 28356 3043 28408 3052
rect 28356 3009 28365 3043
rect 28365 3009 28399 3043
rect 28399 3009 28408 3043
rect 28356 3000 28408 3009
rect 33876 3111 33928 3120
rect 33048 3043 33100 3052
rect 33048 3009 33057 3043
rect 33057 3009 33091 3043
rect 33091 3009 33100 3043
rect 33048 3000 33100 3009
rect 33232 3043 33284 3052
rect 33232 3009 33241 3043
rect 33241 3009 33275 3043
rect 33275 3009 33284 3043
rect 33232 3000 33284 3009
rect 33416 3043 33468 3052
rect 33416 3009 33425 3043
rect 33425 3009 33459 3043
rect 33459 3009 33468 3043
rect 33416 3000 33468 3009
rect 33876 3077 33885 3111
rect 33885 3077 33919 3111
rect 33919 3077 33928 3111
rect 33876 3068 33928 3077
rect 34244 3111 34296 3120
rect 34244 3077 34253 3111
rect 34253 3077 34287 3111
rect 34287 3077 34296 3111
rect 34244 3068 34296 3077
rect 36360 3136 36412 3188
rect 40224 3136 40276 3188
rect 41696 3179 41748 3188
rect 41696 3145 41705 3179
rect 41705 3145 41739 3179
rect 41739 3145 41748 3179
rect 41696 3136 41748 3145
rect 42432 3179 42484 3188
rect 42432 3145 42441 3179
rect 42441 3145 42475 3179
rect 42475 3145 42484 3179
rect 42432 3136 42484 3145
rect 43168 3136 43220 3188
rect 57152 3136 57204 3188
rect 41328 3068 41380 3120
rect 42616 3111 42668 3120
rect 42616 3077 42643 3111
rect 42643 3077 42668 3111
rect 42616 3068 42668 3077
rect 35808 3000 35860 3052
rect 26332 2932 26384 2984
rect 20536 2864 20588 2916
rect 23572 2907 23624 2916
rect 21732 2796 21784 2848
rect 21916 2839 21968 2848
rect 21916 2805 21925 2839
rect 21925 2805 21959 2839
rect 21959 2805 21968 2839
rect 21916 2796 21968 2805
rect 23572 2873 23581 2907
rect 23581 2873 23615 2907
rect 23615 2873 23624 2907
rect 23572 2864 23624 2873
rect 27344 2864 27396 2916
rect 32588 2864 32640 2916
rect 26516 2796 26568 2848
rect 31576 2796 31628 2848
rect 33416 2796 33468 2848
rect 37372 3000 37424 3052
rect 37464 2932 37516 2984
rect 40040 3000 40092 3052
rect 40868 3043 40920 3052
rect 40868 3009 40877 3043
rect 40877 3009 40911 3043
rect 40911 3009 40920 3043
rect 40868 3000 40920 3009
rect 39948 2864 40000 2916
rect 41696 2932 41748 2984
rect 43076 3068 43128 3120
rect 45100 3068 45152 3120
rect 43444 3000 43496 3052
rect 43812 2975 43864 2984
rect 43812 2941 43821 2975
rect 43821 2941 43855 2975
rect 43855 2941 43864 2975
rect 43812 2932 43864 2941
rect 45192 3043 45244 3052
rect 45192 3009 45201 3043
rect 45201 3009 45235 3043
rect 45235 3009 45244 3043
rect 45192 3000 45244 3009
rect 40132 2796 40184 2848
rect 42248 2796 42300 2848
rect 52736 2864 52788 2916
rect 56048 2796 56100 2848
rect 57244 2839 57296 2848
rect 57244 2805 57253 2839
rect 57253 2805 57287 2839
rect 57287 2805 57296 2839
rect 57244 2796 57296 2805
rect 59912 2796 59964 2848
rect 4214 2694 4266 2746
rect 4278 2694 4330 2746
rect 4342 2694 4394 2746
rect 4406 2694 4458 2746
rect 4470 2694 4522 2746
rect 34934 2694 34986 2746
rect 34998 2694 35050 2746
rect 35062 2694 35114 2746
rect 35126 2694 35178 2746
rect 35190 2694 35242 2746
rect 4896 2592 4948 2644
rect 5724 2456 5776 2508
rect 21272 2592 21324 2644
rect 22560 2592 22612 2644
rect 23848 2592 23900 2644
rect 24216 2592 24268 2644
rect 26884 2592 26936 2644
rect 27068 2592 27120 2644
rect 28080 2592 28132 2644
rect 8760 2524 8812 2576
rect 8116 2499 8168 2508
rect 8116 2465 8125 2499
rect 8125 2465 8159 2499
rect 8159 2465 8168 2499
rect 8116 2456 8168 2465
rect 10140 2456 10192 2508
rect 10508 2456 10560 2508
rect 20628 2456 20680 2508
rect 21088 2499 21140 2508
rect 1492 2431 1544 2440
rect 1492 2397 1501 2431
rect 1501 2397 1535 2431
rect 1535 2397 1544 2431
rect 1492 2388 1544 2397
rect 1952 2388 2004 2440
rect 2596 2431 2648 2440
rect 2596 2397 2605 2431
rect 2605 2397 2639 2431
rect 2639 2397 2648 2431
rect 2596 2388 2648 2397
rect 5080 2388 5132 2440
rect 7748 2388 7800 2440
rect 8484 2388 8536 2440
rect 9680 2388 9732 2440
rect 13452 2388 13504 2440
rect 15476 2388 15528 2440
rect 18420 2431 18472 2440
rect 18420 2397 18429 2431
rect 18429 2397 18463 2431
rect 18463 2397 18472 2431
rect 18420 2388 18472 2397
rect 19156 2388 19208 2440
rect 20812 2431 20864 2440
rect 19984 2320 20036 2372
rect 20812 2397 20821 2431
rect 20821 2397 20855 2431
rect 20855 2397 20864 2431
rect 20812 2388 20864 2397
rect 21088 2465 21097 2499
rect 21097 2465 21131 2499
rect 21131 2465 21140 2499
rect 21088 2456 21140 2465
rect 21916 2388 21968 2440
rect 3884 2252 3936 2304
rect 11612 2252 11664 2304
rect 12532 2295 12584 2304
rect 12532 2261 12541 2295
rect 12541 2261 12575 2295
rect 12575 2261 12584 2295
rect 12532 2252 12584 2261
rect 13544 2252 13596 2304
rect 18052 2252 18104 2304
rect 20168 2295 20220 2304
rect 20168 2261 20177 2295
rect 20177 2261 20211 2295
rect 20211 2261 20220 2295
rect 20168 2252 20220 2261
rect 23664 2456 23716 2508
rect 25780 2456 25832 2508
rect 25964 2499 26016 2508
rect 25964 2465 25973 2499
rect 25973 2465 26007 2499
rect 26007 2465 26016 2499
rect 25964 2456 26016 2465
rect 23756 2431 23808 2440
rect 23756 2397 23765 2431
rect 23765 2397 23799 2431
rect 23799 2397 23808 2431
rect 23756 2388 23808 2397
rect 25872 2431 25924 2440
rect 25872 2397 25881 2431
rect 25881 2397 25915 2431
rect 25915 2397 25924 2431
rect 25872 2388 25924 2397
rect 26332 2456 26384 2508
rect 26700 2456 26752 2508
rect 26884 2456 26936 2508
rect 33048 2592 33100 2644
rect 39948 2635 40000 2644
rect 39948 2601 39957 2635
rect 39957 2601 39991 2635
rect 39991 2601 40000 2635
rect 39948 2592 40000 2601
rect 46112 2592 46164 2644
rect 50988 2592 51040 2644
rect 51172 2635 51224 2644
rect 51172 2601 51181 2635
rect 51181 2601 51215 2635
rect 51215 2601 51224 2635
rect 51172 2592 51224 2601
rect 52368 2592 52420 2644
rect 55864 2592 55916 2644
rect 32680 2524 32732 2576
rect 48504 2524 48556 2576
rect 26516 2388 26568 2440
rect 26976 2431 27028 2440
rect 26976 2397 26985 2431
rect 26985 2397 27019 2431
rect 27019 2397 27028 2431
rect 26976 2388 27028 2397
rect 27712 2388 27764 2440
rect 28448 2388 28500 2440
rect 31576 2431 31628 2440
rect 23848 2320 23900 2372
rect 26700 2320 26752 2372
rect 27252 2320 27304 2372
rect 29644 2320 29696 2372
rect 31576 2397 31585 2431
rect 31585 2397 31619 2431
rect 31619 2397 31628 2431
rect 31576 2388 31628 2397
rect 32588 2431 32640 2440
rect 32588 2397 32597 2431
rect 32597 2397 32631 2431
rect 32631 2397 32640 2431
rect 32588 2388 32640 2397
rect 33232 2431 33284 2440
rect 33232 2397 33241 2431
rect 33241 2397 33275 2431
rect 33275 2397 33284 2431
rect 33232 2388 33284 2397
rect 33416 2431 33468 2440
rect 33416 2397 33425 2431
rect 33425 2397 33459 2431
rect 33459 2397 33468 2431
rect 33416 2388 33468 2397
rect 30104 2295 30156 2304
rect 30104 2261 30113 2295
rect 30113 2261 30147 2295
rect 30147 2261 30156 2295
rect 30104 2252 30156 2261
rect 32680 2252 32732 2304
rect 36084 2388 36136 2440
rect 40132 2431 40184 2440
rect 40132 2397 40141 2431
rect 40141 2397 40175 2431
rect 40175 2397 40184 2431
rect 40132 2388 40184 2397
rect 40224 2431 40276 2440
rect 40224 2397 40233 2431
rect 40233 2397 40267 2431
rect 40267 2397 40276 2431
rect 40224 2388 40276 2397
rect 41604 2388 41656 2440
rect 43352 2388 43404 2440
rect 42708 2363 42760 2372
rect 42708 2329 42717 2363
rect 42717 2329 42751 2363
rect 42751 2329 42760 2363
rect 42708 2320 42760 2329
rect 46112 2431 46164 2440
rect 46112 2397 46121 2431
rect 46121 2397 46155 2431
rect 46155 2397 46164 2431
rect 46112 2388 46164 2397
rect 52552 2524 52604 2576
rect 51172 2388 51224 2440
rect 52736 2431 52788 2440
rect 52736 2397 52745 2431
rect 52745 2397 52779 2431
rect 52779 2397 52788 2431
rect 52736 2388 52788 2397
rect 54208 2388 54260 2440
rect 56048 2388 56100 2440
rect 57888 2431 57940 2440
rect 57888 2397 57897 2431
rect 57897 2397 57931 2431
rect 57931 2397 57940 2431
rect 57888 2388 57940 2397
rect 49792 2320 49844 2372
rect 57244 2363 57296 2372
rect 57244 2329 57253 2363
rect 57253 2329 57287 2363
rect 57287 2329 57296 2363
rect 57244 2320 57296 2329
rect 34152 2295 34204 2304
rect 34152 2261 34161 2295
rect 34161 2261 34195 2295
rect 34195 2261 34204 2295
rect 34152 2252 34204 2261
rect 37556 2295 37608 2304
rect 37556 2261 37565 2295
rect 37565 2261 37599 2295
rect 37599 2261 37608 2295
rect 37556 2252 37608 2261
rect 38016 2252 38068 2304
rect 40040 2252 40092 2304
rect 41880 2295 41932 2304
rect 41880 2261 41889 2295
rect 41889 2261 41923 2295
rect 41923 2261 41932 2295
rect 41880 2252 41932 2261
rect 43352 2295 43404 2304
rect 43352 2261 43361 2295
rect 43361 2261 43395 2295
rect 43395 2261 43404 2295
rect 43352 2252 43404 2261
rect 43812 2252 43864 2304
rect 45744 2252 45796 2304
rect 47676 2252 47728 2304
rect 50160 2252 50212 2304
rect 52184 2252 52236 2304
rect 57980 2252 58032 2304
rect 19574 2150 19626 2202
rect 19638 2150 19690 2202
rect 19702 2150 19754 2202
rect 19766 2150 19818 2202
rect 19830 2150 19882 2202
rect 50294 2150 50346 2202
rect 50358 2150 50410 2202
rect 50422 2150 50474 2202
rect 50486 2150 50538 2202
rect 50550 2150 50602 2202
rect 5172 2048 5224 2100
rect 37556 2048 37608 2100
rect 48504 2048 48556 2100
rect 54576 2048 54628 2100
rect 12532 1980 12584 2032
rect 46480 1980 46532 2032
rect 18420 1912 18472 1964
rect 26608 1912 26660 1964
rect 42708 1912 42760 1964
rect 48780 1912 48832 1964
rect 14188 1844 14240 1896
rect 30104 1844 30156 1896
rect 20168 1776 20220 1828
rect 43352 1776 43404 1828
rect 26240 1708 26292 1760
rect 26976 1708 27028 1760
rect 27528 1708 27580 1760
rect 49792 1708 49844 1760
<< metal2 >>
rect 18 39200 74 40000
rect 1950 39200 2006 40000
rect 3882 39200 3938 40000
rect 5814 39200 5870 40000
rect 7746 39200 7802 40000
rect 9678 39200 9734 40000
rect 12254 39200 12310 40000
rect 14186 39200 14242 40000
rect 16118 39200 16174 40000
rect 16224 39222 16528 39250
rect 32 37126 60 39200
rect 1490 38176 1546 38185
rect 1490 38111 1546 38120
rect 20 37120 72 37126
rect 20 37062 72 37068
rect 1504 36922 1532 38111
rect 1964 37126 1992 39200
rect 3896 37262 3924 39200
rect 4214 37564 4522 37584
rect 4214 37562 4220 37564
rect 4276 37562 4300 37564
rect 4356 37562 4380 37564
rect 4436 37562 4460 37564
rect 4516 37562 4522 37564
rect 4276 37510 4278 37562
rect 4458 37510 4460 37562
rect 4214 37508 4220 37510
rect 4276 37508 4300 37510
rect 4356 37508 4380 37510
rect 4436 37508 4460 37510
rect 4516 37508 4522 37510
rect 4214 37488 4522 37508
rect 5724 37392 5776 37398
rect 5724 37334 5776 37340
rect 5828 37346 5856 39200
rect 4620 37324 4672 37330
rect 4620 37266 4672 37272
rect 2412 37256 2464 37262
rect 2412 37198 2464 37204
rect 3884 37256 3936 37262
rect 3884 37198 3936 37204
rect 1952 37120 2004 37126
rect 1952 37062 2004 37068
rect 1492 36916 1544 36922
rect 1492 36858 1544 36864
rect 2044 36780 2096 36786
rect 2044 36722 2096 36728
rect 1676 36168 1728 36174
rect 1490 36136 1546 36145
rect 1676 36110 1728 36116
rect 1490 36071 1546 36080
rect 1504 36038 1532 36071
rect 1492 36032 1544 36038
rect 1492 35974 1544 35980
rect 1584 33516 1636 33522
rect 1584 33458 1636 33464
rect 1596 33425 1624 33458
rect 1582 33416 1638 33425
rect 1582 33351 1638 33360
rect 1596 33114 1624 33351
rect 1584 33108 1636 33114
rect 1584 33050 1636 33056
rect 1688 32026 1716 36110
rect 1768 33312 1820 33318
rect 1768 33254 1820 33260
rect 1676 32020 1728 32026
rect 1676 31962 1728 31968
rect 1584 31748 1636 31754
rect 1584 31690 1636 31696
rect 1596 31414 1624 31690
rect 1584 31408 1636 31414
rect 1582 31376 1584 31385
rect 1636 31376 1638 31385
rect 1582 31311 1638 31320
rect 1492 29504 1544 29510
rect 1492 29446 1544 29452
rect 1504 29345 1532 29446
rect 1490 29336 1546 29345
rect 1490 29271 1546 29280
rect 1400 21548 1452 21554
rect 1400 21490 1452 21496
rect 1412 21185 1440 21490
rect 1584 21344 1636 21350
rect 1584 21286 1636 21292
rect 1398 21176 1454 21185
rect 1398 21111 1400 21120
rect 1452 21111 1454 21120
rect 1400 21082 1452 21088
rect 1492 20528 1544 20534
rect 1492 20470 1544 20476
rect 1400 19372 1452 19378
rect 1400 19314 1452 19320
rect 1412 19145 1440 19314
rect 1398 19136 1454 19145
rect 1398 19071 1454 19080
rect 1412 18970 1440 19071
rect 1400 18964 1452 18970
rect 1400 18906 1452 18912
rect 1504 14618 1532 20470
rect 1596 18766 1624 21286
rect 1584 18760 1636 18766
rect 1584 18702 1636 18708
rect 1596 18358 1624 18702
rect 1584 18352 1636 18358
rect 1584 18294 1636 18300
rect 1584 17604 1636 17610
rect 1584 17546 1636 17552
rect 1492 14612 1544 14618
rect 1492 14554 1544 14560
rect 1400 14408 1452 14414
rect 1398 14376 1400 14385
rect 1452 14376 1454 14385
rect 1398 14311 1454 14320
rect 1596 12986 1624 17546
rect 1780 16250 1808 33254
rect 1952 31816 2004 31822
rect 1952 31758 2004 31764
rect 1858 27296 1914 27305
rect 1858 27231 1914 27240
rect 1872 27062 1900 27231
rect 1860 27056 1912 27062
rect 1860 26998 1912 27004
rect 1872 26586 1900 26998
rect 1860 26580 1912 26586
rect 1860 26522 1912 26528
rect 1858 25256 1914 25265
rect 1858 25191 1860 25200
rect 1912 25191 1914 25200
rect 1860 25162 1912 25168
rect 1872 24954 1900 25162
rect 1860 24948 1912 24954
rect 1860 24890 1912 24896
rect 1858 23216 1914 23225
rect 1858 23151 1914 23160
rect 1872 23118 1900 23151
rect 1860 23112 1912 23118
rect 1860 23054 1912 23060
rect 1872 22778 1900 23054
rect 1860 22772 1912 22778
rect 1860 22714 1912 22720
rect 1964 20262 1992 31758
rect 2056 27606 2084 36722
rect 2228 32564 2280 32570
rect 2228 32506 2280 32512
rect 2240 29850 2268 32506
rect 2228 29844 2280 29850
rect 2228 29786 2280 29792
rect 2240 29646 2268 29786
rect 2228 29640 2280 29646
rect 2228 29582 2280 29588
rect 2044 27600 2096 27606
rect 2044 27542 2096 27548
rect 2042 23080 2098 23089
rect 2042 23015 2044 23024
rect 2096 23015 2098 23024
rect 2044 22986 2096 22992
rect 2136 22024 2188 22030
rect 2136 21966 2188 21972
rect 2148 20466 2176 21966
rect 2228 21548 2280 21554
rect 2228 21490 2280 21496
rect 2240 20534 2268 21490
rect 2228 20528 2280 20534
rect 2228 20470 2280 20476
rect 2136 20460 2188 20466
rect 2136 20402 2188 20408
rect 1952 20256 2004 20262
rect 1952 20198 2004 20204
rect 2424 18426 2452 37198
rect 3896 36922 3924 37198
rect 3884 36916 3936 36922
rect 3884 36858 3936 36864
rect 4068 36916 4120 36922
rect 4068 36858 4120 36864
rect 3240 31816 3292 31822
rect 3240 31758 3292 31764
rect 3252 31385 3280 31758
rect 3238 31376 3294 31385
rect 3238 31311 3294 31320
rect 3332 29708 3384 29714
rect 3332 29650 3384 29656
rect 3344 29170 3372 29650
rect 3332 29164 3384 29170
rect 3332 29106 3384 29112
rect 3344 28014 3372 29106
rect 2964 28008 3016 28014
rect 2964 27950 3016 27956
rect 3056 28008 3108 28014
rect 3056 27950 3108 27956
rect 3332 28008 3384 28014
rect 3332 27950 3384 27956
rect 2780 27532 2832 27538
rect 2780 27474 2832 27480
rect 2792 26042 2820 27474
rect 2780 26036 2832 26042
rect 2780 25978 2832 25984
rect 2504 25288 2556 25294
rect 2504 25230 2556 25236
rect 2516 24818 2544 25230
rect 2596 25220 2648 25226
rect 2596 25162 2648 25168
rect 2608 24818 2636 25162
rect 2504 24812 2556 24818
rect 2504 24754 2556 24760
rect 2596 24812 2648 24818
rect 2596 24754 2648 24760
rect 2516 23730 2544 24754
rect 2608 23798 2636 24754
rect 2596 23792 2648 23798
rect 2596 23734 2648 23740
rect 2504 23724 2556 23730
rect 2504 23666 2556 23672
rect 2504 20936 2556 20942
rect 2504 20878 2556 20884
rect 2516 20466 2544 20878
rect 2504 20460 2556 20466
rect 2504 20402 2556 20408
rect 2412 18420 2464 18426
rect 2412 18362 2464 18368
rect 2044 18284 2096 18290
rect 2044 18226 2096 18232
rect 2056 17610 2084 18226
rect 2044 17604 2096 17610
rect 2044 17546 2096 17552
rect 1860 16992 1912 16998
rect 1860 16934 1912 16940
rect 1872 16522 1900 16934
rect 1860 16516 1912 16522
rect 1860 16458 1912 16464
rect 1872 16425 1900 16458
rect 1858 16416 1914 16425
rect 1858 16351 1914 16360
rect 1768 16244 1820 16250
rect 1768 16186 1820 16192
rect 1584 12980 1636 12986
rect 1584 12922 1636 12928
rect 1400 12844 1452 12850
rect 1400 12786 1452 12792
rect 1412 12374 1440 12786
rect 2608 12782 2636 23734
rect 2780 22024 2832 22030
rect 2780 21966 2832 21972
rect 2688 21888 2740 21894
rect 2688 21830 2740 21836
rect 2700 20942 2728 21830
rect 2792 21486 2820 21966
rect 2872 21956 2924 21962
rect 2872 21898 2924 21904
rect 2884 21690 2912 21898
rect 2872 21684 2924 21690
rect 2872 21626 2924 21632
rect 2780 21480 2832 21486
rect 2780 21422 2832 21428
rect 2688 20936 2740 20942
rect 2688 20878 2740 20884
rect 2872 19780 2924 19786
rect 2872 19722 2924 19728
rect 2884 19514 2912 19722
rect 2872 19508 2924 19514
rect 2872 19450 2924 19456
rect 2688 19168 2740 19174
rect 2688 19110 2740 19116
rect 2700 18873 2728 19110
rect 2686 18864 2742 18873
rect 2686 18799 2742 18808
rect 2780 18284 2832 18290
rect 2780 18226 2832 18232
rect 2792 16454 2820 18226
rect 2872 17128 2924 17134
rect 2872 17070 2924 17076
rect 2884 16726 2912 17070
rect 2872 16720 2924 16726
rect 2872 16662 2924 16668
rect 2780 16448 2832 16454
rect 2780 16390 2832 16396
rect 2688 16176 2740 16182
rect 2688 16118 2740 16124
rect 2700 15706 2728 16118
rect 2780 16108 2832 16114
rect 2780 16050 2832 16056
rect 2688 15700 2740 15706
rect 2688 15642 2740 15648
rect 2700 15094 2728 15642
rect 2688 15088 2740 15094
rect 2688 15030 2740 15036
rect 2792 15026 2820 16050
rect 2884 15978 2912 16662
rect 2872 15972 2924 15978
rect 2872 15914 2924 15920
rect 2780 15020 2832 15026
rect 2780 14962 2832 14968
rect 2596 12776 2648 12782
rect 2596 12718 2648 12724
rect 1400 12368 1452 12374
rect 1398 12336 1400 12345
rect 1452 12336 1454 12345
rect 1398 12271 1454 12280
rect 2792 10810 2820 14962
rect 2872 12844 2924 12850
rect 2872 12786 2924 12792
rect 2884 11354 2912 12786
rect 2872 11348 2924 11354
rect 2872 11290 2924 11296
rect 2872 11144 2924 11150
rect 2872 11086 2924 11092
rect 2780 10804 2832 10810
rect 2780 10746 2832 10752
rect 1400 10668 1452 10674
rect 1400 10610 1452 10616
rect 1412 10305 1440 10610
rect 1398 10296 1454 10305
rect 1398 10231 1400 10240
rect 1452 10231 1454 10240
rect 1400 10202 1452 10208
rect 2884 10062 2912 11086
rect 2872 10056 2924 10062
rect 2872 9998 2924 10004
rect 2976 8634 3004 27950
rect 3068 27674 3096 27950
rect 3056 27668 3108 27674
rect 3056 27610 3108 27616
rect 3148 26580 3200 26586
rect 3148 26522 3200 26528
rect 3160 25922 3188 26522
rect 3068 25906 3188 25922
rect 3068 25900 3200 25906
rect 3068 25894 3148 25900
rect 3068 25430 3096 25894
rect 3148 25842 3200 25848
rect 3148 25764 3200 25770
rect 3148 25706 3200 25712
rect 3056 25424 3108 25430
rect 3056 25366 3108 25372
rect 3068 24954 3096 25366
rect 3160 25294 3188 25706
rect 3148 25288 3200 25294
rect 3148 25230 3200 25236
rect 3056 24948 3108 24954
rect 3056 24890 3108 24896
rect 3160 24818 3188 25230
rect 3148 24812 3200 24818
rect 3148 24754 3200 24760
rect 3160 22094 3188 24754
rect 3160 22066 3280 22094
rect 3148 21888 3200 21894
rect 3148 21830 3200 21836
rect 3160 21146 3188 21830
rect 3148 21140 3200 21146
rect 3148 21082 3200 21088
rect 3056 18284 3108 18290
rect 3056 18226 3108 18232
rect 3068 17338 3096 18226
rect 3056 17332 3108 17338
rect 3056 17274 3108 17280
rect 3252 13462 3280 22066
rect 3344 16794 3372 27950
rect 3976 27464 4028 27470
rect 3976 27406 4028 27412
rect 3988 25770 4016 27406
rect 4080 26586 4108 36858
rect 4214 36476 4522 36496
rect 4214 36474 4220 36476
rect 4276 36474 4300 36476
rect 4356 36474 4380 36476
rect 4436 36474 4460 36476
rect 4516 36474 4522 36476
rect 4276 36422 4278 36474
rect 4458 36422 4460 36474
rect 4214 36420 4220 36422
rect 4276 36420 4300 36422
rect 4356 36420 4380 36422
rect 4436 36420 4460 36422
rect 4516 36420 4522 36422
rect 4214 36400 4522 36420
rect 4214 35388 4522 35408
rect 4214 35386 4220 35388
rect 4276 35386 4300 35388
rect 4356 35386 4380 35388
rect 4436 35386 4460 35388
rect 4516 35386 4522 35388
rect 4276 35334 4278 35386
rect 4458 35334 4460 35386
rect 4214 35332 4220 35334
rect 4276 35332 4300 35334
rect 4356 35332 4380 35334
rect 4436 35332 4460 35334
rect 4516 35332 4522 35334
rect 4214 35312 4522 35332
rect 4214 34300 4522 34320
rect 4214 34298 4220 34300
rect 4276 34298 4300 34300
rect 4356 34298 4380 34300
rect 4436 34298 4460 34300
rect 4516 34298 4522 34300
rect 4276 34246 4278 34298
rect 4458 34246 4460 34298
rect 4214 34244 4220 34246
rect 4276 34244 4300 34246
rect 4356 34244 4380 34246
rect 4436 34244 4460 34246
rect 4516 34244 4522 34246
rect 4214 34224 4522 34244
rect 4214 33212 4522 33232
rect 4214 33210 4220 33212
rect 4276 33210 4300 33212
rect 4356 33210 4380 33212
rect 4436 33210 4460 33212
rect 4516 33210 4522 33212
rect 4276 33158 4278 33210
rect 4458 33158 4460 33210
rect 4214 33156 4220 33158
rect 4276 33156 4300 33158
rect 4356 33156 4380 33158
rect 4436 33156 4460 33158
rect 4516 33156 4522 33158
rect 4214 33136 4522 33156
rect 4214 32124 4522 32144
rect 4214 32122 4220 32124
rect 4276 32122 4300 32124
rect 4356 32122 4380 32124
rect 4436 32122 4460 32124
rect 4516 32122 4522 32124
rect 4276 32070 4278 32122
rect 4458 32070 4460 32122
rect 4214 32068 4220 32070
rect 4276 32068 4300 32070
rect 4356 32068 4380 32070
rect 4436 32068 4460 32070
rect 4516 32068 4522 32070
rect 4214 32048 4522 32068
rect 4214 31036 4522 31056
rect 4214 31034 4220 31036
rect 4276 31034 4300 31036
rect 4356 31034 4380 31036
rect 4436 31034 4460 31036
rect 4516 31034 4522 31036
rect 4276 30982 4278 31034
rect 4458 30982 4460 31034
rect 4214 30980 4220 30982
rect 4276 30980 4300 30982
rect 4356 30980 4380 30982
rect 4436 30980 4460 30982
rect 4516 30980 4522 30982
rect 4214 30960 4522 30980
rect 4214 29948 4522 29968
rect 4214 29946 4220 29948
rect 4276 29946 4300 29948
rect 4356 29946 4380 29948
rect 4436 29946 4460 29948
rect 4516 29946 4522 29948
rect 4276 29894 4278 29946
rect 4458 29894 4460 29946
rect 4214 29892 4220 29894
rect 4276 29892 4300 29894
rect 4356 29892 4380 29894
rect 4436 29892 4460 29894
rect 4516 29892 4522 29894
rect 4214 29872 4522 29892
rect 4344 29504 4396 29510
rect 4344 29446 4396 29452
rect 4356 29238 4384 29446
rect 4344 29232 4396 29238
rect 4344 29174 4396 29180
rect 4214 28860 4522 28880
rect 4214 28858 4220 28860
rect 4276 28858 4300 28860
rect 4356 28858 4380 28860
rect 4436 28858 4460 28860
rect 4516 28858 4522 28860
rect 4276 28806 4278 28858
rect 4458 28806 4460 28858
rect 4214 28804 4220 28806
rect 4276 28804 4300 28806
rect 4356 28804 4380 28806
rect 4436 28804 4460 28806
rect 4516 28804 4522 28806
rect 4214 28784 4522 28804
rect 4214 27772 4522 27792
rect 4214 27770 4220 27772
rect 4276 27770 4300 27772
rect 4356 27770 4380 27772
rect 4436 27770 4460 27772
rect 4516 27770 4522 27772
rect 4276 27718 4278 27770
rect 4458 27718 4460 27770
rect 4214 27716 4220 27718
rect 4276 27716 4300 27718
rect 4356 27716 4380 27718
rect 4436 27716 4460 27718
rect 4516 27716 4522 27718
rect 4214 27696 4522 27716
rect 4214 26684 4522 26704
rect 4214 26682 4220 26684
rect 4276 26682 4300 26684
rect 4356 26682 4380 26684
rect 4436 26682 4460 26684
rect 4516 26682 4522 26684
rect 4276 26630 4278 26682
rect 4458 26630 4460 26682
rect 4214 26628 4220 26630
rect 4276 26628 4300 26630
rect 4356 26628 4380 26630
rect 4436 26628 4460 26630
rect 4516 26628 4522 26630
rect 4214 26608 4522 26628
rect 4068 26580 4120 26586
rect 4068 26522 4120 26528
rect 4068 26036 4120 26042
rect 4068 25978 4120 25984
rect 3976 25764 4028 25770
rect 3976 25706 4028 25712
rect 3424 25696 3476 25702
rect 3424 25638 3476 25644
rect 3436 24818 3464 25638
rect 3516 25424 3568 25430
rect 3516 25366 3568 25372
rect 3424 24812 3476 24818
rect 3424 24754 3476 24760
rect 3528 22094 3556 25366
rect 3988 25362 4016 25706
rect 4080 25362 4108 25978
rect 4214 25596 4522 25616
rect 4214 25594 4220 25596
rect 4276 25594 4300 25596
rect 4356 25594 4380 25596
rect 4436 25594 4460 25596
rect 4516 25594 4522 25596
rect 4276 25542 4278 25594
rect 4458 25542 4460 25594
rect 4214 25540 4220 25542
rect 4276 25540 4300 25542
rect 4356 25540 4380 25542
rect 4436 25540 4460 25542
rect 4516 25540 4522 25542
rect 4214 25520 4522 25540
rect 3976 25356 4028 25362
rect 3976 25298 4028 25304
rect 4068 25356 4120 25362
rect 4068 25298 4120 25304
rect 3792 25288 3844 25294
rect 4252 25288 4304 25294
rect 4172 25248 4252 25276
rect 4172 25242 4200 25248
rect 3792 25230 3844 25236
rect 3804 24750 3832 25230
rect 4080 25214 4200 25242
rect 4252 25230 4304 25236
rect 3884 24948 3936 24954
rect 3884 24890 3936 24896
rect 3792 24744 3844 24750
rect 3792 24686 3844 24692
rect 3608 24608 3660 24614
rect 3608 24550 3660 24556
rect 3620 22642 3648 24550
rect 3896 24410 3924 24890
rect 3884 24404 3936 24410
rect 3884 24346 3936 24352
rect 4080 23798 4108 25214
rect 4214 24508 4522 24528
rect 4214 24506 4220 24508
rect 4276 24506 4300 24508
rect 4356 24506 4380 24508
rect 4436 24506 4460 24508
rect 4516 24506 4522 24508
rect 4276 24454 4278 24506
rect 4458 24454 4460 24506
rect 4214 24452 4220 24454
rect 4276 24452 4300 24454
rect 4356 24452 4380 24454
rect 4436 24452 4460 24454
rect 4516 24452 4522 24454
rect 4214 24432 4522 24452
rect 4068 23792 4120 23798
rect 4068 23734 4120 23740
rect 4080 22710 4108 23734
rect 4214 23420 4522 23440
rect 4214 23418 4220 23420
rect 4276 23418 4300 23420
rect 4356 23418 4380 23420
rect 4436 23418 4460 23420
rect 4516 23418 4522 23420
rect 4276 23366 4278 23418
rect 4458 23366 4460 23418
rect 4214 23364 4220 23366
rect 4276 23364 4300 23366
rect 4356 23364 4380 23366
rect 4436 23364 4460 23366
rect 4516 23364 4522 23366
rect 4214 23344 4522 23364
rect 4632 23118 4660 37266
rect 5540 35556 5592 35562
rect 5540 35498 5592 35504
rect 5448 30252 5500 30258
rect 5448 30194 5500 30200
rect 5460 29646 5488 30194
rect 5448 29640 5500 29646
rect 5448 29582 5500 29588
rect 4896 29504 4948 29510
rect 4896 29446 4948 29452
rect 4908 27946 4936 29446
rect 4896 27940 4948 27946
rect 4896 27882 4948 27888
rect 5460 26858 5488 29582
rect 5552 27470 5580 35498
rect 5736 29714 5764 37334
rect 5828 37318 5948 37346
rect 5816 37256 5868 37262
rect 5816 37198 5868 37204
rect 5828 36718 5856 37198
rect 5920 37126 5948 37318
rect 7760 37262 7788 39200
rect 9692 37262 9720 39200
rect 12268 37330 12296 39200
rect 14200 37330 14228 39200
rect 16132 39114 16160 39200
rect 16224 39114 16252 39222
rect 16132 39086 16252 39114
rect 12256 37324 12308 37330
rect 12256 37266 12308 37272
rect 14188 37324 14240 37330
rect 14188 37266 14240 37272
rect 7748 37256 7800 37262
rect 7748 37198 7800 37204
rect 9680 37256 9732 37262
rect 9680 37198 9732 37204
rect 7104 37188 7156 37194
rect 7104 37130 7156 37136
rect 5908 37120 5960 37126
rect 5908 37062 5960 37068
rect 6736 36780 6788 36786
rect 6736 36722 6788 36728
rect 5816 36712 5868 36718
rect 5816 36654 5868 36660
rect 6644 36576 6696 36582
rect 6644 36518 6696 36524
rect 6656 36310 6684 36518
rect 6644 36304 6696 36310
rect 6644 36246 6696 36252
rect 6656 35834 6684 36246
rect 6748 35834 6776 36722
rect 7116 36718 7144 37130
rect 8024 37120 8076 37126
rect 8024 37062 8076 37068
rect 11520 37120 11572 37126
rect 11520 37062 11572 37068
rect 7472 36780 7524 36786
rect 7472 36722 7524 36728
rect 7104 36712 7156 36718
rect 7104 36654 7156 36660
rect 6644 35828 6696 35834
rect 6644 35770 6696 35776
rect 6736 35828 6788 35834
rect 6736 35770 6788 35776
rect 7484 35766 7512 36722
rect 8036 36174 8064 37062
rect 8300 36780 8352 36786
rect 8300 36722 8352 36728
rect 8576 36780 8628 36786
rect 8576 36722 8628 36728
rect 8312 36378 8340 36722
rect 8300 36372 8352 36378
rect 8300 36314 8352 36320
rect 8588 36310 8616 36722
rect 8944 36372 8996 36378
rect 8944 36314 8996 36320
rect 8576 36304 8628 36310
rect 8576 36246 8628 36252
rect 8024 36168 8076 36174
rect 8024 36110 8076 36116
rect 8036 35766 8064 36110
rect 7012 35760 7064 35766
rect 7012 35702 7064 35708
rect 7472 35760 7524 35766
rect 7472 35702 7524 35708
rect 8024 35760 8076 35766
rect 8024 35702 8076 35708
rect 7024 35290 7052 35702
rect 7748 35692 7800 35698
rect 7748 35634 7800 35640
rect 8116 35692 8168 35698
rect 8116 35634 8168 35640
rect 8300 35692 8352 35698
rect 8300 35634 8352 35640
rect 7760 35290 7788 35634
rect 7932 35488 7984 35494
rect 7932 35430 7984 35436
rect 7012 35284 7064 35290
rect 7012 35226 7064 35232
rect 7748 35284 7800 35290
rect 7748 35226 7800 35232
rect 7012 35148 7064 35154
rect 7012 35090 7064 35096
rect 7024 34542 7052 35090
rect 7944 35086 7972 35430
rect 7932 35080 7984 35086
rect 7932 35022 7984 35028
rect 8024 35080 8076 35086
rect 8128 35068 8156 35634
rect 8312 35154 8340 35634
rect 8300 35148 8352 35154
rect 8300 35090 8352 35096
rect 8076 35040 8156 35068
rect 8024 35022 8076 35028
rect 8036 34932 8064 35022
rect 7944 34904 8064 34932
rect 7840 34604 7892 34610
rect 7840 34546 7892 34552
rect 7012 34536 7064 34542
rect 7012 34478 7064 34484
rect 7656 34400 7708 34406
rect 7656 34342 7708 34348
rect 7288 33856 7340 33862
rect 7288 33798 7340 33804
rect 7104 33380 7156 33386
rect 7104 33322 7156 33328
rect 7116 32910 7144 33322
rect 7300 32910 7328 33798
rect 7668 33386 7696 34342
rect 7852 33998 7880 34546
rect 7944 34542 7972 34904
rect 8312 34746 8340 35090
rect 8300 34740 8352 34746
rect 8300 34682 8352 34688
rect 7932 34536 7984 34542
rect 7932 34478 7984 34484
rect 7840 33992 7892 33998
rect 7840 33934 7892 33940
rect 7656 33380 7708 33386
rect 7656 33322 7708 33328
rect 7668 32978 7696 33322
rect 7656 32972 7708 32978
rect 7656 32914 7708 32920
rect 7104 32904 7156 32910
rect 7104 32846 7156 32852
rect 7288 32904 7340 32910
rect 7288 32846 7340 32852
rect 7116 31770 7144 32846
rect 7196 31816 7248 31822
rect 7116 31764 7196 31770
rect 7116 31758 7248 31764
rect 7116 31742 7236 31758
rect 7300 31754 7328 32846
rect 7380 32768 7432 32774
rect 7380 32710 7432 32716
rect 7392 32434 7420 32710
rect 7380 32428 7432 32434
rect 7380 32370 7432 32376
rect 7288 31748 7340 31754
rect 7116 31414 7144 31742
rect 7288 31690 7340 31696
rect 7104 31408 7156 31414
rect 7104 31350 7156 31356
rect 7196 31340 7248 31346
rect 7300 31328 7328 31690
rect 7248 31300 7328 31328
rect 7196 31282 7248 31288
rect 7564 31204 7616 31210
rect 7564 31146 7616 31152
rect 7288 30728 7340 30734
rect 7288 30670 7340 30676
rect 6920 30252 6972 30258
rect 6920 30194 6972 30200
rect 5724 29708 5776 29714
rect 5724 29650 5776 29656
rect 5736 29102 5764 29650
rect 6932 29238 6960 30194
rect 6920 29232 6972 29238
rect 6920 29174 6972 29180
rect 5724 29096 5776 29102
rect 5724 29038 5776 29044
rect 6736 28484 6788 28490
rect 6736 28426 6788 28432
rect 6748 27878 6776 28426
rect 7012 28416 7064 28422
rect 7012 28358 7064 28364
rect 7024 28150 7052 28358
rect 7012 28144 7064 28150
rect 7012 28086 7064 28092
rect 6460 27872 6512 27878
rect 6460 27814 6512 27820
rect 6736 27872 6788 27878
rect 6736 27814 6788 27820
rect 6472 27470 6500 27814
rect 5540 27464 5592 27470
rect 5540 27406 5592 27412
rect 6460 27464 6512 27470
rect 6460 27406 6512 27412
rect 5632 27396 5684 27402
rect 5632 27338 5684 27344
rect 5644 27130 5672 27338
rect 6276 27328 6328 27334
rect 6276 27270 6328 27276
rect 5632 27124 5684 27130
rect 5632 27066 5684 27072
rect 6288 26926 6316 27270
rect 6644 27124 6696 27130
rect 6644 27066 6696 27072
rect 6276 26920 6328 26926
rect 6276 26862 6328 26868
rect 5448 26852 5500 26858
rect 5448 26794 5500 26800
rect 5460 23730 5488 26794
rect 6288 26382 6316 26862
rect 6656 26790 6684 27066
rect 6748 27062 6776 27814
rect 7196 27328 7248 27334
rect 7196 27270 7248 27276
rect 6736 27056 6788 27062
rect 6736 26998 6788 27004
rect 6828 26988 6880 26994
rect 6828 26930 6880 26936
rect 7104 26988 7156 26994
rect 7208 26976 7236 27270
rect 7300 27130 7328 30670
rect 7380 29844 7432 29850
rect 7380 29786 7432 29792
rect 7392 29646 7420 29786
rect 7380 29640 7432 29646
rect 7380 29582 7432 29588
rect 7392 28966 7420 29582
rect 7472 29572 7524 29578
rect 7472 29514 7524 29520
rect 7484 29306 7512 29514
rect 7472 29300 7524 29306
rect 7472 29242 7524 29248
rect 7380 28960 7432 28966
rect 7380 28902 7432 28908
rect 7472 27872 7524 27878
rect 7472 27814 7524 27820
rect 7484 27606 7512 27814
rect 7472 27600 7524 27606
rect 7472 27542 7524 27548
rect 7288 27124 7340 27130
rect 7288 27066 7340 27072
rect 7156 26948 7236 26976
rect 7104 26930 7156 26936
rect 6644 26784 6696 26790
rect 6644 26726 6696 26732
rect 6656 26450 6684 26726
rect 6840 26586 6868 26930
rect 6828 26580 6880 26586
rect 6828 26522 6880 26528
rect 6644 26444 6696 26450
rect 6644 26386 6696 26392
rect 6276 26376 6328 26382
rect 6276 26318 6328 26324
rect 6288 26042 6316 26318
rect 6276 26036 6328 26042
rect 6276 25978 6328 25984
rect 6288 25226 6316 25978
rect 6656 25770 6684 26386
rect 6920 25900 6972 25906
rect 6920 25842 6972 25848
rect 6644 25764 6696 25770
rect 6644 25706 6696 25712
rect 6656 25498 6684 25706
rect 6644 25492 6696 25498
rect 6644 25434 6696 25440
rect 6276 25220 6328 25226
rect 6276 25162 6328 25168
rect 6828 25220 6880 25226
rect 6828 25162 6880 25168
rect 5448 23724 5500 23730
rect 5448 23666 5500 23672
rect 4804 23520 4856 23526
rect 4804 23462 4856 23468
rect 4620 23112 4672 23118
rect 4620 23054 4672 23060
rect 4632 22778 4660 23054
rect 4816 23050 4844 23462
rect 6840 23322 6868 25162
rect 6932 24206 6960 25842
rect 7012 25152 7064 25158
rect 7012 25094 7064 25100
rect 7024 24818 7052 25094
rect 7208 24818 7236 26948
rect 7470 25528 7526 25537
rect 7470 25463 7526 25472
rect 7484 24818 7512 25463
rect 7012 24812 7064 24818
rect 7012 24754 7064 24760
rect 7196 24812 7248 24818
rect 7196 24754 7248 24760
rect 7288 24812 7340 24818
rect 7288 24754 7340 24760
rect 7472 24812 7524 24818
rect 7472 24754 7524 24760
rect 7208 24614 7236 24754
rect 7196 24608 7248 24614
rect 7196 24550 7248 24556
rect 6920 24200 6972 24206
rect 6920 24142 6972 24148
rect 7012 23656 7064 23662
rect 7012 23598 7064 23604
rect 6828 23316 6880 23322
rect 6828 23258 6880 23264
rect 6184 23180 6236 23186
rect 6184 23122 6236 23128
rect 4804 23044 4856 23050
rect 4804 22986 4856 22992
rect 4620 22772 4672 22778
rect 4620 22714 4672 22720
rect 4068 22704 4120 22710
rect 4068 22646 4120 22652
rect 3608 22636 3660 22642
rect 3608 22578 3660 22584
rect 4620 22432 4672 22438
rect 4620 22374 4672 22380
rect 4214 22332 4522 22352
rect 4214 22330 4220 22332
rect 4276 22330 4300 22332
rect 4356 22330 4380 22332
rect 4436 22330 4460 22332
rect 4516 22330 4522 22332
rect 4276 22278 4278 22330
rect 4458 22278 4460 22330
rect 4214 22276 4220 22278
rect 4276 22276 4300 22278
rect 4356 22276 4380 22278
rect 4436 22276 4460 22278
rect 4516 22276 4522 22278
rect 4214 22256 4522 22276
rect 3436 22066 3556 22094
rect 3436 17066 3464 22066
rect 4160 21888 4212 21894
rect 4160 21830 4212 21836
rect 4172 21554 4200 21830
rect 4632 21690 4660 22374
rect 4620 21684 4672 21690
rect 4620 21626 4672 21632
rect 4160 21548 4212 21554
rect 4160 21490 4212 21496
rect 4620 21548 4672 21554
rect 4620 21490 4672 21496
rect 4214 21244 4522 21264
rect 4214 21242 4220 21244
rect 4276 21242 4300 21244
rect 4356 21242 4380 21244
rect 4436 21242 4460 21244
rect 4516 21242 4522 21244
rect 4276 21190 4278 21242
rect 4458 21190 4460 21242
rect 4214 21188 4220 21190
rect 4276 21188 4300 21190
rect 4356 21188 4380 21190
rect 4436 21188 4460 21190
rect 4516 21188 4522 21190
rect 4214 21168 4522 21188
rect 4632 21010 4660 21490
rect 4620 21004 4672 21010
rect 4620 20946 4672 20952
rect 3976 20392 4028 20398
rect 3976 20334 4028 20340
rect 3988 20058 4016 20334
rect 4068 20324 4120 20330
rect 4068 20266 4120 20272
rect 3976 20052 4028 20058
rect 3976 19994 4028 20000
rect 4080 19854 4108 20266
rect 4214 20156 4522 20176
rect 4214 20154 4220 20156
rect 4276 20154 4300 20156
rect 4356 20154 4380 20156
rect 4436 20154 4460 20156
rect 4516 20154 4522 20156
rect 4276 20102 4278 20154
rect 4458 20102 4460 20154
rect 4214 20100 4220 20102
rect 4276 20100 4300 20102
rect 4356 20100 4380 20102
rect 4436 20100 4460 20102
rect 4516 20100 4522 20102
rect 4214 20080 4522 20100
rect 4068 19848 4120 19854
rect 4068 19790 4120 19796
rect 3976 19304 4028 19310
rect 3976 19246 4028 19252
rect 3988 17882 4016 19246
rect 4068 19168 4120 19174
rect 4068 19110 4120 19116
rect 4080 18970 4108 19110
rect 4214 19068 4522 19088
rect 4214 19066 4220 19068
rect 4276 19066 4300 19068
rect 4356 19066 4380 19068
rect 4436 19066 4460 19068
rect 4516 19066 4522 19068
rect 4276 19014 4278 19066
rect 4458 19014 4460 19066
rect 4214 19012 4220 19014
rect 4276 19012 4300 19014
rect 4356 19012 4380 19014
rect 4436 19012 4460 19014
rect 4516 19012 4522 19014
rect 4214 18992 4522 19012
rect 4068 18964 4120 18970
rect 4068 18906 4120 18912
rect 4080 18766 4108 18906
rect 4068 18760 4120 18766
rect 4068 18702 4120 18708
rect 4214 17980 4522 18000
rect 4214 17978 4220 17980
rect 4276 17978 4300 17980
rect 4356 17978 4380 17980
rect 4436 17978 4460 17980
rect 4516 17978 4522 17980
rect 4276 17926 4278 17978
rect 4458 17926 4460 17978
rect 4214 17924 4220 17926
rect 4276 17924 4300 17926
rect 4356 17924 4380 17926
rect 4436 17924 4460 17926
rect 4516 17924 4522 17926
rect 4214 17904 4522 17924
rect 3976 17876 4028 17882
rect 3976 17818 4028 17824
rect 3988 17746 4016 17818
rect 3976 17740 4028 17746
rect 3976 17682 4028 17688
rect 3516 17332 3568 17338
rect 3516 17274 3568 17280
rect 3424 17060 3476 17066
rect 3424 17002 3476 17008
rect 3332 16788 3384 16794
rect 3332 16730 3384 16736
rect 3436 16658 3464 17002
rect 3424 16652 3476 16658
rect 3424 16594 3476 16600
rect 3436 15026 3464 16594
rect 3528 16114 3556 17274
rect 4214 16892 4522 16912
rect 4214 16890 4220 16892
rect 4276 16890 4300 16892
rect 4356 16890 4380 16892
rect 4436 16890 4460 16892
rect 4516 16890 4522 16892
rect 4276 16838 4278 16890
rect 4458 16838 4460 16890
rect 4214 16836 4220 16838
rect 4276 16836 4300 16838
rect 4356 16836 4380 16838
rect 4436 16836 4460 16838
rect 4516 16836 4522 16838
rect 4214 16816 4522 16836
rect 4160 16584 4212 16590
rect 4160 16526 4212 16532
rect 4620 16584 4672 16590
rect 4620 16526 4672 16532
rect 4172 16250 4200 16526
rect 4160 16244 4212 16250
rect 4160 16186 4212 16192
rect 3516 16108 3568 16114
rect 3516 16050 3568 16056
rect 3792 15972 3844 15978
rect 3792 15914 3844 15920
rect 3804 15502 3832 15914
rect 4214 15804 4522 15824
rect 4214 15802 4220 15804
rect 4276 15802 4300 15804
rect 4356 15802 4380 15804
rect 4436 15802 4460 15804
rect 4516 15802 4522 15804
rect 4276 15750 4278 15802
rect 4458 15750 4460 15802
rect 4214 15748 4220 15750
rect 4276 15748 4300 15750
rect 4356 15748 4380 15750
rect 4436 15748 4460 15750
rect 4516 15748 4522 15750
rect 4214 15728 4522 15748
rect 4632 15502 4660 16526
rect 3792 15496 3844 15502
rect 3792 15438 3844 15444
rect 4620 15496 4672 15502
rect 4620 15438 4672 15444
rect 3792 15360 3844 15366
rect 3792 15302 3844 15308
rect 3804 15094 3832 15302
rect 3516 15088 3568 15094
rect 3516 15030 3568 15036
rect 3792 15088 3844 15094
rect 3792 15030 3844 15036
rect 3424 15020 3476 15026
rect 3424 14962 3476 14968
rect 3528 14346 3556 15030
rect 3884 15020 3936 15026
rect 3884 14962 3936 14968
rect 3896 14618 3924 14962
rect 4214 14716 4522 14736
rect 4214 14714 4220 14716
rect 4276 14714 4300 14716
rect 4356 14714 4380 14716
rect 4436 14714 4460 14716
rect 4516 14714 4522 14716
rect 4276 14662 4278 14714
rect 4458 14662 4460 14714
rect 4214 14660 4220 14662
rect 4276 14660 4300 14662
rect 4356 14660 4380 14662
rect 4436 14660 4460 14662
rect 4516 14660 4522 14662
rect 4214 14640 4522 14660
rect 3884 14612 3936 14618
rect 3884 14554 3936 14560
rect 3516 14340 3568 14346
rect 3516 14282 3568 14288
rect 3528 13938 3556 14282
rect 4160 14272 4212 14278
rect 4160 14214 4212 14220
rect 4172 14006 4200 14214
rect 4160 14000 4212 14006
rect 4160 13942 4212 13948
rect 3516 13932 3568 13938
rect 3516 13874 3568 13880
rect 3240 13456 3292 13462
rect 3240 13398 3292 13404
rect 3148 13320 3200 13326
rect 3148 13262 3200 13268
rect 3056 13252 3108 13258
rect 3056 13194 3108 13200
rect 3068 12918 3096 13194
rect 3056 12912 3108 12918
rect 3056 12854 3108 12860
rect 3056 12640 3108 12646
rect 3056 12582 3108 12588
rect 3068 9586 3096 12582
rect 3160 12442 3188 13262
rect 3240 12912 3292 12918
rect 3240 12854 3292 12860
rect 3148 12436 3200 12442
rect 3148 12378 3200 12384
rect 3252 11762 3280 12854
rect 3240 11756 3292 11762
rect 3240 11698 3292 11704
rect 3240 10600 3292 10606
rect 3240 10542 3292 10548
rect 3148 10056 3200 10062
rect 3148 9998 3200 10004
rect 3056 9580 3108 9586
rect 3056 9522 3108 9528
rect 3056 9444 3108 9450
rect 3056 9386 3108 9392
rect 3068 8906 3096 9386
rect 3160 8974 3188 9998
rect 3252 9178 3280 10542
rect 3424 9920 3476 9926
rect 3424 9862 3476 9868
rect 3436 9586 3464 9862
rect 3424 9580 3476 9586
rect 3424 9522 3476 9528
rect 3240 9172 3292 9178
rect 3240 9114 3292 9120
rect 3148 8968 3200 8974
rect 3148 8910 3200 8916
rect 3056 8900 3108 8906
rect 3056 8842 3108 8848
rect 2964 8628 3016 8634
rect 2964 8570 3016 8576
rect 3068 8362 3096 8842
rect 1492 8356 1544 8362
rect 1492 8298 1544 8304
rect 3056 8356 3108 8362
rect 3056 8298 3108 8304
rect 1504 8265 1532 8298
rect 1490 8256 1546 8265
rect 1490 8191 1546 8200
rect 1584 6316 1636 6322
rect 1584 6258 1636 6264
rect 1596 6225 1624 6258
rect 1582 6216 1638 6225
rect 1582 6151 1638 6160
rect 2044 6180 2096 6186
rect 1596 5914 1624 6151
rect 2044 6122 2096 6128
rect 1584 5908 1636 5914
rect 1584 5850 1636 5856
rect 1492 4480 1544 4486
rect 1492 4422 1544 4428
rect 1504 4185 1532 4422
rect 1490 4176 1546 4185
rect 1490 4111 1546 4120
rect 2056 3602 2084 6122
rect 3068 5302 3096 8298
rect 3528 6390 3556 13874
rect 4632 13802 4660 15438
rect 4712 14816 4764 14822
rect 4712 14758 4764 14764
rect 4724 14278 4752 14758
rect 4712 14272 4764 14278
rect 4712 14214 4764 14220
rect 4620 13796 4672 13802
rect 4620 13738 4672 13744
rect 4214 13628 4522 13648
rect 4214 13626 4220 13628
rect 4276 13626 4300 13628
rect 4356 13626 4380 13628
rect 4436 13626 4460 13628
rect 4516 13626 4522 13628
rect 4276 13574 4278 13626
rect 4458 13574 4460 13626
rect 4214 13572 4220 13574
rect 4276 13572 4300 13574
rect 4356 13572 4380 13574
rect 4436 13572 4460 13574
rect 4516 13572 4522 13574
rect 4214 13552 4522 13572
rect 4214 12540 4522 12560
rect 4214 12538 4220 12540
rect 4276 12538 4300 12540
rect 4356 12538 4380 12540
rect 4436 12538 4460 12540
rect 4516 12538 4522 12540
rect 4276 12486 4278 12538
rect 4458 12486 4460 12538
rect 4214 12484 4220 12486
rect 4276 12484 4300 12486
rect 4356 12484 4380 12486
rect 4436 12484 4460 12486
rect 4516 12484 4522 12486
rect 4214 12464 4522 12484
rect 4816 12434 4844 22986
rect 6196 22778 6224 23122
rect 5264 22772 5316 22778
rect 5264 22714 5316 22720
rect 6184 22772 6236 22778
rect 6184 22714 6236 22720
rect 4896 22024 4948 22030
rect 4896 21966 4948 21972
rect 5080 22024 5132 22030
rect 5080 21966 5132 21972
rect 4908 20942 4936 21966
rect 5092 21622 5120 21966
rect 5172 21684 5224 21690
rect 5172 21626 5224 21632
rect 5080 21616 5132 21622
rect 5080 21558 5132 21564
rect 5092 21010 5120 21558
rect 5080 21004 5132 21010
rect 5080 20946 5132 20952
rect 4896 20936 4948 20942
rect 4896 20878 4948 20884
rect 4896 20256 4948 20262
rect 4896 20198 4948 20204
rect 4908 18766 4936 20198
rect 4896 18760 4948 18766
rect 4896 18702 4948 18708
rect 4988 18692 5040 18698
rect 4988 18634 5040 18640
rect 5000 17678 5028 18634
rect 4988 17672 5040 17678
rect 4988 17614 5040 17620
rect 5000 17270 5028 17614
rect 4988 17264 5040 17270
rect 4988 17206 5040 17212
rect 4988 14884 5040 14890
rect 4988 14826 5040 14832
rect 4816 12406 4936 12434
rect 4252 12232 4304 12238
rect 4252 12174 4304 12180
rect 4264 11898 4292 12174
rect 4252 11892 4304 11898
rect 4252 11834 4304 11840
rect 3608 11824 3660 11830
rect 3608 11766 3660 11772
rect 3620 11354 3648 11766
rect 3792 11756 3844 11762
rect 3792 11698 3844 11704
rect 3884 11756 3936 11762
rect 3884 11698 3936 11704
rect 3700 11552 3752 11558
rect 3700 11494 3752 11500
rect 3608 11348 3660 11354
rect 3608 11290 3660 11296
rect 3712 10674 3740 11494
rect 3804 11014 3832 11698
rect 3896 11218 3924 11698
rect 4264 11642 4292 11834
rect 4080 11614 4292 11642
rect 3884 11212 3936 11218
rect 3884 11154 3936 11160
rect 3792 11008 3844 11014
rect 3792 10950 3844 10956
rect 3700 10668 3752 10674
rect 3700 10610 3752 10616
rect 3608 8968 3660 8974
rect 3608 8910 3660 8916
rect 3620 8294 3648 8910
rect 3608 8288 3660 8294
rect 3608 8230 3660 8236
rect 3712 7970 3740 10610
rect 3804 9926 3832 10950
rect 3896 10810 3924 11154
rect 4080 11150 4108 11614
rect 4214 11452 4522 11472
rect 4214 11450 4220 11452
rect 4276 11450 4300 11452
rect 4356 11450 4380 11452
rect 4436 11450 4460 11452
rect 4516 11450 4522 11452
rect 4276 11398 4278 11450
rect 4458 11398 4460 11450
rect 4214 11396 4220 11398
rect 4276 11396 4300 11398
rect 4356 11396 4380 11398
rect 4436 11396 4460 11398
rect 4516 11396 4522 11398
rect 4214 11376 4522 11396
rect 4068 11144 4120 11150
rect 4068 11086 4120 11092
rect 4068 11008 4120 11014
rect 4068 10950 4120 10956
rect 3884 10804 3936 10810
rect 3884 10746 3936 10752
rect 4080 10674 4108 10950
rect 4068 10668 4120 10674
rect 4068 10610 4120 10616
rect 4080 9994 4108 10610
rect 4214 10364 4522 10384
rect 4214 10362 4220 10364
rect 4276 10362 4300 10364
rect 4356 10362 4380 10364
rect 4436 10362 4460 10364
rect 4516 10362 4522 10364
rect 4276 10310 4278 10362
rect 4458 10310 4460 10362
rect 4214 10308 4220 10310
rect 4276 10308 4300 10310
rect 4356 10308 4380 10310
rect 4436 10308 4460 10310
rect 4516 10308 4522 10310
rect 4214 10288 4522 10308
rect 4068 9988 4120 9994
rect 4068 9930 4120 9936
rect 3792 9920 3844 9926
rect 3792 9862 3844 9868
rect 3804 9586 3832 9862
rect 3792 9580 3844 9586
rect 3792 9522 3844 9528
rect 4080 9178 4108 9930
rect 4620 9580 4672 9586
rect 4620 9522 4672 9528
rect 4214 9276 4522 9296
rect 4214 9274 4220 9276
rect 4276 9274 4300 9276
rect 4356 9274 4380 9276
rect 4436 9274 4460 9276
rect 4516 9274 4522 9276
rect 4276 9222 4278 9274
rect 4458 9222 4460 9274
rect 4214 9220 4220 9222
rect 4276 9220 4300 9222
rect 4356 9220 4380 9222
rect 4436 9220 4460 9222
rect 4516 9220 4522 9222
rect 4214 9200 4522 9220
rect 4068 9172 4120 9178
rect 4068 9114 4120 9120
rect 3792 8900 3844 8906
rect 3792 8842 3844 8848
rect 3884 8900 3936 8906
rect 3884 8842 3936 8848
rect 3804 8090 3832 8842
rect 3896 8498 3924 8842
rect 4632 8634 4660 9522
rect 4712 9376 4764 9382
rect 4712 9318 4764 9324
rect 4620 8628 4672 8634
rect 4620 8570 4672 8576
rect 3884 8492 3936 8498
rect 3884 8434 3936 8440
rect 4528 8492 4580 8498
rect 4528 8434 4580 8440
rect 3976 8424 4028 8430
rect 3976 8366 4028 8372
rect 4540 8378 4568 8434
rect 4632 8378 4660 8570
rect 3884 8288 3936 8294
rect 3884 8230 3936 8236
rect 3792 8084 3844 8090
rect 3792 8026 3844 8032
rect 3712 7942 3832 7970
rect 3516 6384 3568 6390
rect 3516 6326 3568 6332
rect 3424 6316 3476 6322
rect 3424 6258 3476 6264
rect 3436 5370 3464 6258
rect 3424 5364 3476 5370
rect 3424 5306 3476 5312
rect 3056 5296 3108 5302
rect 3056 5238 3108 5244
rect 3804 5234 3832 7942
rect 3240 5228 3292 5234
rect 3240 5170 3292 5176
rect 3792 5228 3844 5234
rect 3792 5170 3844 5176
rect 3252 4758 3280 5170
rect 3240 4752 3292 4758
rect 3240 4694 3292 4700
rect 3896 4622 3924 8230
rect 3988 8022 4016 8366
rect 4068 8356 4120 8362
rect 4540 8350 4660 8378
rect 4068 8298 4120 8304
rect 3976 8016 4028 8022
rect 3976 7958 4028 7964
rect 4080 7970 4108 8298
rect 4214 8188 4522 8208
rect 4214 8186 4220 8188
rect 4276 8186 4300 8188
rect 4356 8186 4380 8188
rect 4436 8186 4460 8188
rect 4516 8186 4522 8188
rect 4276 8134 4278 8186
rect 4458 8134 4460 8186
rect 4214 8132 4220 8134
rect 4276 8132 4300 8134
rect 4356 8132 4380 8134
rect 4436 8132 4460 8134
rect 4516 8132 4522 8134
rect 4214 8112 4522 8132
rect 4080 7942 4292 7970
rect 4264 7818 4292 7942
rect 4252 7812 4304 7818
rect 4252 7754 4304 7760
rect 4264 7342 4292 7754
rect 4252 7336 4304 7342
rect 4252 7278 4304 7284
rect 4214 7100 4522 7120
rect 4214 7098 4220 7100
rect 4276 7098 4300 7100
rect 4356 7098 4380 7100
rect 4436 7098 4460 7100
rect 4516 7098 4522 7100
rect 4276 7046 4278 7098
rect 4458 7046 4460 7098
rect 4214 7044 4220 7046
rect 4276 7044 4300 7046
rect 4356 7044 4380 7046
rect 4436 7044 4460 7046
rect 4516 7044 4522 7046
rect 4214 7024 4522 7044
rect 4214 6012 4522 6032
rect 4214 6010 4220 6012
rect 4276 6010 4300 6012
rect 4356 6010 4380 6012
rect 4436 6010 4460 6012
rect 4516 6010 4522 6012
rect 4276 5958 4278 6010
rect 4458 5958 4460 6010
rect 4214 5956 4220 5958
rect 4276 5956 4300 5958
rect 4356 5956 4380 5958
rect 4436 5956 4460 5958
rect 4516 5956 4522 5958
rect 4214 5936 4522 5956
rect 4632 5778 4660 8350
rect 4724 6390 4752 9318
rect 4712 6384 4764 6390
rect 4712 6326 4764 6332
rect 4620 5772 4672 5778
rect 4620 5714 4672 5720
rect 3976 5228 4028 5234
rect 3976 5170 4028 5176
rect 3988 4826 4016 5170
rect 4214 4924 4522 4944
rect 4214 4922 4220 4924
rect 4276 4922 4300 4924
rect 4356 4922 4380 4924
rect 4436 4922 4460 4924
rect 4516 4922 4522 4924
rect 4276 4870 4278 4922
rect 4458 4870 4460 4922
rect 4214 4868 4220 4870
rect 4276 4868 4300 4870
rect 4356 4868 4380 4870
rect 4436 4868 4460 4870
rect 4516 4868 4522 4870
rect 4214 4848 4522 4868
rect 3976 4820 4028 4826
rect 3976 4762 4028 4768
rect 3884 4616 3936 4622
rect 3884 4558 3936 4564
rect 4214 3836 4522 3856
rect 4214 3834 4220 3836
rect 4276 3834 4300 3836
rect 4356 3834 4380 3836
rect 4436 3834 4460 3836
rect 4516 3834 4522 3836
rect 4276 3782 4278 3834
rect 4458 3782 4460 3834
rect 4214 3780 4220 3782
rect 4276 3780 4300 3782
rect 4356 3780 4380 3782
rect 4436 3780 4460 3782
rect 4516 3780 4522 3782
rect 4214 3760 4522 3780
rect 2044 3596 2096 3602
rect 2044 3538 2096 3544
rect 1400 3392 1452 3398
rect 1400 3334 1452 3340
rect 1412 3058 1440 3334
rect 1400 3052 1452 3058
rect 1400 2994 1452 3000
rect 20 2848 72 2854
rect 20 2790 72 2796
rect 32 800 60 2790
rect 1412 2145 1440 2994
rect 1492 2848 1544 2854
rect 1492 2790 1544 2796
rect 2596 2848 2648 2854
rect 2596 2790 2648 2796
rect 1504 2446 1532 2790
rect 2608 2446 2636 2790
rect 4214 2748 4522 2768
rect 4214 2746 4220 2748
rect 4276 2746 4300 2748
rect 4356 2746 4380 2748
rect 4436 2746 4460 2748
rect 4516 2746 4522 2748
rect 4276 2694 4278 2746
rect 4458 2694 4460 2746
rect 4214 2692 4220 2694
rect 4276 2692 4300 2694
rect 4356 2692 4380 2694
rect 4436 2692 4460 2694
rect 4516 2692 4522 2694
rect 4214 2672 4522 2692
rect 4908 2650 4936 12406
rect 5000 3194 5028 14826
rect 4988 3188 5040 3194
rect 4988 3130 5040 3136
rect 5080 2916 5132 2922
rect 5080 2858 5132 2864
rect 4896 2644 4948 2650
rect 4896 2586 4948 2592
rect 5092 2446 5120 2858
rect 1492 2440 1544 2446
rect 1492 2382 1544 2388
rect 1952 2440 2004 2446
rect 1952 2382 2004 2388
rect 2596 2440 2648 2446
rect 2596 2382 2648 2388
rect 5080 2440 5132 2446
rect 5080 2382 5132 2388
rect 1398 2136 1454 2145
rect 1398 2071 1454 2080
rect 1964 800 1992 2382
rect 3884 2304 3936 2310
rect 3884 2246 3936 2252
rect 3896 800 3924 2246
rect 5184 2106 5212 21626
rect 5276 20602 5304 22714
rect 6840 22642 6868 23258
rect 7024 23186 7052 23598
rect 7300 23322 7328 24754
rect 7288 23316 7340 23322
rect 7288 23258 7340 23264
rect 7012 23180 7064 23186
rect 7012 23122 7064 23128
rect 6828 22636 6880 22642
rect 6828 22578 6880 22584
rect 7472 22160 7524 22166
rect 7472 22102 7524 22108
rect 7104 22024 7156 22030
rect 7104 21966 7156 21972
rect 6736 21888 6788 21894
rect 6736 21830 6788 21836
rect 6748 21554 6776 21830
rect 6736 21548 6788 21554
rect 6736 21490 6788 21496
rect 5816 21344 5868 21350
rect 5816 21286 5868 21292
rect 5828 21078 5856 21286
rect 5816 21072 5868 21078
rect 5816 21014 5868 21020
rect 6748 21010 6776 21490
rect 6736 21004 6788 21010
rect 6736 20946 6788 20952
rect 6460 20800 6512 20806
rect 6460 20742 6512 20748
rect 5264 20596 5316 20602
rect 5264 20538 5316 20544
rect 5276 19922 5304 20538
rect 6472 20466 6500 20742
rect 6460 20460 6512 20466
rect 6460 20402 6512 20408
rect 5448 20052 5500 20058
rect 5448 19994 5500 20000
rect 5264 19916 5316 19922
rect 5264 19858 5316 19864
rect 5460 19514 5488 19994
rect 6920 19984 6972 19990
rect 6920 19926 6972 19932
rect 5540 19848 5592 19854
rect 5540 19790 5592 19796
rect 5448 19508 5500 19514
rect 5448 19450 5500 19456
rect 5552 19378 5580 19790
rect 6276 19712 6328 19718
rect 6276 19654 6328 19660
rect 6288 19378 6316 19654
rect 5540 19372 5592 19378
rect 5540 19314 5592 19320
rect 6276 19372 6328 19378
rect 6276 19314 6328 19320
rect 6288 18698 6316 19314
rect 6932 19310 6960 19926
rect 7116 19854 7144 21966
rect 7484 21010 7512 22102
rect 7576 21554 7604 31146
rect 7656 30252 7708 30258
rect 7656 30194 7708 30200
rect 7668 29714 7696 30194
rect 7656 29708 7708 29714
rect 7656 29650 7708 29656
rect 7656 24336 7708 24342
rect 7656 24278 7708 24284
rect 7668 23798 7696 24278
rect 7656 23792 7708 23798
rect 7656 23734 7708 23740
rect 7748 23724 7800 23730
rect 7748 23666 7800 23672
rect 7760 23254 7788 23666
rect 7748 23248 7800 23254
rect 7748 23190 7800 23196
rect 7656 22636 7708 22642
rect 7656 22578 7708 22584
rect 7668 22030 7696 22578
rect 7656 22024 7708 22030
rect 7656 21966 7708 21972
rect 7564 21548 7616 21554
rect 7564 21490 7616 21496
rect 7472 21004 7524 21010
rect 7472 20946 7524 20952
rect 7484 20602 7512 20946
rect 7576 20942 7604 21490
rect 7564 20936 7616 20942
rect 7564 20878 7616 20884
rect 7840 20868 7892 20874
rect 7840 20810 7892 20816
rect 7472 20596 7524 20602
rect 7472 20538 7524 20544
rect 7104 19848 7156 19854
rect 7104 19790 7156 19796
rect 7484 19378 7512 20538
rect 7852 20466 7880 20810
rect 7840 20460 7892 20466
rect 7840 20402 7892 20408
rect 7852 19854 7880 20402
rect 7840 19848 7892 19854
rect 7760 19796 7840 19802
rect 7760 19790 7892 19796
rect 7760 19774 7880 19790
rect 7760 19446 7788 19774
rect 7840 19712 7892 19718
rect 7840 19654 7892 19660
rect 7748 19440 7800 19446
rect 7748 19382 7800 19388
rect 7196 19372 7248 19378
rect 7196 19314 7248 19320
rect 7472 19372 7524 19378
rect 7472 19314 7524 19320
rect 6920 19304 6972 19310
rect 6920 19246 6972 19252
rect 7208 18766 7236 19314
rect 7484 18834 7512 19314
rect 7748 19304 7800 19310
rect 7748 19246 7800 19252
rect 7656 19236 7708 19242
rect 7656 19178 7708 19184
rect 7472 18828 7524 18834
rect 7472 18770 7524 18776
rect 7196 18760 7248 18766
rect 7196 18702 7248 18708
rect 7564 18760 7616 18766
rect 7564 18702 7616 18708
rect 6276 18692 6328 18698
rect 6276 18634 6328 18640
rect 7576 18426 7604 18702
rect 7564 18420 7616 18426
rect 7564 18362 7616 18368
rect 7668 18290 7696 19178
rect 7760 18970 7788 19246
rect 7748 18964 7800 18970
rect 7748 18906 7800 18912
rect 7852 18290 7880 19654
rect 7196 18284 7248 18290
rect 7196 18226 7248 18232
rect 7656 18284 7708 18290
rect 7656 18226 7708 18232
rect 7840 18284 7892 18290
rect 7840 18226 7892 18232
rect 6000 18080 6052 18086
rect 6000 18022 6052 18028
rect 6012 17678 6040 18022
rect 7012 17876 7064 17882
rect 7012 17818 7064 17824
rect 6000 17672 6052 17678
rect 6000 17614 6052 17620
rect 7024 16794 7052 17818
rect 7208 17814 7236 18226
rect 7472 18080 7524 18086
rect 7472 18022 7524 18028
rect 7196 17808 7248 17814
rect 7196 17750 7248 17756
rect 7288 17604 7340 17610
rect 7288 17546 7340 17552
rect 7300 17134 7328 17546
rect 7484 17270 7512 18022
rect 7668 17882 7696 18226
rect 7656 17876 7708 17882
rect 7656 17818 7708 17824
rect 7748 17672 7800 17678
rect 7852 17660 7880 18226
rect 7800 17632 7880 17660
rect 7748 17614 7800 17620
rect 7472 17264 7524 17270
rect 7472 17206 7524 17212
rect 7288 17128 7340 17134
rect 7288 17070 7340 17076
rect 7012 16788 7064 16794
rect 7012 16730 7064 16736
rect 7484 16590 7512 17206
rect 7840 16992 7892 16998
rect 7840 16934 7892 16940
rect 7852 16794 7880 16934
rect 7840 16788 7892 16794
rect 7840 16730 7892 16736
rect 7472 16584 7524 16590
rect 7472 16526 7524 16532
rect 7562 16144 7618 16153
rect 7196 16108 7248 16114
rect 7562 16079 7564 16088
rect 7196 16050 7248 16056
rect 7616 16079 7618 16088
rect 7564 16050 7616 16056
rect 6920 15972 6972 15978
rect 6920 15914 6972 15920
rect 6932 15502 6960 15914
rect 6920 15496 6972 15502
rect 6920 15438 6972 15444
rect 6644 15088 6696 15094
rect 6644 15030 6696 15036
rect 5816 15020 5868 15026
rect 5816 14962 5868 14968
rect 5356 14272 5408 14278
rect 5356 14214 5408 14220
rect 5368 13870 5396 14214
rect 5356 13864 5408 13870
rect 5356 13806 5408 13812
rect 5368 7857 5396 13806
rect 5724 12164 5776 12170
rect 5724 12106 5776 12112
rect 5736 11898 5764 12106
rect 5724 11892 5776 11898
rect 5724 11834 5776 11840
rect 5354 7848 5410 7857
rect 5354 7783 5410 7792
rect 5828 2774 5856 14962
rect 6656 14346 6684 15030
rect 6932 14618 6960 15438
rect 7208 15026 7236 16050
rect 7748 15496 7800 15502
rect 7748 15438 7800 15444
rect 7760 15162 7788 15438
rect 7748 15156 7800 15162
rect 7748 15098 7800 15104
rect 7196 15020 7248 15026
rect 7196 14962 7248 14968
rect 6920 14612 6972 14618
rect 6920 14554 6972 14560
rect 6644 14340 6696 14346
rect 6644 14282 6696 14288
rect 6368 13320 6420 13326
rect 6368 13262 6420 13268
rect 6276 13252 6328 13258
rect 6276 13194 6328 13200
rect 5908 12640 5960 12646
rect 5908 12582 5960 12588
rect 5920 12442 5948 12582
rect 5908 12436 5960 12442
rect 6288 12434 6316 13194
rect 6380 12918 6408 13262
rect 6368 12912 6420 12918
rect 6368 12854 6420 12860
rect 6552 12844 6604 12850
rect 6552 12786 6604 12792
rect 6288 12406 6500 12434
rect 5908 12378 5960 12384
rect 6472 12238 6500 12406
rect 6564 12306 6592 12786
rect 6552 12300 6604 12306
rect 6552 12242 6604 12248
rect 6460 12232 6512 12238
rect 6460 12174 6512 12180
rect 6184 12164 6236 12170
rect 6184 12106 6236 12112
rect 6196 11762 6224 12106
rect 6184 11756 6236 11762
rect 6184 11698 6236 11704
rect 6368 11756 6420 11762
rect 6368 11698 6420 11704
rect 6380 10810 6408 11698
rect 6472 11626 6500 12174
rect 6460 11620 6512 11626
rect 6460 11562 6512 11568
rect 6368 10804 6420 10810
rect 6368 10746 6420 10752
rect 6000 10600 6052 10606
rect 6000 10542 6052 10548
rect 6012 10266 6040 10542
rect 6656 10538 6684 14282
rect 7380 13864 7432 13870
rect 7380 13806 7432 13812
rect 7392 13326 7420 13806
rect 7944 13530 7972 34478
rect 8208 33992 8260 33998
rect 8208 33934 8260 33940
rect 8220 33522 8248 33934
rect 8300 33924 8352 33930
rect 8300 33866 8352 33872
rect 8312 33522 8340 33866
rect 8208 33516 8260 33522
rect 8208 33458 8260 33464
rect 8300 33516 8352 33522
rect 8300 33458 8352 33464
rect 8312 33402 8340 33458
rect 8116 33380 8168 33386
rect 8116 33322 8168 33328
rect 8220 33374 8340 33402
rect 8128 32910 8156 33322
rect 8116 32904 8168 32910
rect 8116 32846 8168 32852
rect 8116 32768 8168 32774
rect 8116 32710 8168 32716
rect 8128 32434 8156 32710
rect 8116 32428 8168 32434
rect 8116 32370 8168 32376
rect 8128 31346 8156 32370
rect 8220 31822 8248 33374
rect 8392 32292 8444 32298
rect 8392 32234 8444 32240
rect 8404 32026 8432 32234
rect 8392 32020 8444 32026
rect 8392 31962 8444 31968
rect 8208 31816 8260 31822
rect 8208 31758 8260 31764
rect 8116 31340 8168 31346
rect 8116 31282 8168 31288
rect 8220 28150 8248 31758
rect 8208 28144 8260 28150
rect 8208 28086 8260 28092
rect 8484 28076 8536 28082
rect 8484 28018 8536 28024
rect 8024 27940 8076 27946
rect 8024 27882 8076 27888
rect 8036 27470 8064 27882
rect 8496 27470 8524 28018
rect 8024 27464 8076 27470
rect 8024 27406 8076 27412
rect 8484 27464 8536 27470
rect 8484 27406 8536 27412
rect 8036 27062 8064 27406
rect 8116 27328 8168 27334
rect 8116 27270 8168 27276
rect 8024 27056 8076 27062
rect 8024 26998 8076 27004
rect 8036 26518 8064 26998
rect 8128 26994 8156 27270
rect 8116 26988 8168 26994
rect 8116 26930 8168 26936
rect 8024 26512 8076 26518
rect 8024 26454 8076 26460
rect 8024 26376 8076 26382
rect 8024 26318 8076 26324
rect 8036 24818 8064 26318
rect 8300 24948 8352 24954
rect 8300 24890 8352 24896
rect 8484 24948 8536 24954
rect 8484 24890 8536 24896
rect 8208 24880 8260 24886
rect 8208 24822 8260 24828
rect 8024 24812 8076 24818
rect 8024 24754 8076 24760
rect 8220 24410 8248 24822
rect 8208 24404 8260 24410
rect 8208 24346 8260 24352
rect 8024 23520 8076 23526
rect 8024 23462 8076 23468
rect 8036 23118 8064 23462
rect 8024 23112 8076 23118
rect 8024 23054 8076 23060
rect 8036 22030 8064 23054
rect 8312 22642 8340 24890
rect 8392 24744 8444 24750
rect 8392 24686 8444 24692
rect 8404 24410 8432 24686
rect 8392 24404 8444 24410
rect 8392 24346 8444 24352
rect 8392 24200 8444 24206
rect 8390 24168 8392 24177
rect 8444 24168 8446 24177
rect 8390 24103 8446 24112
rect 8496 22778 8524 24890
rect 8484 22772 8536 22778
rect 8484 22714 8536 22720
rect 8300 22636 8352 22642
rect 8300 22578 8352 22584
rect 8024 22024 8076 22030
rect 8024 21966 8076 21972
rect 8036 21418 8064 21966
rect 8024 21412 8076 21418
rect 8024 21354 8076 21360
rect 8300 20936 8352 20942
rect 8300 20878 8352 20884
rect 8116 20868 8168 20874
rect 8116 20810 8168 20816
rect 8024 20460 8076 20466
rect 8024 20402 8076 20408
rect 8036 19786 8064 20402
rect 8128 19990 8156 20810
rect 8208 20596 8260 20602
rect 8208 20538 8260 20544
rect 8220 20058 8248 20538
rect 8208 20052 8260 20058
rect 8208 19994 8260 20000
rect 8116 19984 8168 19990
rect 8116 19926 8168 19932
rect 8024 19780 8076 19786
rect 8024 19722 8076 19728
rect 8036 19378 8064 19722
rect 8024 19372 8076 19378
rect 8024 19314 8076 19320
rect 8036 18834 8064 19314
rect 8024 18828 8076 18834
rect 8024 18770 8076 18776
rect 8024 18284 8076 18290
rect 8024 18226 8076 18232
rect 8036 17678 8064 18226
rect 8312 18086 8340 20878
rect 8300 18080 8352 18086
rect 8300 18022 8352 18028
rect 8024 17672 8076 17678
rect 8024 17614 8076 17620
rect 8208 17536 8260 17542
rect 8208 17478 8260 17484
rect 8220 17270 8248 17478
rect 8024 17264 8076 17270
rect 8208 17264 8260 17270
rect 8076 17212 8156 17218
rect 8024 17206 8156 17212
rect 8208 17206 8260 17212
rect 8036 17190 8156 17206
rect 8128 16114 8156 17190
rect 8220 17066 8248 17206
rect 8208 17060 8260 17066
rect 8208 17002 8260 17008
rect 8484 16992 8536 16998
rect 8484 16934 8536 16940
rect 8496 16590 8524 16934
rect 8484 16584 8536 16590
rect 8484 16526 8536 16532
rect 8208 16516 8260 16522
rect 8208 16458 8260 16464
rect 8220 16250 8248 16458
rect 8208 16244 8260 16250
rect 8208 16186 8260 16192
rect 8116 16108 8168 16114
rect 8116 16050 8168 16056
rect 7932 13524 7984 13530
rect 7932 13466 7984 13472
rect 7380 13320 7432 13326
rect 7380 13262 7432 13268
rect 7288 12844 7340 12850
rect 7288 12786 7340 12792
rect 7104 12232 7156 12238
rect 7104 12174 7156 12180
rect 7116 11762 7144 12174
rect 7300 12170 7328 12786
rect 7840 12640 7892 12646
rect 7840 12582 7892 12588
rect 7852 12434 7880 12582
rect 7852 12406 8064 12434
rect 8036 12238 8064 12406
rect 8024 12232 8076 12238
rect 8024 12174 8076 12180
rect 7288 12164 7340 12170
rect 7288 12106 7340 12112
rect 7300 11898 7328 12106
rect 7288 11892 7340 11898
rect 7288 11834 7340 11840
rect 7104 11756 7156 11762
rect 7104 11698 7156 11704
rect 8036 11694 8064 12174
rect 8024 11688 8076 11694
rect 7102 11656 7158 11665
rect 8024 11630 8076 11636
rect 7102 11591 7104 11600
rect 7156 11591 7158 11600
rect 7104 11562 7156 11568
rect 6828 10668 6880 10674
rect 6828 10610 6880 10616
rect 6644 10532 6696 10538
rect 6644 10474 6696 10480
rect 6840 10266 6868 10610
rect 6000 10260 6052 10266
rect 6000 10202 6052 10208
rect 6828 10260 6880 10266
rect 6828 10202 6880 10208
rect 6920 10192 6972 10198
rect 6920 10134 6972 10140
rect 6368 10124 6420 10130
rect 6368 10066 6420 10072
rect 6380 9722 6408 10066
rect 6368 9716 6420 9722
rect 6368 9658 6420 9664
rect 6932 9654 6960 10134
rect 6920 9648 6972 9654
rect 6920 9590 6972 9596
rect 6552 9512 6604 9518
rect 6552 9454 6604 9460
rect 7012 9512 7064 9518
rect 7012 9454 7064 9460
rect 6564 9178 6592 9454
rect 6552 9172 6604 9178
rect 6552 9114 6604 9120
rect 6460 8968 6512 8974
rect 6920 8968 6972 8974
rect 6512 8916 6592 8922
rect 6460 8910 6592 8916
rect 6920 8910 6972 8916
rect 6472 8894 6592 8910
rect 6564 8498 6592 8894
rect 6552 8492 6604 8498
rect 6552 8434 6604 8440
rect 6564 8090 6592 8434
rect 6932 8430 6960 8910
rect 7024 8498 7052 9454
rect 7012 8492 7064 8498
rect 7012 8434 7064 8440
rect 6920 8424 6972 8430
rect 6920 8366 6972 8372
rect 7656 8424 7708 8430
rect 7656 8366 7708 8372
rect 7668 8090 7696 8366
rect 6552 8084 6604 8090
rect 6552 8026 6604 8032
rect 7656 8084 7708 8090
rect 7656 8026 7708 8032
rect 6736 7404 6788 7410
rect 6736 7346 6788 7352
rect 6748 6934 6776 7346
rect 6828 7336 6880 7342
rect 6828 7278 6880 7284
rect 6736 6928 6788 6934
rect 6736 6870 6788 6876
rect 6748 5778 6776 6870
rect 6840 6458 6868 7278
rect 6828 6452 6880 6458
rect 6828 6394 6880 6400
rect 6840 5846 6868 6394
rect 7196 6112 7248 6118
rect 7196 6054 7248 6060
rect 6828 5840 6880 5846
rect 6828 5782 6880 5788
rect 7208 5778 7236 6054
rect 6736 5772 6788 5778
rect 6736 5714 6788 5720
rect 7196 5772 7248 5778
rect 7196 5714 7248 5720
rect 6736 5636 6788 5642
rect 6736 5578 6788 5584
rect 6748 5302 6776 5578
rect 6828 5568 6880 5574
rect 6828 5510 6880 5516
rect 6736 5296 6788 5302
rect 6736 5238 6788 5244
rect 6460 5228 6512 5234
rect 6460 5170 6512 5176
rect 6276 5024 6328 5030
rect 6276 4966 6328 4972
rect 6288 4690 6316 4966
rect 6276 4684 6328 4690
rect 6276 4626 6328 4632
rect 6288 4214 6316 4626
rect 6472 4622 6500 5170
rect 6644 5160 6696 5166
rect 6644 5102 6696 5108
rect 6656 4826 6684 5102
rect 6840 5098 6868 5510
rect 7288 5228 7340 5234
rect 7288 5170 7340 5176
rect 6828 5092 6880 5098
rect 6828 5034 6880 5040
rect 7300 4826 7328 5170
rect 6644 4820 6696 4826
rect 6644 4762 6696 4768
rect 7104 4820 7156 4826
rect 7104 4762 7156 4768
rect 7288 4820 7340 4826
rect 7288 4762 7340 4768
rect 6460 4616 6512 4622
rect 6460 4558 6512 4564
rect 6736 4616 6788 4622
rect 7116 4604 7144 4762
rect 7380 4684 7432 4690
rect 7380 4626 7432 4632
rect 7288 4616 7340 4622
rect 7116 4576 7288 4604
rect 6736 4558 6788 4564
rect 7288 4558 7340 4564
rect 6472 4282 6500 4558
rect 6460 4276 6512 4282
rect 6460 4218 6512 4224
rect 6748 4214 6776 4558
rect 6276 4208 6328 4214
rect 6276 4150 6328 4156
rect 6736 4208 6788 4214
rect 6736 4150 6788 4156
rect 7392 2922 7420 4626
rect 7380 2916 7432 2922
rect 7380 2858 7432 2864
rect 5736 2746 5856 2774
rect 5736 2514 5764 2746
rect 8128 2514 8156 16050
rect 8208 10056 8260 10062
rect 8208 9998 8260 10004
rect 8220 9178 8248 9998
rect 8588 9602 8616 36246
rect 8852 36168 8904 36174
rect 8852 36110 8904 36116
rect 8760 36032 8812 36038
rect 8760 35974 8812 35980
rect 8772 35698 8800 35974
rect 8760 35692 8812 35698
rect 8760 35634 8812 35640
rect 8864 35630 8892 36110
rect 8956 35698 8984 36314
rect 9586 35728 9642 35737
rect 8944 35692 8996 35698
rect 9586 35663 9642 35672
rect 8944 35634 8996 35640
rect 8852 35624 8904 35630
rect 8852 35566 8904 35572
rect 8864 35494 8892 35566
rect 8852 35488 8904 35494
rect 8852 35430 8904 35436
rect 8760 32020 8812 32026
rect 8760 31962 8812 31968
rect 8668 24812 8720 24818
rect 8668 24754 8720 24760
rect 8680 24614 8708 24754
rect 8668 24608 8720 24614
rect 8668 24550 8720 24556
rect 8772 22710 8800 31962
rect 8760 22704 8812 22710
rect 8760 22646 8812 22652
rect 8668 18624 8720 18630
rect 8668 18566 8720 18572
rect 8680 16250 8708 18566
rect 8668 16244 8720 16250
rect 8668 16186 8720 16192
rect 8668 12844 8720 12850
rect 8668 12786 8720 12792
rect 8680 12442 8708 12786
rect 8668 12436 8720 12442
rect 8668 12378 8720 12384
rect 8588 9574 8708 9602
rect 8208 9172 8260 9178
rect 8208 9114 8260 9120
rect 8576 9036 8628 9042
rect 8576 8978 8628 8984
rect 8588 8634 8616 8978
rect 8576 8628 8628 8634
rect 8576 8570 8628 8576
rect 8680 6769 8708 9574
rect 8666 6760 8722 6769
rect 8666 6695 8722 6704
rect 8484 2848 8536 2854
rect 8484 2790 8536 2796
rect 5724 2508 5776 2514
rect 5724 2450 5776 2456
rect 8116 2508 8168 2514
rect 8116 2450 8168 2456
rect 8496 2446 8524 2790
rect 8772 2582 8800 22646
rect 8864 13802 8892 35430
rect 9600 35290 9628 35663
rect 9588 35284 9640 35290
rect 9588 35226 9640 35232
rect 11532 35086 11560 37062
rect 14200 36854 14228 37266
rect 16500 37210 16528 39222
rect 18050 39200 18106 40000
rect 19982 39200 20038 40000
rect 21914 39200 21970 40000
rect 23846 39200 23902 40000
rect 25778 39200 25834 40000
rect 28354 39200 28410 40000
rect 30286 39200 30342 40000
rect 32218 39200 32274 40000
rect 34150 39200 34206 40000
rect 36082 39200 36138 40000
rect 38014 39200 38070 40000
rect 39946 39200 40002 40000
rect 41878 39200 41934 40000
rect 44454 39200 44510 40000
rect 46386 39200 46442 40000
rect 46492 39222 46888 39250
rect 16672 37256 16724 37262
rect 16500 37182 16620 37210
rect 16672 37198 16724 37204
rect 16592 37126 16620 37182
rect 16580 37120 16632 37126
rect 16580 37062 16632 37068
rect 14188 36848 14240 36854
rect 14188 36790 14240 36796
rect 16580 35828 16632 35834
rect 16580 35770 16632 35776
rect 11704 35692 11756 35698
rect 11704 35634 11756 35640
rect 11888 35692 11940 35698
rect 11888 35634 11940 35640
rect 11520 35080 11572 35086
rect 11520 35022 11572 35028
rect 11532 34610 11560 35022
rect 9496 34604 9548 34610
rect 9496 34546 9548 34552
rect 11520 34604 11572 34610
rect 11520 34546 11572 34552
rect 9128 33992 9180 33998
rect 9128 33934 9180 33940
rect 9140 33590 9168 33934
rect 9508 33930 9536 34546
rect 11612 34536 11664 34542
rect 11612 34478 11664 34484
rect 11152 34468 11204 34474
rect 11152 34410 11204 34416
rect 11164 33998 11192 34410
rect 11624 33998 11652 34478
rect 11716 34202 11744 35634
rect 11900 35290 11928 35634
rect 12348 35556 12400 35562
rect 12348 35498 12400 35504
rect 11888 35284 11940 35290
rect 11888 35226 11940 35232
rect 11704 34196 11756 34202
rect 11704 34138 11756 34144
rect 11796 34128 11848 34134
rect 11796 34070 11848 34076
rect 9772 33992 9824 33998
rect 9772 33934 9824 33940
rect 11152 33992 11204 33998
rect 11152 33934 11204 33940
rect 11612 33992 11664 33998
rect 11612 33934 11664 33940
rect 9496 33924 9548 33930
rect 9496 33866 9548 33872
rect 9128 33584 9180 33590
rect 9128 33526 9180 33532
rect 9784 33522 9812 33934
rect 9772 33516 9824 33522
rect 9772 33458 9824 33464
rect 8944 33448 8996 33454
rect 8944 33390 8996 33396
rect 8956 33114 8984 33390
rect 8944 33108 8996 33114
rect 8944 33050 8996 33056
rect 8956 32502 8984 33050
rect 8944 32496 8996 32502
rect 8944 32438 8996 32444
rect 9312 32496 9364 32502
rect 9312 32438 9364 32444
rect 9324 32026 9352 32438
rect 9312 32020 9364 32026
rect 9312 31962 9364 31968
rect 9784 31890 9812 33458
rect 11164 32910 11192 33934
rect 11808 33658 11836 34070
rect 11900 34066 11928 35226
rect 12164 35080 12216 35086
rect 12164 35022 12216 35028
rect 12176 34134 12204 35022
rect 12360 34610 12388 35498
rect 12440 35488 12492 35494
rect 12440 35430 12492 35436
rect 12452 35154 12480 35430
rect 16592 35290 16620 35770
rect 16580 35284 16632 35290
rect 16580 35226 16632 35232
rect 12440 35148 12492 35154
rect 12440 35090 12492 35096
rect 12452 34678 12480 35090
rect 12716 35080 12768 35086
rect 12716 35022 12768 35028
rect 12532 34944 12584 34950
rect 12532 34886 12584 34892
rect 12440 34672 12492 34678
rect 12440 34614 12492 34620
rect 12544 34610 12572 34886
rect 12348 34604 12400 34610
rect 12348 34546 12400 34552
rect 12532 34604 12584 34610
rect 12532 34546 12584 34552
rect 12164 34128 12216 34134
rect 12164 34070 12216 34076
rect 11888 34060 11940 34066
rect 11888 34002 11940 34008
rect 12072 34060 12124 34066
rect 12072 34002 12124 34008
rect 11796 33652 11848 33658
rect 11796 33594 11848 33600
rect 12084 33590 12112 34002
rect 12728 33930 12756 35022
rect 16592 35018 16620 35226
rect 12900 35012 12952 35018
rect 12900 34954 12952 34960
rect 16580 35012 16632 35018
rect 16580 34954 16632 34960
rect 12912 33998 12940 34954
rect 15292 34672 15344 34678
rect 15292 34614 15344 34620
rect 16488 34672 16540 34678
rect 16488 34614 16540 34620
rect 15200 34536 15252 34542
rect 15200 34478 15252 34484
rect 14096 34400 14148 34406
rect 14096 34342 14148 34348
rect 12900 33992 12952 33998
rect 12900 33934 12952 33940
rect 12716 33924 12768 33930
rect 12716 33866 12768 33872
rect 13728 33924 13780 33930
rect 13728 33866 13780 33872
rect 12072 33584 12124 33590
rect 12072 33526 12124 33532
rect 11612 33516 11664 33522
rect 11612 33458 11664 33464
rect 11624 32910 11652 33458
rect 12164 33448 12216 33454
rect 12164 33390 12216 33396
rect 12176 32910 12204 33390
rect 11152 32904 11204 32910
rect 11152 32846 11204 32852
rect 11612 32904 11664 32910
rect 11612 32846 11664 32852
rect 11980 32904 12032 32910
rect 11980 32846 12032 32852
rect 12164 32904 12216 32910
rect 12164 32846 12216 32852
rect 10876 32836 10928 32842
rect 10876 32778 10928 32784
rect 10416 32428 10468 32434
rect 10416 32370 10468 32376
rect 10232 32360 10284 32366
rect 10232 32302 10284 32308
rect 10048 32020 10100 32026
rect 10048 31962 10100 31968
rect 9772 31884 9824 31890
rect 9772 31826 9824 31832
rect 9956 31884 10008 31890
rect 9956 31826 10008 31832
rect 8944 31680 8996 31686
rect 8944 31622 8996 31628
rect 8956 31414 8984 31622
rect 8944 31408 8996 31414
rect 8944 31350 8996 31356
rect 9496 31272 9548 31278
rect 9496 31214 9548 31220
rect 9508 30326 9536 31214
rect 9496 30320 9548 30326
rect 9496 30262 9548 30268
rect 9128 30184 9180 30190
rect 9128 30126 9180 30132
rect 9140 29238 9168 30126
rect 9680 29844 9732 29850
rect 9680 29786 9732 29792
rect 9692 29646 9720 29786
rect 9680 29640 9732 29646
rect 9680 29582 9732 29588
rect 9128 29232 9180 29238
rect 9128 29174 9180 29180
rect 8944 29164 8996 29170
rect 8944 29106 8996 29112
rect 8956 28558 8984 29106
rect 9140 28558 9168 29174
rect 9692 28558 9720 29582
rect 9784 29102 9812 31826
rect 9864 31136 9916 31142
rect 9864 31078 9916 31084
rect 9876 30734 9904 31078
rect 9864 30728 9916 30734
rect 9864 30670 9916 30676
rect 9876 29850 9904 30670
rect 9864 29844 9916 29850
rect 9864 29786 9916 29792
rect 9864 29504 9916 29510
rect 9864 29446 9916 29452
rect 9772 29096 9824 29102
rect 9772 29038 9824 29044
rect 9876 29034 9904 29446
rect 9864 29028 9916 29034
rect 9864 28970 9916 28976
rect 9876 28694 9904 28970
rect 9864 28688 9916 28694
rect 9864 28630 9916 28636
rect 8944 28552 8996 28558
rect 8944 28494 8996 28500
rect 9128 28552 9180 28558
rect 9128 28494 9180 28500
rect 9680 28552 9732 28558
rect 9680 28494 9732 28500
rect 8956 28014 8984 28494
rect 9692 28082 9720 28494
rect 9680 28076 9732 28082
rect 9680 28018 9732 28024
rect 8944 28008 8996 28014
rect 8944 27950 8996 27956
rect 8944 27464 8996 27470
rect 8944 27406 8996 27412
rect 8956 27334 8984 27406
rect 8944 27328 8996 27334
rect 8944 27270 8996 27276
rect 8956 24177 8984 27270
rect 9772 26988 9824 26994
rect 9772 26930 9824 26936
rect 9784 25906 9812 26930
rect 9864 26784 9916 26790
rect 9864 26726 9916 26732
rect 9876 26382 9904 26726
rect 9864 26376 9916 26382
rect 9864 26318 9916 26324
rect 9404 25900 9456 25906
rect 9404 25842 9456 25848
rect 9772 25900 9824 25906
rect 9772 25842 9824 25848
rect 9416 25702 9444 25842
rect 9680 25832 9732 25838
rect 9680 25774 9732 25780
rect 9404 25696 9456 25702
rect 9404 25638 9456 25644
rect 9416 25362 9444 25638
rect 9404 25356 9456 25362
rect 9404 25298 9456 25304
rect 9220 24200 9272 24206
rect 8942 24168 8998 24177
rect 9220 24142 9272 24148
rect 8942 24103 8998 24112
rect 9232 23594 9260 24142
rect 9312 24132 9364 24138
rect 9312 24074 9364 24080
rect 9324 23730 9352 24074
rect 9416 23866 9444 25298
rect 9692 24818 9720 25774
rect 9876 25498 9904 26318
rect 9968 26042 9996 31826
rect 10060 31822 10088 31962
rect 10048 31816 10100 31822
rect 10048 31758 10100 31764
rect 10140 31816 10192 31822
rect 10140 31758 10192 31764
rect 10060 31482 10088 31758
rect 10048 31476 10100 31482
rect 10048 31418 10100 31424
rect 10048 31340 10100 31346
rect 10048 31282 10100 31288
rect 10060 30598 10088 31282
rect 10152 30938 10180 31758
rect 10140 30932 10192 30938
rect 10140 30874 10192 30880
rect 10048 30592 10100 30598
rect 10048 30534 10100 30540
rect 10060 30326 10088 30534
rect 10048 30320 10100 30326
rect 10048 30262 10100 30268
rect 10244 29458 10272 32302
rect 10428 32026 10456 32370
rect 10692 32360 10744 32366
rect 10692 32302 10744 32308
rect 10508 32224 10560 32230
rect 10508 32166 10560 32172
rect 10416 32020 10468 32026
rect 10416 31962 10468 31968
rect 10520 31822 10548 32166
rect 10704 31890 10732 32302
rect 10692 31884 10744 31890
rect 10692 31826 10744 31832
rect 10508 31816 10560 31822
rect 10508 31758 10560 31764
rect 10600 31272 10652 31278
rect 10600 31214 10652 31220
rect 10324 31136 10376 31142
rect 10324 31078 10376 31084
rect 10336 30870 10364 31078
rect 10324 30864 10376 30870
rect 10324 30806 10376 30812
rect 10336 30394 10364 30806
rect 10612 30802 10640 31214
rect 10600 30796 10652 30802
rect 10600 30738 10652 30744
rect 10324 30388 10376 30394
rect 10324 30330 10376 30336
rect 10784 30388 10836 30394
rect 10784 30330 10836 30336
rect 10692 30252 10744 30258
rect 10692 30194 10744 30200
rect 10508 30048 10560 30054
rect 10508 29990 10560 29996
rect 10152 29430 10272 29458
rect 10152 27130 10180 29430
rect 10520 29238 10548 29990
rect 10704 29850 10732 30194
rect 10796 29850 10824 30330
rect 10692 29844 10744 29850
rect 10692 29786 10744 29792
rect 10784 29844 10836 29850
rect 10784 29786 10836 29792
rect 10508 29232 10560 29238
rect 10508 29174 10560 29180
rect 10600 29164 10652 29170
rect 10600 29106 10652 29112
rect 10416 29028 10468 29034
rect 10416 28970 10468 28976
rect 10428 28150 10456 28970
rect 10612 28762 10640 29106
rect 10600 28756 10652 28762
rect 10600 28698 10652 28704
rect 10704 28694 10732 29786
rect 10782 29064 10838 29073
rect 10782 28999 10838 29008
rect 10796 28762 10824 28999
rect 10784 28756 10836 28762
rect 10784 28698 10836 28704
rect 10692 28688 10744 28694
rect 10692 28630 10744 28636
rect 10508 28484 10560 28490
rect 10508 28426 10560 28432
rect 10692 28484 10744 28490
rect 10692 28426 10744 28432
rect 10416 28144 10468 28150
rect 10416 28086 10468 28092
rect 10520 27946 10548 28426
rect 10508 27940 10560 27946
rect 10508 27882 10560 27888
rect 10140 27124 10192 27130
rect 10140 27066 10192 27072
rect 10048 27056 10100 27062
rect 10048 26998 10100 27004
rect 9956 26036 10008 26042
rect 9956 25978 10008 25984
rect 9864 25492 9916 25498
rect 9864 25434 9916 25440
rect 9680 24812 9732 24818
rect 9680 24754 9732 24760
rect 9876 24698 9904 25434
rect 10060 25226 10088 26998
rect 10324 26784 10376 26790
rect 10324 26726 10376 26732
rect 10336 26382 10364 26726
rect 10140 26376 10192 26382
rect 10140 26318 10192 26324
rect 10324 26376 10376 26382
rect 10324 26318 10376 26324
rect 10152 25770 10180 26318
rect 10232 26240 10284 26246
rect 10232 26182 10284 26188
rect 10244 25906 10272 26182
rect 10232 25900 10284 25906
rect 10232 25842 10284 25848
rect 10324 25832 10376 25838
rect 10324 25774 10376 25780
rect 10140 25764 10192 25770
rect 10140 25706 10192 25712
rect 10336 25498 10364 25774
rect 10324 25492 10376 25498
rect 10324 25434 10376 25440
rect 10048 25220 10100 25226
rect 10048 25162 10100 25168
rect 10060 24818 10088 25162
rect 10048 24812 10100 24818
rect 9784 24670 9904 24698
rect 9968 24772 10048 24800
rect 9680 24608 9732 24614
rect 9680 24550 9732 24556
rect 9404 23860 9456 23866
rect 9404 23802 9456 23808
rect 9312 23724 9364 23730
rect 9312 23666 9364 23672
rect 9220 23588 9272 23594
rect 9220 23530 9272 23536
rect 9324 23322 9352 23666
rect 9312 23316 9364 23322
rect 9312 23258 9364 23264
rect 9416 22030 9444 23802
rect 9496 23316 9548 23322
rect 9496 23258 9548 23264
rect 9404 22024 9456 22030
rect 9404 21966 9456 21972
rect 9312 21888 9364 21894
rect 9312 21830 9364 21836
rect 9324 20942 9352 21830
rect 9508 21622 9536 23258
rect 9692 21622 9720 24550
rect 9784 24138 9812 24670
rect 9772 24132 9824 24138
rect 9772 24074 9824 24080
rect 9968 23798 9996 24772
rect 10048 24754 10100 24760
rect 10324 24200 10376 24206
rect 10324 24142 10376 24148
rect 10336 23866 10364 24142
rect 10324 23860 10376 23866
rect 10324 23802 10376 23808
rect 9956 23792 10008 23798
rect 9956 23734 10008 23740
rect 10140 23724 10192 23730
rect 10520 23712 10548 27882
rect 10704 27402 10732 28426
rect 10692 27396 10744 27402
rect 10692 27338 10744 27344
rect 10704 26042 10732 27338
rect 10600 26036 10652 26042
rect 10600 25978 10652 25984
rect 10692 26036 10744 26042
rect 10692 25978 10744 25984
rect 10612 25906 10640 25978
rect 10600 25900 10652 25906
rect 10600 25842 10652 25848
rect 10140 23666 10192 23672
rect 10336 23684 10548 23712
rect 10152 23118 10180 23666
rect 9864 23112 9916 23118
rect 9864 23054 9916 23060
rect 10140 23112 10192 23118
rect 10140 23054 10192 23060
rect 9876 22710 9904 23054
rect 9864 22704 9916 22710
rect 9864 22646 9916 22652
rect 9772 22432 9824 22438
rect 9772 22374 9824 22380
rect 9496 21616 9548 21622
rect 9496 21558 9548 21564
rect 9680 21616 9732 21622
rect 9784 21593 9812 22374
rect 9876 22098 9904 22646
rect 9864 22092 9916 22098
rect 9864 22034 9916 22040
rect 9680 21558 9732 21564
rect 9770 21584 9826 21593
rect 9508 21146 9536 21558
rect 9876 21554 9904 22034
rect 9956 22024 10008 22030
rect 9956 21966 10008 21972
rect 10048 22024 10100 22030
rect 10048 21966 10100 21972
rect 9968 21690 9996 21966
rect 10060 21894 10088 21966
rect 10048 21888 10100 21894
rect 10048 21830 10100 21836
rect 9956 21684 10008 21690
rect 9956 21626 10008 21632
rect 9770 21519 9772 21528
rect 9824 21519 9826 21528
rect 9864 21548 9916 21554
rect 9772 21490 9824 21496
rect 9864 21490 9916 21496
rect 9784 21146 9812 21490
rect 9496 21140 9548 21146
rect 9496 21082 9548 21088
rect 9772 21140 9824 21146
rect 9772 21082 9824 21088
rect 9312 20936 9364 20942
rect 9312 20878 9364 20884
rect 10336 20466 10364 23684
rect 10612 23526 10640 25842
rect 10704 25226 10732 25978
rect 10692 25220 10744 25226
rect 10692 25162 10744 25168
rect 10784 24676 10836 24682
rect 10784 24618 10836 24624
rect 10796 24138 10824 24618
rect 10888 24410 10916 32778
rect 10968 30388 11020 30394
rect 10968 30330 11020 30336
rect 10980 26586 11008 30330
rect 11060 30048 11112 30054
rect 11058 30016 11060 30025
rect 11112 30016 11114 30025
rect 11058 29951 11114 29960
rect 11072 29782 11100 29951
rect 11060 29776 11112 29782
rect 11060 29718 11112 29724
rect 11164 29170 11192 32846
rect 11244 30660 11296 30666
rect 11244 30602 11296 30608
rect 11152 29164 11204 29170
rect 11152 29106 11204 29112
rect 11164 28558 11192 29106
rect 11152 28552 11204 28558
rect 11152 28494 11204 28500
rect 11256 27538 11284 30602
rect 11992 28966 12020 32846
rect 13740 32774 13768 33866
rect 13268 32768 13320 32774
rect 13268 32710 13320 32716
rect 13728 32768 13780 32774
rect 13728 32710 13780 32716
rect 13280 32434 13308 32710
rect 13740 32434 13768 32710
rect 13268 32428 13320 32434
rect 13268 32370 13320 32376
rect 13728 32428 13780 32434
rect 13728 32370 13780 32376
rect 13544 31816 13596 31822
rect 13544 31758 13596 31764
rect 13360 31748 13412 31754
rect 13360 31690 13412 31696
rect 13176 31680 13228 31686
rect 13176 31622 13228 31628
rect 13188 31142 13216 31622
rect 13372 31414 13400 31690
rect 13556 31414 13584 31758
rect 13360 31408 13412 31414
rect 13360 31350 13412 31356
rect 13544 31408 13596 31414
rect 13544 31350 13596 31356
rect 13176 31136 13228 31142
rect 13176 31078 13228 31084
rect 12900 30932 12952 30938
rect 12900 30874 12952 30880
rect 12716 30796 12768 30802
rect 12716 30738 12768 30744
rect 12728 30598 12756 30738
rect 12716 30592 12768 30598
rect 12716 30534 12768 30540
rect 12912 30258 12940 30874
rect 12992 30728 13044 30734
rect 12992 30670 13044 30676
rect 13084 30728 13136 30734
rect 13084 30670 13136 30676
rect 13004 30258 13032 30670
rect 13096 30598 13124 30670
rect 13084 30592 13136 30598
rect 13084 30534 13136 30540
rect 13188 30326 13216 31078
rect 13372 30870 13400 31350
rect 13360 30864 13412 30870
rect 13360 30806 13412 30812
rect 13268 30796 13320 30802
rect 13268 30738 13320 30744
rect 13176 30320 13228 30326
rect 13176 30262 13228 30268
rect 12900 30252 12952 30258
rect 12900 30194 12952 30200
rect 12992 30252 13044 30258
rect 12992 30194 13044 30200
rect 12440 30184 12492 30190
rect 12440 30126 12492 30132
rect 12452 29646 12480 30126
rect 13004 29850 13032 30194
rect 13280 30190 13308 30738
rect 13556 30598 13584 31350
rect 13544 30592 13596 30598
rect 13544 30534 13596 30540
rect 13268 30184 13320 30190
rect 13268 30126 13320 30132
rect 13820 30116 13872 30122
rect 13820 30058 13872 30064
rect 12992 29844 13044 29850
rect 12992 29786 13044 29792
rect 12440 29640 12492 29646
rect 12440 29582 12492 29588
rect 13636 29640 13688 29646
rect 13636 29582 13688 29588
rect 12624 29572 12676 29578
rect 12624 29514 12676 29520
rect 12256 29504 12308 29510
rect 12256 29446 12308 29452
rect 12348 29504 12400 29510
rect 12348 29446 12400 29452
rect 11980 28960 12032 28966
rect 11980 28902 12032 28908
rect 11992 28626 12020 28902
rect 12164 28756 12216 28762
rect 12164 28698 12216 28704
rect 11980 28620 12032 28626
rect 11980 28562 12032 28568
rect 12176 28558 12204 28698
rect 11428 28552 11480 28558
rect 11428 28494 11480 28500
rect 12164 28552 12216 28558
rect 12164 28494 12216 28500
rect 11244 27532 11296 27538
rect 11244 27474 11296 27480
rect 11440 26994 11468 28494
rect 12268 27878 12296 29446
rect 12360 28762 12388 29446
rect 12636 29306 12664 29514
rect 13082 29336 13138 29345
rect 12624 29300 12676 29306
rect 13082 29271 13084 29280
rect 12624 29242 12676 29248
rect 13136 29271 13138 29280
rect 13452 29300 13504 29306
rect 13084 29242 13136 29248
rect 13452 29242 13504 29248
rect 12348 28756 12400 28762
rect 12348 28698 12400 28704
rect 12256 27872 12308 27878
rect 12256 27814 12308 27820
rect 11796 27464 11848 27470
rect 11796 27406 11848 27412
rect 11428 26988 11480 26994
rect 11428 26930 11480 26936
rect 10968 26580 11020 26586
rect 10968 26522 11020 26528
rect 11440 26314 11468 26930
rect 11244 26308 11296 26314
rect 11244 26250 11296 26256
rect 11428 26308 11480 26314
rect 11428 26250 11480 26256
rect 11256 25974 11284 26250
rect 11244 25968 11296 25974
rect 11244 25910 11296 25916
rect 11808 25906 11836 27406
rect 12268 27062 12296 27814
rect 13096 27470 13124 29242
rect 13464 28558 13492 29242
rect 13648 29209 13676 29582
rect 13728 29504 13780 29510
rect 13728 29446 13780 29452
rect 13634 29200 13690 29209
rect 13634 29135 13690 29144
rect 13648 29034 13676 29135
rect 13740 29034 13768 29446
rect 13636 29028 13688 29034
rect 13636 28970 13688 28976
rect 13728 29028 13780 29034
rect 13728 28970 13780 28976
rect 13452 28552 13504 28558
rect 13452 28494 13504 28500
rect 13268 27600 13320 27606
rect 13268 27542 13320 27548
rect 13084 27464 13136 27470
rect 13084 27406 13136 27412
rect 13280 27062 13308 27542
rect 12256 27056 12308 27062
rect 12256 26998 12308 27004
rect 13268 27056 13320 27062
rect 13268 26998 13320 27004
rect 11888 26852 11940 26858
rect 11888 26794 11940 26800
rect 11900 26450 11928 26794
rect 11888 26444 11940 26450
rect 11888 26386 11940 26392
rect 12992 25968 13044 25974
rect 12992 25910 13044 25916
rect 11796 25900 11848 25906
rect 11796 25842 11848 25848
rect 11060 25696 11112 25702
rect 11060 25638 11112 25644
rect 10876 24404 10928 24410
rect 10876 24346 10928 24352
rect 10784 24132 10836 24138
rect 10784 24074 10836 24080
rect 10796 23866 10824 24074
rect 10784 23860 10836 23866
rect 10784 23802 10836 23808
rect 10600 23520 10652 23526
rect 10796 23497 10824 23802
rect 10600 23462 10652 23468
rect 10782 23488 10838 23497
rect 10612 22642 10640 23462
rect 10782 23423 10838 23432
rect 10600 22636 10652 22642
rect 10600 22578 10652 22584
rect 10612 22234 10640 22578
rect 10600 22228 10652 22234
rect 10600 22170 10652 22176
rect 10796 22094 10824 23423
rect 10876 22094 10928 22098
rect 10796 22092 10928 22094
rect 10796 22066 10876 22092
rect 10876 22034 10928 22040
rect 11072 22030 11100 25638
rect 13004 25294 13032 25910
rect 13280 25906 13308 26998
rect 13544 26920 13596 26926
rect 13544 26862 13596 26868
rect 13556 26586 13584 26862
rect 13544 26580 13596 26586
rect 13544 26522 13596 26528
rect 13648 25906 13676 28970
rect 13728 28552 13780 28558
rect 13728 28494 13780 28500
rect 13740 28218 13768 28494
rect 13832 28218 13860 30058
rect 14108 29510 14136 34342
rect 15212 34202 15240 34478
rect 15200 34196 15252 34202
rect 15200 34138 15252 34144
rect 15304 33998 15332 34614
rect 15844 34604 15896 34610
rect 15844 34546 15896 34552
rect 15856 33998 15884 34546
rect 16120 34536 16172 34542
rect 16120 34478 16172 34484
rect 16132 34134 16160 34478
rect 16120 34128 16172 34134
rect 16120 34070 16172 34076
rect 14188 33992 14240 33998
rect 14188 33934 14240 33940
rect 15292 33992 15344 33998
rect 15292 33934 15344 33940
rect 15844 33992 15896 33998
rect 15844 33934 15896 33940
rect 14200 31958 14228 33934
rect 15856 32502 15884 33934
rect 15844 32496 15896 32502
rect 15844 32438 15896 32444
rect 15200 32428 15252 32434
rect 15200 32370 15252 32376
rect 15660 32428 15712 32434
rect 15660 32370 15712 32376
rect 15108 32360 15160 32366
rect 15108 32302 15160 32308
rect 14280 32224 14332 32230
rect 14280 32166 14332 32172
rect 14464 32224 14516 32230
rect 14464 32166 14516 32172
rect 14292 31958 14320 32166
rect 14188 31952 14240 31958
rect 14188 31894 14240 31900
rect 14280 31952 14332 31958
rect 14280 31894 14332 31900
rect 14372 30728 14424 30734
rect 14372 30670 14424 30676
rect 14188 29572 14240 29578
rect 14188 29514 14240 29520
rect 14096 29504 14148 29510
rect 14096 29446 14148 29452
rect 13910 29336 13966 29345
rect 14108 29306 14136 29446
rect 13910 29271 13966 29280
rect 14096 29300 14148 29306
rect 13924 29170 13952 29271
rect 14096 29242 14148 29248
rect 13912 29164 13964 29170
rect 13912 29106 13964 29112
rect 14002 29064 14058 29073
rect 14200 29034 14228 29514
rect 14002 28999 14058 29008
rect 14188 29028 14240 29034
rect 13728 28212 13780 28218
rect 13728 28154 13780 28160
rect 13820 28212 13872 28218
rect 13820 28154 13872 28160
rect 14016 28082 14044 28999
rect 14188 28970 14240 28976
rect 14004 28076 14056 28082
rect 14004 28018 14056 28024
rect 13728 28008 13780 28014
rect 13728 27950 13780 27956
rect 13740 26976 13768 27950
rect 14384 27606 14412 30670
rect 14476 29850 14504 32166
rect 15120 31482 15148 32302
rect 15212 32026 15240 32370
rect 15292 32292 15344 32298
rect 15292 32234 15344 32240
rect 15200 32020 15252 32026
rect 15200 31962 15252 31968
rect 15108 31476 15160 31482
rect 15108 31418 15160 31424
rect 14556 30728 14608 30734
rect 14556 30670 14608 30676
rect 14568 30190 14596 30670
rect 14556 30184 14608 30190
rect 14556 30126 14608 30132
rect 14464 29844 14516 29850
rect 14464 29786 14516 29792
rect 15108 29844 15160 29850
rect 15108 29786 15160 29792
rect 15120 29646 15148 29786
rect 15016 29640 15068 29646
rect 15016 29582 15068 29588
rect 15108 29640 15160 29646
rect 15108 29582 15160 29588
rect 14922 29200 14978 29209
rect 14648 29164 14700 29170
rect 14648 29106 14700 29112
rect 14740 29164 14792 29170
rect 14922 29135 14924 29144
rect 14740 29106 14792 29112
rect 14976 29135 14978 29144
rect 14924 29106 14976 29112
rect 14660 29073 14688 29106
rect 14646 29064 14702 29073
rect 14646 28999 14702 29008
rect 14556 28416 14608 28422
rect 14556 28358 14608 28364
rect 14464 27940 14516 27946
rect 14464 27882 14516 27888
rect 14372 27600 14424 27606
rect 14372 27542 14424 27548
rect 14476 27470 14504 27882
rect 14280 27464 14332 27470
rect 14280 27406 14332 27412
rect 14464 27464 14516 27470
rect 14464 27406 14516 27412
rect 13820 26988 13872 26994
rect 13740 26948 13820 26976
rect 13268 25900 13320 25906
rect 13268 25842 13320 25848
rect 13636 25900 13688 25906
rect 13636 25842 13688 25848
rect 13176 25832 13228 25838
rect 13176 25774 13228 25780
rect 13084 25764 13136 25770
rect 13084 25706 13136 25712
rect 12440 25288 12492 25294
rect 12440 25230 12492 25236
rect 12992 25288 13044 25294
rect 12992 25230 13044 25236
rect 11980 24880 12032 24886
rect 11980 24822 12032 24828
rect 11520 22976 11572 22982
rect 11520 22918 11572 22924
rect 10784 22024 10836 22030
rect 10784 21966 10836 21972
rect 11060 22024 11112 22030
rect 11060 21966 11112 21972
rect 10508 21888 10560 21894
rect 10508 21830 10560 21836
rect 10520 21457 10548 21830
rect 10506 21448 10562 21457
rect 10506 21383 10562 21392
rect 10796 20942 10824 21966
rect 11244 21888 11296 21894
rect 11244 21830 11296 21836
rect 11256 21486 11284 21830
rect 11532 21690 11560 22918
rect 11520 21684 11572 21690
rect 11520 21626 11572 21632
rect 11060 21480 11112 21486
rect 11060 21422 11112 21428
rect 11244 21480 11296 21486
rect 11244 21422 11296 21428
rect 11072 21321 11100 21422
rect 11058 21312 11114 21321
rect 11058 21247 11114 21256
rect 10784 20936 10836 20942
rect 10784 20878 10836 20884
rect 10416 20528 10468 20534
rect 10414 20496 10416 20505
rect 10468 20496 10470 20505
rect 9496 20460 9548 20466
rect 9496 20402 9548 20408
rect 9956 20460 10008 20466
rect 9956 20402 10008 20408
rect 10324 20460 10376 20466
rect 10414 20431 10470 20440
rect 10324 20402 10376 20408
rect 9508 19786 9536 20402
rect 9680 20324 9732 20330
rect 9680 20266 9732 20272
rect 9692 19854 9720 20266
rect 9680 19848 9732 19854
rect 9680 19790 9732 19796
rect 9496 19780 9548 19786
rect 9496 19722 9548 19728
rect 9968 19446 9996 20402
rect 11152 20256 11204 20262
rect 11152 20198 11204 20204
rect 11164 19922 11192 20198
rect 11992 19922 12020 24822
rect 12452 23730 12480 25230
rect 12716 25152 12768 25158
rect 12716 25094 12768 25100
rect 12440 23724 12492 23730
rect 12440 23666 12492 23672
rect 12532 23656 12584 23662
rect 12532 23598 12584 23604
rect 12544 23526 12572 23598
rect 12532 23520 12584 23526
rect 12532 23462 12584 23468
rect 12728 23338 12756 25094
rect 12808 24404 12860 24410
rect 12808 24346 12860 24352
rect 12820 23866 12848 24346
rect 12992 24200 13044 24206
rect 12992 24142 13044 24148
rect 12808 23860 12860 23866
rect 12808 23802 12860 23808
rect 13004 23594 13032 24142
rect 12992 23588 13044 23594
rect 12992 23530 13044 23536
rect 12728 23310 12848 23338
rect 12820 23254 12848 23310
rect 12808 23248 12860 23254
rect 12808 23190 12860 23196
rect 12624 23112 12676 23118
rect 12624 23054 12676 23060
rect 12636 20618 12664 23054
rect 12820 22642 12848 23190
rect 12900 22704 12952 22710
rect 12900 22646 12952 22652
rect 12808 22636 12860 22642
rect 12808 22578 12860 22584
rect 12912 22166 12940 22646
rect 12992 22636 13044 22642
rect 12992 22578 13044 22584
rect 12900 22160 12952 22166
rect 12900 22102 12952 22108
rect 12912 21554 12940 22102
rect 13004 21876 13032 22578
rect 13096 22574 13124 25706
rect 13188 25226 13216 25774
rect 13176 25220 13228 25226
rect 13176 25162 13228 25168
rect 13084 22568 13136 22574
rect 13084 22510 13136 22516
rect 13096 22234 13124 22510
rect 13084 22228 13136 22234
rect 13084 22170 13136 22176
rect 13188 22030 13216 25162
rect 13280 24070 13308 25842
rect 13648 25362 13676 25842
rect 13740 25838 13768 26948
rect 13820 26930 13872 26936
rect 14292 26926 14320 27406
rect 14568 26994 14596 28358
rect 14648 27124 14700 27130
rect 14648 27066 14700 27072
rect 14464 26988 14516 26994
rect 14464 26930 14516 26936
rect 14556 26988 14608 26994
rect 14556 26930 14608 26936
rect 14280 26920 14332 26926
rect 14280 26862 14332 26868
rect 14096 26580 14148 26586
rect 14096 26522 14148 26528
rect 13728 25832 13780 25838
rect 13728 25774 13780 25780
rect 14108 25770 14136 26522
rect 14476 26042 14504 26930
rect 14464 26036 14516 26042
rect 14464 25978 14516 25984
rect 14096 25764 14148 25770
rect 14096 25706 14148 25712
rect 14568 25430 14596 26930
rect 14660 26926 14688 27066
rect 14648 26920 14700 26926
rect 14648 26862 14700 26868
rect 14556 25424 14608 25430
rect 14556 25366 14608 25372
rect 13636 25356 13688 25362
rect 13636 25298 13688 25304
rect 14004 25356 14056 25362
rect 14004 25298 14056 25304
rect 13544 24812 13596 24818
rect 13544 24754 13596 24760
rect 13360 24744 13412 24750
rect 13360 24686 13412 24692
rect 13372 24342 13400 24686
rect 13360 24336 13412 24342
rect 13360 24278 13412 24284
rect 13556 24138 13584 24754
rect 13544 24132 13596 24138
rect 13544 24074 13596 24080
rect 13268 24064 13320 24070
rect 13268 24006 13320 24012
rect 13556 23662 13584 24074
rect 13820 24064 13872 24070
rect 13820 24006 13872 24012
rect 13636 23724 13688 23730
rect 13636 23666 13688 23672
rect 13544 23656 13596 23662
rect 13544 23598 13596 23604
rect 13648 23118 13676 23666
rect 13832 23254 13860 24006
rect 13820 23248 13872 23254
rect 13820 23190 13872 23196
rect 13636 23112 13688 23118
rect 13636 23054 13688 23060
rect 13728 22976 13780 22982
rect 13728 22918 13780 22924
rect 13740 22234 13768 22918
rect 14016 22642 14044 25298
rect 14464 25220 14516 25226
rect 14464 25162 14516 25168
rect 14096 25152 14148 25158
rect 14096 25094 14148 25100
rect 14108 24614 14136 25094
rect 14188 24676 14240 24682
rect 14188 24618 14240 24624
rect 14096 24608 14148 24614
rect 14096 24550 14148 24556
rect 14108 24070 14136 24550
rect 14200 24206 14228 24618
rect 14476 24206 14504 25162
rect 14660 24274 14688 26862
rect 14752 25906 14780 29106
rect 15028 28558 15056 29582
rect 15016 28552 15068 28558
rect 15016 28494 15068 28500
rect 15108 28144 15160 28150
rect 15108 28086 15160 28092
rect 15120 27130 15148 28086
rect 15200 28076 15252 28082
rect 15200 28018 15252 28024
rect 15212 27878 15240 28018
rect 15200 27872 15252 27878
rect 15200 27814 15252 27820
rect 15304 27606 15332 32234
rect 15672 32026 15700 32370
rect 16212 32292 16264 32298
rect 16212 32234 16264 32240
rect 15660 32020 15712 32026
rect 15660 31962 15712 31968
rect 16224 31822 16252 32234
rect 16500 32230 16528 34614
rect 16580 32904 16632 32910
rect 16580 32846 16632 32852
rect 16488 32224 16540 32230
rect 16488 32166 16540 32172
rect 16500 32026 16528 32166
rect 16592 32026 16620 32846
rect 16488 32020 16540 32026
rect 16488 31962 16540 31968
rect 16580 32020 16632 32026
rect 16580 31962 16632 31968
rect 16212 31816 16264 31822
rect 16212 31758 16264 31764
rect 15844 30728 15896 30734
rect 15896 30688 15976 30716
rect 15844 30670 15896 30676
rect 15948 30258 15976 30688
rect 16028 30320 16080 30326
rect 16028 30262 16080 30268
rect 15568 30252 15620 30258
rect 15568 30194 15620 30200
rect 15844 30252 15896 30258
rect 15844 30194 15896 30200
rect 15936 30252 15988 30258
rect 15936 30194 15988 30200
rect 15384 30048 15436 30054
rect 15384 29990 15436 29996
rect 15396 29850 15424 29990
rect 15384 29844 15436 29850
rect 15384 29786 15436 29792
rect 15476 29504 15528 29510
rect 15476 29446 15528 29452
rect 15488 29170 15516 29446
rect 15580 29306 15608 30194
rect 15856 30138 15884 30194
rect 16040 30138 16068 30262
rect 15856 30110 16068 30138
rect 15856 29850 15884 30110
rect 15844 29844 15896 29850
rect 15844 29786 15896 29792
rect 16028 29640 16080 29646
rect 16028 29582 16080 29588
rect 16212 29640 16264 29646
rect 16212 29582 16264 29588
rect 16040 29345 16068 29582
rect 16026 29336 16082 29345
rect 15568 29300 15620 29306
rect 16026 29271 16082 29280
rect 15568 29242 15620 29248
rect 15476 29164 15528 29170
rect 15476 29106 15528 29112
rect 15292 27600 15344 27606
rect 15292 27542 15344 27548
rect 15108 27124 15160 27130
rect 15108 27066 15160 27072
rect 14924 26988 14976 26994
rect 14924 26930 14976 26936
rect 14740 25900 14792 25906
rect 14740 25842 14792 25848
rect 14936 25294 14964 26930
rect 15304 26926 15332 27542
rect 15488 27130 15516 29106
rect 15658 27432 15714 27441
rect 15658 27367 15714 27376
rect 15476 27124 15528 27130
rect 15476 27066 15528 27072
rect 15292 26920 15344 26926
rect 15292 26862 15344 26868
rect 15016 26852 15068 26858
rect 15016 26794 15068 26800
rect 15028 26450 15056 26794
rect 15200 26512 15252 26518
rect 15200 26454 15252 26460
rect 15016 26444 15068 26450
rect 15016 26386 15068 26392
rect 14924 25288 14976 25294
rect 14738 25256 14794 25265
rect 14924 25230 14976 25236
rect 14738 25191 14794 25200
rect 14752 25158 14780 25191
rect 14740 25152 14792 25158
rect 14740 25094 14792 25100
rect 14740 24336 14792 24342
rect 14738 24304 14740 24313
rect 14792 24304 14794 24313
rect 14648 24268 14700 24274
rect 14738 24239 14794 24248
rect 14648 24210 14700 24216
rect 14188 24200 14240 24206
rect 14188 24142 14240 24148
rect 14464 24200 14516 24206
rect 14464 24142 14516 24148
rect 14556 24200 14608 24206
rect 14556 24142 14608 24148
rect 14200 24070 14228 24142
rect 14096 24064 14148 24070
rect 14096 24006 14148 24012
rect 14188 24064 14240 24070
rect 14188 24006 14240 24012
rect 14108 23526 14136 24006
rect 14568 23866 14596 24142
rect 14556 23860 14608 23866
rect 14556 23802 14608 23808
rect 14568 23730 14596 23802
rect 14556 23724 14608 23730
rect 14556 23666 14608 23672
rect 14096 23520 14148 23526
rect 14096 23462 14148 23468
rect 14004 22636 14056 22642
rect 13832 22596 14004 22624
rect 13360 22228 13412 22234
rect 13360 22170 13412 22176
rect 13728 22228 13780 22234
rect 13728 22170 13780 22176
rect 13176 22024 13228 22030
rect 13176 21966 13228 21972
rect 13176 21888 13228 21894
rect 13004 21848 13176 21876
rect 13176 21830 13228 21836
rect 13188 21554 13216 21830
rect 13372 21554 13400 22170
rect 13544 22024 13596 22030
rect 13544 21966 13596 21972
rect 13556 21690 13584 21966
rect 13544 21684 13596 21690
rect 13544 21626 13596 21632
rect 12900 21548 12952 21554
rect 12900 21490 12952 21496
rect 13176 21548 13228 21554
rect 13176 21490 13228 21496
rect 13360 21548 13412 21554
rect 13360 21490 13412 21496
rect 12992 21412 13044 21418
rect 12992 21354 13044 21360
rect 13004 20874 13032 21354
rect 13188 20874 13216 21490
rect 13372 21146 13400 21490
rect 13360 21140 13412 21146
rect 13360 21082 13412 21088
rect 13832 21010 13860 22596
rect 14004 22578 14056 22584
rect 14108 21321 14136 23462
rect 14464 22976 14516 22982
rect 14464 22918 14516 22924
rect 14476 22710 14504 22918
rect 14464 22704 14516 22710
rect 14464 22646 14516 22652
rect 14936 22642 14964 25230
rect 15028 24614 15056 26386
rect 15212 26314 15240 26454
rect 15200 26308 15252 26314
rect 15200 26250 15252 26256
rect 15212 25974 15240 26250
rect 15200 25968 15252 25974
rect 15200 25910 15252 25916
rect 15672 24954 15700 27367
rect 16040 27062 16068 29271
rect 16224 29073 16252 29582
rect 16210 29064 16266 29073
rect 16210 28999 16266 29008
rect 16224 28082 16252 28999
rect 16212 28076 16264 28082
rect 16212 28018 16264 28024
rect 16028 27056 16080 27062
rect 16028 26998 16080 27004
rect 16488 26988 16540 26994
rect 16488 26930 16540 26936
rect 15660 24948 15712 24954
rect 15660 24890 15712 24896
rect 15198 24848 15254 24857
rect 15198 24783 15200 24792
rect 15252 24783 15254 24792
rect 15200 24754 15252 24760
rect 15016 24608 15068 24614
rect 15016 24550 15068 24556
rect 15106 23488 15162 23497
rect 15106 23423 15162 23432
rect 15016 23180 15068 23186
rect 15016 23122 15068 23128
rect 15028 22642 15056 23122
rect 14188 22636 14240 22642
rect 14188 22578 14240 22584
rect 14924 22636 14976 22642
rect 14924 22578 14976 22584
rect 15016 22636 15068 22642
rect 15016 22578 15068 22584
rect 14200 22409 14228 22578
rect 14462 22536 14518 22545
rect 14280 22500 14332 22506
rect 14462 22471 14464 22480
rect 14280 22442 14332 22448
rect 14516 22471 14518 22480
rect 14464 22442 14516 22448
rect 14186 22400 14242 22409
rect 14186 22335 14242 22344
rect 14200 21622 14228 22335
rect 14292 22098 14320 22442
rect 14936 22098 14964 22578
rect 15120 22506 15148 23423
rect 15476 23316 15528 23322
rect 15476 23258 15528 23264
rect 15384 23112 15436 23118
rect 15384 23054 15436 23060
rect 15396 22778 15424 23054
rect 15384 22772 15436 22778
rect 15384 22714 15436 22720
rect 15198 22672 15254 22681
rect 15198 22607 15254 22616
rect 15108 22500 15160 22506
rect 15108 22442 15160 22448
rect 14280 22094 14332 22098
rect 14280 22092 14596 22094
rect 14332 22066 14596 22092
rect 14280 22034 14332 22040
rect 14188 21616 14240 21622
rect 14188 21558 14240 21564
rect 14094 21312 14150 21321
rect 14150 21270 14320 21298
rect 14094 21247 14150 21256
rect 13820 21004 13872 21010
rect 13820 20946 13872 20952
rect 13728 20936 13780 20942
rect 13728 20878 13780 20884
rect 12992 20868 13044 20874
rect 12992 20810 13044 20816
rect 13176 20868 13228 20874
rect 13176 20810 13228 20816
rect 12636 20590 12756 20618
rect 12624 20460 12676 20466
rect 12624 20402 12676 20408
rect 11152 19916 11204 19922
rect 11152 19858 11204 19864
rect 11980 19916 12032 19922
rect 11980 19858 12032 19864
rect 10232 19780 10284 19786
rect 10232 19722 10284 19728
rect 9956 19440 10008 19446
rect 9956 19382 10008 19388
rect 9956 18216 10008 18222
rect 9956 18158 10008 18164
rect 8944 17536 8996 17542
rect 8944 17478 8996 17484
rect 8956 17338 8984 17478
rect 8944 17332 8996 17338
rect 8944 17274 8996 17280
rect 9128 17332 9180 17338
rect 9128 17274 9180 17280
rect 9036 17128 9088 17134
rect 9036 17070 9088 17076
rect 9048 16794 9076 17070
rect 9036 16788 9088 16794
rect 9036 16730 9088 16736
rect 9140 16726 9168 17274
rect 9968 17202 9996 18158
rect 9956 17196 10008 17202
rect 9956 17138 10008 17144
rect 10140 17196 10192 17202
rect 10140 17138 10192 17144
rect 9968 16810 9996 17138
rect 10152 16998 10180 17138
rect 10140 16992 10192 16998
rect 10140 16934 10192 16940
rect 9968 16794 10088 16810
rect 9968 16788 10100 16794
rect 9968 16782 10048 16788
rect 10048 16730 10100 16736
rect 9128 16720 9180 16726
rect 9128 16662 9180 16668
rect 9956 16720 10008 16726
rect 9956 16662 10008 16668
rect 9036 16584 9088 16590
rect 9036 16526 9088 16532
rect 9680 16584 9732 16590
rect 9680 16526 9732 16532
rect 9048 16114 9076 16526
rect 9220 16516 9272 16522
rect 9220 16458 9272 16464
rect 9312 16516 9364 16522
rect 9312 16458 9364 16464
rect 9232 16114 9260 16458
rect 9324 16250 9352 16458
rect 9312 16244 9364 16250
rect 9312 16186 9364 16192
rect 9588 16244 9640 16250
rect 9588 16186 9640 16192
rect 9036 16108 9088 16114
rect 9036 16050 9088 16056
rect 9220 16108 9272 16114
rect 9220 16050 9272 16056
rect 9048 15706 9076 16050
rect 9036 15700 9088 15706
rect 9036 15642 9088 15648
rect 9232 15570 9260 16050
rect 9220 15564 9272 15570
rect 9220 15506 9272 15512
rect 8944 15360 8996 15366
rect 8944 15302 8996 15308
rect 8956 14890 8984 15302
rect 9232 15162 9260 15506
rect 9600 15450 9628 16186
rect 9692 15638 9720 16526
rect 9968 16114 9996 16662
rect 10152 16522 10180 16934
rect 10140 16516 10192 16522
rect 10140 16458 10192 16464
rect 9956 16108 10008 16114
rect 9956 16050 10008 16056
rect 10048 16040 10100 16046
rect 10048 15982 10100 15988
rect 9680 15632 9732 15638
rect 9680 15574 9732 15580
rect 10060 15502 10088 15982
rect 9680 15496 9732 15502
rect 9600 15444 9680 15450
rect 9600 15438 9732 15444
rect 10048 15496 10100 15502
rect 10048 15438 10100 15444
rect 9600 15422 9720 15438
rect 9220 15156 9272 15162
rect 9220 15098 9272 15104
rect 10060 15094 10088 15438
rect 10048 15088 10100 15094
rect 10048 15030 10100 15036
rect 8944 14884 8996 14890
rect 8944 14826 8996 14832
rect 8956 14482 8984 14826
rect 10060 14618 10088 15030
rect 10140 15020 10192 15026
rect 10140 14962 10192 14968
rect 10048 14612 10100 14618
rect 10048 14554 10100 14560
rect 10152 14498 10180 14962
rect 10244 14634 10272 19722
rect 11164 19310 11192 19858
rect 11152 19304 11204 19310
rect 11152 19246 11204 19252
rect 10508 19236 10560 19242
rect 10508 19178 10560 19184
rect 10520 18902 10548 19178
rect 11164 18986 11192 19246
rect 11072 18970 11192 18986
rect 11060 18964 11192 18970
rect 11112 18958 11192 18964
rect 11060 18906 11112 18912
rect 10508 18896 10560 18902
rect 10508 18838 10560 18844
rect 11072 18766 11100 18906
rect 11060 18760 11112 18766
rect 11060 18702 11112 18708
rect 10692 18284 10744 18290
rect 10692 18226 10744 18232
rect 10416 17264 10468 17270
rect 10416 17206 10468 17212
rect 10428 16522 10456 17206
rect 10416 16516 10468 16522
rect 10416 16458 10468 16464
rect 10600 16448 10652 16454
rect 10600 16390 10652 16396
rect 10508 15972 10560 15978
rect 10508 15914 10560 15920
rect 10416 15428 10468 15434
rect 10416 15370 10468 15376
rect 10428 14890 10456 15370
rect 10416 14884 10468 14890
rect 10416 14826 10468 14832
rect 10244 14606 10456 14634
rect 8944 14476 8996 14482
rect 10152 14470 10364 14498
rect 8944 14418 8996 14424
rect 10336 14414 10364 14470
rect 10324 14408 10376 14414
rect 10324 14350 10376 14356
rect 9680 13932 9732 13938
rect 9680 13874 9732 13880
rect 8852 13796 8904 13802
rect 8852 13738 8904 13744
rect 9692 13530 9720 13874
rect 9680 13524 9732 13530
rect 9680 13466 9732 13472
rect 9864 13456 9916 13462
rect 9864 13398 9916 13404
rect 9680 13184 9732 13190
rect 9680 13126 9732 13132
rect 9692 12918 9720 13126
rect 9680 12912 9732 12918
rect 9680 12854 9732 12860
rect 8852 12844 8904 12850
rect 8852 12786 8904 12792
rect 8864 12306 8892 12786
rect 8852 12300 8904 12306
rect 8852 12242 8904 12248
rect 9876 12238 9904 13398
rect 8944 12232 8996 12238
rect 8944 12174 8996 12180
rect 9864 12232 9916 12238
rect 9864 12174 9916 12180
rect 8956 11898 8984 12174
rect 9680 12164 9732 12170
rect 9680 12106 9732 12112
rect 8944 11892 8996 11898
rect 8944 11834 8996 11840
rect 9692 11830 9720 12106
rect 9680 11824 9732 11830
rect 9680 11766 9732 11772
rect 9312 11756 9364 11762
rect 9312 11698 9364 11704
rect 9324 10810 9352 11698
rect 9876 11558 9904 12174
rect 10232 12096 10284 12102
rect 10232 12038 10284 12044
rect 10048 11824 10100 11830
rect 10048 11766 10100 11772
rect 9864 11552 9916 11558
rect 9864 11494 9916 11500
rect 9312 10804 9364 10810
rect 9312 10746 9364 10752
rect 9496 10600 9548 10606
rect 9496 10542 9548 10548
rect 9508 10266 9536 10542
rect 9496 10260 9548 10266
rect 9496 10202 9548 10208
rect 8852 10124 8904 10130
rect 8852 10066 8904 10072
rect 8864 9586 8892 10066
rect 9876 10033 9904 11494
rect 10060 10810 10088 11766
rect 10244 11694 10272 12038
rect 10232 11688 10284 11694
rect 10232 11630 10284 11636
rect 10140 11008 10192 11014
rect 10140 10950 10192 10956
rect 10048 10804 10100 10810
rect 10048 10746 10100 10752
rect 10152 10674 10180 10950
rect 10140 10668 10192 10674
rect 10140 10610 10192 10616
rect 10244 10169 10272 11630
rect 10230 10160 10286 10169
rect 10230 10095 10286 10104
rect 9862 10024 9918 10033
rect 9862 9959 9918 9968
rect 9588 9920 9640 9926
rect 9588 9862 9640 9868
rect 9600 9654 9628 9862
rect 9588 9648 9640 9654
rect 9588 9590 9640 9596
rect 8852 9580 8904 9586
rect 8852 9522 8904 9528
rect 8864 9178 8892 9522
rect 9600 9489 9628 9590
rect 9586 9480 9642 9489
rect 9586 9415 9642 9424
rect 8852 9172 8904 9178
rect 8852 9114 8904 9120
rect 10048 9036 10100 9042
rect 10048 8978 10100 8984
rect 10060 8945 10088 8978
rect 10046 8936 10102 8945
rect 10046 8871 10048 8880
rect 10100 8871 10102 8880
rect 10048 8842 10100 8848
rect 9588 7812 9640 7818
rect 9588 7754 9640 7760
rect 9600 7002 9628 7754
rect 9588 6996 9640 7002
rect 9588 6938 9640 6944
rect 10048 6860 10100 6866
rect 10048 6802 10100 6808
rect 10060 6322 10088 6802
rect 10140 6724 10192 6730
rect 10140 6666 10192 6672
rect 10152 6322 10180 6666
rect 10232 6384 10284 6390
rect 10232 6326 10284 6332
rect 10048 6316 10100 6322
rect 10048 6258 10100 6264
rect 10140 6316 10192 6322
rect 10140 6258 10192 6264
rect 9680 6112 9732 6118
rect 9680 6054 9732 6060
rect 9692 5370 9720 6054
rect 10060 5914 10088 6258
rect 10048 5908 10100 5914
rect 10048 5850 10100 5856
rect 9680 5364 9732 5370
rect 9680 5306 9732 5312
rect 10048 5228 10100 5234
rect 10048 5170 10100 5176
rect 9680 5092 9732 5098
rect 9680 5034 9732 5040
rect 9692 4146 9720 5034
rect 9680 4140 9732 4146
rect 9680 4082 9732 4088
rect 9692 2922 9720 4082
rect 9772 4072 9824 4078
rect 9772 4014 9824 4020
rect 9784 3738 9812 4014
rect 10060 3738 10088 5170
rect 10244 4690 10272 6326
rect 10336 5522 10364 14350
rect 10428 12374 10456 14606
rect 10520 12434 10548 15914
rect 10612 15638 10640 16390
rect 10600 15632 10652 15638
rect 10600 15574 10652 15580
rect 10704 15450 10732 18226
rect 11888 16720 11940 16726
rect 11888 16662 11940 16668
rect 11900 16153 11928 16662
rect 11886 16144 11942 16153
rect 10968 16108 11020 16114
rect 11886 16079 11942 16088
rect 10968 16050 11020 16056
rect 10612 15422 10732 15450
rect 10784 15496 10836 15502
rect 10784 15438 10836 15444
rect 10612 14822 10640 15422
rect 10692 15360 10744 15366
rect 10692 15302 10744 15308
rect 10704 15026 10732 15302
rect 10692 15020 10744 15026
rect 10692 14962 10744 14968
rect 10600 14816 10652 14822
rect 10600 14758 10652 14764
rect 10796 14618 10824 15438
rect 10980 14822 11008 16050
rect 11336 15972 11388 15978
rect 11336 15914 11388 15920
rect 11348 15570 11376 15914
rect 11336 15564 11388 15570
rect 11336 15506 11388 15512
rect 11888 15020 11940 15026
rect 11888 14962 11940 14968
rect 11900 14906 11928 14962
rect 11808 14878 11928 14906
rect 11808 14822 11836 14878
rect 10968 14816 11020 14822
rect 10968 14758 11020 14764
rect 11796 14816 11848 14822
rect 11796 14758 11848 14764
rect 10784 14612 10836 14618
rect 10784 14554 10836 14560
rect 10968 13864 11020 13870
rect 10968 13806 11020 13812
rect 10876 13184 10928 13190
rect 10876 13126 10928 13132
rect 10888 12646 10916 13126
rect 10980 12986 11008 13806
rect 10968 12980 11020 12986
rect 10968 12922 11020 12928
rect 10876 12640 10928 12646
rect 10980 12617 11008 12922
rect 11992 12850 12020 19858
rect 12636 17882 12664 20402
rect 12624 17876 12676 17882
rect 12624 17818 12676 17824
rect 12440 17740 12492 17746
rect 12440 17682 12492 17688
rect 12452 17134 12480 17682
rect 12636 17678 12664 17818
rect 12624 17672 12676 17678
rect 12624 17614 12676 17620
rect 12440 17128 12492 17134
rect 12440 17070 12492 17076
rect 12440 16516 12492 16522
rect 12440 16458 12492 16464
rect 12452 16182 12480 16458
rect 12440 16176 12492 16182
rect 12440 16118 12492 16124
rect 12348 15156 12400 15162
rect 12348 15098 12400 15104
rect 12072 15088 12124 15094
rect 12072 15030 12124 15036
rect 12084 14793 12112 15030
rect 12360 15008 12388 15098
rect 12440 15020 12492 15026
rect 12360 14980 12440 15008
rect 12070 14784 12126 14793
rect 12070 14719 12126 14728
rect 12360 14618 12388 14980
rect 12440 14962 12492 14968
rect 12624 15020 12676 15026
rect 12624 14962 12676 14968
rect 12532 14884 12584 14890
rect 12532 14826 12584 14832
rect 12348 14612 12400 14618
rect 12348 14554 12400 14560
rect 12544 14006 12572 14826
rect 12636 14793 12664 14962
rect 12622 14784 12678 14793
rect 12622 14719 12678 14728
rect 12532 14000 12584 14006
rect 12532 13942 12584 13948
rect 12348 13456 12400 13462
rect 12348 13398 12400 13404
rect 11980 12844 12032 12850
rect 11980 12786 12032 12792
rect 10876 12582 10928 12588
rect 10966 12608 11022 12617
rect 10520 12406 10640 12434
rect 10416 12368 10468 12374
rect 10416 12310 10468 12316
rect 10612 9110 10640 12406
rect 10888 10713 10916 12582
rect 10966 12543 11022 12552
rect 11888 12096 11940 12102
rect 11888 12038 11940 12044
rect 11900 11762 11928 12038
rect 12360 11762 12388 13398
rect 12728 12850 12756 20590
rect 13004 20058 13032 20810
rect 13740 20466 13768 20878
rect 13832 20534 13860 20946
rect 13820 20528 13872 20534
rect 13820 20470 13872 20476
rect 13360 20460 13412 20466
rect 13360 20402 13412 20408
rect 13728 20460 13780 20466
rect 13728 20402 13780 20408
rect 13082 20360 13138 20369
rect 13082 20295 13084 20304
rect 13136 20295 13138 20304
rect 13084 20266 13136 20272
rect 12992 20052 13044 20058
rect 12992 19994 13044 20000
rect 12992 19168 13044 19174
rect 12992 19110 13044 19116
rect 12808 18624 12860 18630
rect 12808 18566 12860 18572
rect 12820 18290 12848 18566
rect 12808 18284 12860 18290
rect 12808 18226 12860 18232
rect 12820 18086 12848 18226
rect 13004 18154 13032 19110
rect 12992 18148 13044 18154
rect 12992 18090 13044 18096
rect 12808 18080 12860 18086
rect 12808 18022 12860 18028
rect 12716 12844 12768 12850
rect 12716 12786 12768 12792
rect 12440 12776 12492 12782
rect 12440 12718 12492 12724
rect 12452 12306 12480 12718
rect 12440 12300 12492 12306
rect 12440 12242 12492 12248
rect 12624 11824 12676 11830
rect 12624 11766 12676 11772
rect 11888 11756 11940 11762
rect 11888 11698 11940 11704
rect 12348 11756 12400 11762
rect 12348 11698 12400 11704
rect 11900 11218 11928 11698
rect 11888 11212 11940 11218
rect 11888 11154 11940 11160
rect 12360 11150 12388 11698
rect 12348 11144 12400 11150
rect 12348 11086 12400 11092
rect 12348 11008 12400 11014
rect 12348 10950 12400 10956
rect 10874 10704 10930 10713
rect 12360 10674 12388 10950
rect 10874 10639 10930 10648
rect 12164 10668 12216 10674
rect 12164 10610 12216 10616
rect 12348 10668 12400 10674
rect 12348 10610 12400 10616
rect 10692 10600 10744 10606
rect 10690 10568 10692 10577
rect 10744 10568 10746 10577
rect 10690 10503 10746 10512
rect 11520 10464 11572 10470
rect 11520 10406 11572 10412
rect 11532 9586 11560 10406
rect 12176 10266 12204 10610
rect 12440 10464 12492 10470
rect 12440 10406 12492 10412
rect 12164 10260 12216 10266
rect 12164 10202 12216 10208
rect 12452 9586 12480 10406
rect 12636 10130 12664 11766
rect 12624 10124 12676 10130
rect 12624 10066 12676 10072
rect 12636 9586 12664 10066
rect 11520 9580 11572 9586
rect 11520 9522 11572 9528
rect 12440 9580 12492 9586
rect 12440 9522 12492 9528
rect 12624 9580 12676 9586
rect 12624 9522 12676 9528
rect 10876 9376 10928 9382
rect 10876 9318 10928 9324
rect 10600 9104 10652 9110
rect 10600 9046 10652 9052
rect 10888 8974 10916 9318
rect 10968 9036 11020 9042
rect 10968 8978 11020 8984
rect 10876 8968 10928 8974
rect 10876 8910 10928 8916
rect 10888 8090 10916 8910
rect 10876 8084 10928 8090
rect 10876 8026 10928 8032
rect 10980 7954 11008 8978
rect 12440 8288 12492 8294
rect 12440 8230 12492 8236
rect 10968 7948 11020 7954
rect 10968 7890 11020 7896
rect 10416 7812 10468 7818
rect 10416 7754 10468 7760
rect 10428 7410 10456 7754
rect 10508 7744 10560 7750
rect 10508 7686 10560 7692
rect 10416 7404 10468 7410
rect 10416 7346 10468 7352
rect 10428 6798 10456 7346
rect 10520 7002 10548 7686
rect 10980 7546 11008 7890
rect 11428 7880 11480 7886
rect 11428 7822 11480 7828
rect 11612 7880 11664 7886
rect 11612 7822 11664 7828
rect 11440 7546 11468 7822
rect 11520 7744 11572 7750
rect 11520 7686 11572 7692
rect 10968 7540 11020 7546
rect 10968 7482 11020 7488
rect 11428 7540 11480 7546
rect 11428 7482 11480 7488
rect 11532 7342 11560 7686
rect 11520 7336 11572 7342
rect 11520 7278 11572 7284
rect 11624 7002 11652 7822
rect 12452 7546 12480 8230
rect 12440 7540 12492 7546
rect 12440 7482 12492 7488
rect 10508 6996 10560 7002
rect 10508 6938 10560 6944
rect 11612 6996 11664 7002
rect 11612 6938 11664 6944
rect 10416 6792 10468 6798
rect 10416 6734 10468 6740
rect 10428 6390 10456 6734
rect 10416 6384 10468 6390
rect 10416 6326 10468 6332
rect 10416 6248 10468 6254
rect 10416 6190 10468 6196
rect 10428 5710 10456 6190
rect 10520 5778 10548 6938
rect 11624 6798 11652 6938
rect 12820 6866 12848 18022
rect 13372 17746 13400 20402
rect 13636 20324 13688 20330
rect 13636 20266 13688 20272
rect 13544 20256 13596 20262
rect 13544 20198 13596 20204
rect 13556 20058 13584 20198
rect 13544 20052 13596 20058
rect 13544 19994 13596 20000
rect 13648 19938 13676 20266
rect 13556 19910 13676 19938
rect 13556 19310 13584 19910
rect 13636 19780 13688 19786
rect 13636 19722 13688 19728
rect 13648 19378 13676 19722
rect 14188 19712 14240 19718
rect 14188 19654 14240 19660
rect 14200 19446 14228 19654
rect 14188 19440 14240 19446
rect 14188 19382 14240 19388
rect 13636 19372 13688 19378
rect 13636 19314 13688 19320
rect 13544 19304 13596 19310
rect 13544 19246 13596 19252
rect 13556 18834 13584 19246
rect 13544 18828 13596 18834
rect 13544 18770 13596 18776
rect 13452 18148 13504 18154
rect 13452 18090 13504 18096
rect 13360 17740 13412 17746
rect 13360 17682 13412 17688
rect 12900 17264 12952 17270
rect 12900 17206 12952 17212
rect 12912 16794 12940 17206
rect 12900 16788 12952 16794
rect 12900 16730 12952 16736
rect 13360 16040 13412 16046
rect 13360 15982 13412 15988
rect 13372 15638 13400 15982
rect 13360 15632 13412 15638
rect 13360 15574 13412 15580
rect 13464 15026 13492 18090
rect 13542 16824 13598 16833
rect 13542 16759 13598 16768
rect 13556 16726 13584 16759
rect 13544 16720 13596 16726
rect 13544 16662 13596 16668
rect 13556 16250 13584 16662
rect 13544 16244 13596 16250
rect 13544 16186 13596 16192
rect 13556 15638 13584 16186
rect 13648 16182 13676 19314
rect 13728 17672 13780 17678
rect 13728 17614 13780 17620
rect 13740 17270 13768 17614
rect 14004 17536 14056 17542
rect 14004 17478 14056 17484
rect 13728 17264 13780 17270
rect 13728 17206 13780 17212
rect 13636 16176 13688 16182
rect 13636 16118 13688 16124
rect 13726 15872 13782 15881
rect 13726 15807 13782 15816
rect 13740 15706 13768 15807
rect 13728 15700 13780 15706
rect 13728 15642 13780 15648
rect 13544 15632 13596 15638
rect 13544 15574 13596 15580
rect 13556 15434 13584 15574
rect 13544 15428 13596 15434
rect 13544 15370 13596 15376
rect 13452 15020 13504 15026
rect 13452 14962 13504 14968
rect 13360 14884 13412 14890
rect 13360 14826 13412 14832
rect 13372 13734 13400 14826
rect 13464 14618 13492 14962
rect 13452 14612 13504 14618
rect 13452 14554 13504 14560
rect 13360 13728 13412 13734
rect 13360 13670 13412 13676
rect 13084 13252 13136 13258
rect 13084 13194 13136 13200
rect 13176 13252 13228 13258
rect 13176 13194 13228 13200
rect 13096 12986 13124 13194
rect 13084 12980 13136 12986
rect 13084 12922 13136 12928
rect 13188 12850 13216 13194
rect 13176 12844 13228 12850
rect 13176 12786 13228 12792
rect 13542 12472 13598 12481
rect 13542 12407 13598 12416
rect 13556 12374 13584 12407
rect 13544 12368 13596 12374
rect 13544 12310 13596 12316
rect 13176 11552 13228 11558
rect 13176 11494 13228 11500
rect 13188 10674 13216 11494
rect 13176 10668 13228 10674
rect 13176 10610 13228 10616
rect 13084 9920 13136 9926
rect 13084 9862 13136 9868
rect 13096 9586 13124 9862
rect 14016 9722 14044 17478
rect 14096 17196 14148 17202
rect 14096 17138 14148 17144
rect 14108 16726 14136 17138
rect 14096 16720 14148 16726
rect 14096 16662 14148 16668
rect 14188 16108 14240 16114
rect 14188 16050 14240 16056
rect 14200 15502 14228 16050
rect 14188 15496 14240 15502
rect 14188 15438 14240 15444
rect 14200 15162 14228 15438
rect 14292 15366 14320 21270
rect 14568 21078 14596 22066
rect 14924 22092 14976 22098
rect 14924 22034 14976 22040
rect 15016 22092 15068 22098
rect 15016 22034 15068 22040
rect 14936 21554 14964 22034
rect 14924 21548 14976 21554
rect 14924 21490 14976 21496
rect 15028 21434 15056 22034
rect 15212 21894 15240 22607
rect 15488 22137 15516 23258
rect 15474 22128 15530 22137
rect 15474 22063 15530 22072
rect 15200 21888 15252 21894
rect 15200 21830 15252 21836
rect 14936 21406 15056 21434
rect 14648 21140 14700 21146
rect 14648 21082 14700 21088
rect 14832 21140 14884 21146
rect 14832 21082 14884 21088
rect 14556 21072 14608 21078
rect 14556 21014 14608 21020
rect 14372 19508 14424 19514
rect 14372 19450 14424 19456
rect 14384 18766 14412 19450
rect 14372 18760 14424 18766
rect 14372 18702 14424 18708
rect 14464 17876 14516 17882
rect 14464 17818 14516 17824
rect 14372 17808 14424 17814
rect 14372 17750 14424 17756
rect 14384 17202 14412 17750
rect 14372 17196 14424 17202
rect 14372 17138 14424 17144
rect 14476 16794 14504 17818
rect 14568 17320 14596 21014
rect 14660 20788 14688 21082
rect 14844 20942 14872 21082
rect 14936 20942 14964 21406
rect 15014 21040 15070 21049
rect 15014 20975 15070 20984
rect 14832 20936 14884 20942
rect 14832 20878 14884 20884
rect 14924 20936 14976 20942
rect 14924 20878 14976 20884
rect 14936 20788 14964 20878
rect 15028 20874 15056 20975
rect 15016 20868 15068 20874
rect 15016 20810 15068 20816
rect 14660 20760 14964 20788
rect 14660 20602 14688 20760
rect 14648 20596 14700 20602
rect 14648 20538 14700 20544
rect 15200 20324 15252 20330
rect 15200 20266 15252 20272
rect 14648 20052 14700 20058
rect 14648 19994 14700 20000
rect 14660 19378 14688 19994
rect 15212 19378 15240 20266
rect 14648 19372 14700 19378
rect 14648 19314 14700 19320
rect 14832 19372 14884 19378
rect 14832 19314 14884 19320
rect 15200 19372 15252 19378
rect 15200 19314 15252 19320
rect 14740 19304 14792 19310
rect 14740 19246 14792 19252
rect 14752 18850 14780 19246
rect 14660 18822 14780 18850
rect 14660 18358 14688 18822
rect 14740 18692 14792 18698
rect 14740 18634 14792 18640
rect 14648 18352 14700 18358
rect 14648 18294 14700 18300
rect 14752 18290 14780 18634
rect 14844 18290 14872 19314
rect 15212 18834 15240 19314
rect 15200 18828 15252 18834
rect 15200 18770 15252 18776
rect 14924 18760 14976 18766
rect 14922 18728 14924 18737
rect 14976 18728 14978 18737
rect 14922 18663 14978 18672
rect 15212 18426 15240 18770
rect 15292 18760 15344 18766
rect 15292 18702 15344 18708
rect 15304 18426 15332 18702
rect 15200 18420 15252 18426
rect 15200 18362 15252 18368
rect 15292 18420 15344 18426
rect 15292 18362 15344 18368
rect 15108 18352 15160 18358
rect 15108 18294 15160 18300
rect 14740 18284 14792 18290
rect 14740 18226 14792 18232
rect 14832 18284 14884 18290
rect 14832 18226 14884 18232
rect 14568 17292 14688 17320
rect 14556 17196 14608 17202
rect 14556 17138 14608 17144
rect 14464 16788 14516 16794
rect 14464 16730 14516 16736
rect 14476 16522 14504 16730
rect 14568 16590 14596 17138
rect 14556 16584 14608 16590
rect 14556 16526 14608 16532
rect 14464 16516 14516 16522
rect 14464 16458 14516 16464
rect 14568 15706 14596 16526
rect 14660 15858 14688 17292
rect 14752 17202 14780 18226
rect 14740 17196 14792 17202
rect 14740 17138 14792 17144
rect 14844 16658 14872 18226
rect 15016 17604 15068 17610
rect 15016 17546 15068 17552
rect 15028 16998 15056 17546
rect 15120 17218 15148 18294
rect 15200 18080 15252 18086
rect 15200 18022 15252 18028
rect 15212 17678 15240 18022
rect 15200 17672 15252 17678
rect 15200 17614 15252 17620
rect 15566 17640 15622 17649
rect 15566 17575 15568 17584
rect 15620 17575 15622 17584
rect 15568 17546 15620 17552
rect 15120 17202 15240 17218
rect 15120 17196 15252 17202
rect 15120 17190 15200 17196
rect 15016 16992 15068 16998
rect 15016 16934 15068 16940
rect 14832 16652 14884 16658
rect 14832 16594 14884 16600
rect 14924 16040 14976 16046
rect 14924 15982 14976 15988
rect 14660 15830 14780 15858
rect 14556 15700 14608 15706
rect 14556 15642 14608 15648
rect 14648 15700 14700 15706
rect 14648 15642 14700 15648
rect 14464 15496 14516 15502
rect 14464 15438 14516 15444
rect 14280 15360 14332 15366
rect 14280 15302 14332 15308
rect 14188 15156 14240 15162
rect 14188 15098 14240 15104
rect 14096 14476 14148 14482
rect 14096 14418 14148 14424
rect 14004 9716 14056 9722
rect 14004 9658 14056 9664
rect 13728 9648 13780 9654
rect 13728 9590 13780 9596
rect 13084 9580 13136 9586
rect 13084 9522 13136 9528
rect 13740 7546 13768 9590
rect 13728 7540 13780 7546
rect 13728 7482 13780 7488
rect 13740 7313 13768 7482
rect 13726 7304 13782 7313
rect 13726 7239 13782 7248
rect 12900 7200 12952 7206
rect 12900 7142 12952 7148
rect 12912 6934 12940 7142
rect 12900 6928 12952 6934
rect 12900 6870 12952 6876
rect 12808 6860 12860 6866
rect 12808 6802 12860 6808
rect 12912 6798 12940 6870
rect 11612 6792 11664 6798
rect 11612 6734 11664 6740
rect 12900 6792 12952 6798
rect 12900 6734 12952 6740
rect 14108 6746 14136 14418
rect 14292 13938 14320 15302
rect 14476 14890 14504 15438
rect 14464 14884 14516 14890
rect 14464 14826 14516 14832
rect 14568 14618 14596 15642
rect 14660 15570 14688 15642
rect 14648 15564 14700 15570
rect 14648 15506 14700 15512
rect 14648 14816 14700 14822
rect 14648 14758 14700 14764
rect 14556 14612 14608 14618
rect 14556 14554 14608 14560
rect 14372 14544 14424 14550
rect 14372 14486 14424 14492
rect 14384 14006 14412 14486
rect 14372 14000 14424 14006
rect 14372 13942 14424 13948
rect 14280 13932 14332 13938
rect 14280 13874 14332 13880
rect 14568 13326 14596 14554
rect 14660 14482 14688 14758
rect 14648 14476 14700 14482
rect 14648 14418 14700 14424
rect 14556 13320 14608 13326
rect 14556 13262 14608 13268
rect 14752 12850 14780 15830
rect 14832 13184 14884 13190
rect 14832 13126 14884 13132
rect 14740 12844 14792 12850
rect 14740 12786 14792 12792
rect 14844 11626 14872 13126
rect 14936 12986 14964 15982
rect 15120 15502 15148 17190
rect 15200 17138 15252 17144
rect 15292 17060 15344 17066
rect 15292 17002 15344 17008
rect 15304 16726 15332 17002
rect 15476 16992 15528 16998
rect 15476 16934 15528 16940
rect 15292 16720 15344 16726
rect 15292 16662 15344 16668
rect 15488 16590 15516 16934
rect 15476 16584 15528 16590
rect 15476 16526 15528 16532
rect 15292 15904 15344 15910
rect 15292 15846 15344 15852
rect 15108 15496 15160 15502
rect 15108 15438 15160 15444
rect 15198 15464 15254 15473
rect 15198 15399 15254 15408
rect 15016 15088 15068 15094
rect 15016 15030 15068 15036
rect 15028 14278 15056 15030
rect 15212 15026 15240 15399
rect 15200 15020 15252 15026
rect 15200 14962 15252 14968
rect 15304 14822 15332 15846
rect 15476 15496 15528 15502
rect 15476 15438 15528 15444
rect 15488 14958 15516 15438
rect 15568 15020 15620 15026
rect 15568 14962 15620 14968
rect 15476 14952 15528 14958
rect 15580 14929 15608 14962
rect 15476 14894 15528 14900
rect 15566 14920 15622 14929
rect 15566 14855 15622 14864
rect 15292 14816 15344 14822
rect 15292 14758 15344 14764
rect 15568 14408 15620 14414
rect 15568 14350 15620 14356
rect 15016 14272 15068 14278
rect 15016 14214 15068 14220
rect 14924 12980 14976 12986
rect 14924 12922 14976 12928
rect 14832 11620 14884 11626
rect 14832 11562 14884 11568
rect 14280 11076 14332 11082
rect 14280 11018 14332 11024
rect 14292 7426 14320 11018
rect 14924 10056 14976 10062
rect 14924 9998 14976 10004
rect 14936 8974 14964 9998
rect 14924 8968 14976 8974
rect 14924 8910 14976 8916
rect 14464 8832 14516 8838
rect 14464 8774 14516 8780
rect 14476 7886 14504 8774
rect 15028 8294 15056 14214
rect 15580 13938 15608 14350
rect 15568 13932 15620 13938
rect 15568 13874 15620 13880
rect 15672 13530 15700 24890
rect 16500 24886 16528 26930
rect 16488 24880 16540 24886
rect 16488 24822 16540 24828
rect 16488 24608 16540 24614
rect 16488 24550 16540 24556
rect 16500 24274 16528 24550
rect 16488 24268 16540 24274
rect 16488 24210 16540 24216
rect 16580 24200 16632 24206
rect 16580 24142 16632 24148
rect 16488 24132 16540 24138
rect 16488 24074 16540 24080
rect 16500 23186 16528 24074
rect 16592 23730 16620 24142
rect 16580 23724 16632 23730
rect 16580 23666 16632 23672
rect 16488 23180 16540 23186
rect 16488 23122 16540 23128
rect 16396 23112 16448 23118
rect 16396 23054 16448 23060
rect 16120 23044 16172 23050
rect 16120 22986 16172 22992
rect 15936 22432 15988 22438
rect 15936 22374 15988 22380
rect 15752 22228 15804 22234
rect 15752 22170 15804 22176
rect 15764 21962 15792 22170
rect 15752 21956 15804 21962
rect 15752 21898 15804 21904
rect 15948 21690 15976 22374
rect 15936 21684 15988 21690
rect 15936 21626 15988 21632
rect 16132 21321 16160 22986
rect 16304 22024 16356 22030
rect 16408 21978 16436 23054
rect 16488 22636 16540 22642
rect 16488 22578 16540 22584
rect 16500 22234 16528 22578
rect 16488 22228 16540 22234
rect 16488 22170 16540 22176
rect 16684 22094 16712 37198
rect 18064 37126 18092 39200
rect 19996 37262 20024 39200
rect 21928 37346 21956 39200
rect 23860 37398 23888 39200
rect 23848 37392 23900 37398
rect 21928 37318 22232 37346
rect 23848 37334 23900 37340
rect 19984 37256 20036 37262
rect 19984 37198 20036 37204
rect 22204 37194 22232 37318
rect 25792 37262 25820 39200
rect 28368 37262 28396 39200
rect 30300 37330 30328 39200
rect 28908 37324 28960 37330
rect 28908 37266 28960 37272
rect 30288 37324 30340 37330
rect 30288 37266 30340 37272
rect 25780 37256 25832 37262
rect 25780 37198 25832 37204
rect 28356 37256 28408 37262
rect 28356 37198 28408 37204
rect 20260 37188 20312 37194
rect 20260 37130 20312 37136
rect 22192 37188 22244 37194
rect 22192 37130 22244 37136
rect 28632 37188 28684 37194
rect 28632 37130 28684 37136
rect 18052 37120 18104 37126
rect 18052 37062 18104 37068
rect 19574 37020 19882 37040
rect 19574 37018 19580 37020
rect 19636 37018 19660 37020
rect 19716 37018 19740 37020
rect 19796 37018 19820 37020
rect 19876 37018 19882 37020
rect 19636 36966 19638 37018
rect 19818 36966 19820 37018
rect 19574 36964 19580 36966
rect 19636 36964 19660 36966
rect 19716 36964 19740 36966
rect 19796 36964 19820 36966
rect 19876 36964 19882 36966
rect 19574 36944 19882 36964
rect 19432 36712 19484 36718
rect 19432 36654 19484 36660
rect 19444 36378 19472 36654
rect 19432 36372 19484 36378
rect 19432 36314 19484 36320
rect 20076 36236 20128 36242
rect 20076 36178 20128 36184
rect 19248 36168 19300 36174
rect 19248 36110 19300 36116
rect 19340 36168 19392 36174
rect 19340 36110 19392 36116
rect 17776 35828 17828 35834
rect 17776 35770 17828 35776
rect 17408 34604 17460 34610
rect 17408 34546 17460 34552
rect 17420 34202 17448 34546
rect 17408 34196 17460 34202
rect 17408 34138 17460 34144
rect 17788 33658 17816 35770
rect 19260 35766 19288 36110
rect 18144 35760 18196 35766
rect 18144 35702 18196 35708
rect 19248 35760 19300 35766
rect 19248 35702 19300 35708
rect 17868 35012 17920 35018
rect 17868 34954 17920 34960
rect 17880 34610 17908 34954
rect 18156 34746 18184 35702
rect 19352 35630 19380 36110
rect 19574 35932 19882 35952
rect 19574 35930 19580 35932
rect 19636 35930 19660 35932
rect 19716 35930 19740 35932
rect 19796 35930 19820 35932
rect 19876 35930 19882 35932
rect 19636 35878 19638 35930
rect 19818 35878 19820 35930
rect 19574 35876 19580 35878
rect 19636 35876 19660 35878
rect 19716 35876 19740 35878
rect 19796 35876 19820 35878
rect 19876 35876 19882 35878
rect 19574 35856 19882 35876
rect 19340 35624 19392 35630
rect 19340 35566 19392 35572
rect 18696 35488 18748 35494
rect 18696 35430 18748 35436
rect 18708 35290 18736 35430
rect 18328 35284 18380 35290
rect 18328 35226 18380 35232
rect 18696 35284 18748 35290
rect 18696 35226 18748 35232
rect 18144 34740 18196 34746
rect 18144 34682 18196 34688
rect 18340 34610 18368 35226
rect 18420 34944 18472 34950
rect 18420 34886 18472 34892
rect 18432 34610 18460 34886
rect 19352 34746 19380 35566
rect 20088 35494 20116 36178
rect 20076 35488 20128 35494
rect 20076 35430 20128 35436
rect 19574 34844 19882 34864
rect 19574 34842 19580 34844
rect 19636 34842 19660 34844
rect 19716 34842 19740 34844
rect 19796 34842 19820 34844
rect 19876 34842 19882 34844
rect 19636 34790 19638 34842
rect 19818 34790 19820 34842
rect 19574 34788 19580 34790
rect 19636 34788 19660 34790
rect 19716 34788 19740 34790
rect 19796 34788 19820 34790
rect 19876 34788 19882 34790
rect 19574 34768 19882 34788
rect 19340 34740 19392 34746
rect 19340 34682 19392 34688
rect 17868 34604 17920 34610
rect 17868 34546 17920 34552
rect 18328 34604 18380 34610
rect 18328 34546 18380 34552
rect 18420 34604 18472 34610
rect 18420 34546 18472 34552
rect 20168 34604 20220 34610
rect 20168 34546 20220 34552
rect 18340 34474 18368 34546
rect 18328 34468 18380 34474
rect 18328 34410 18380 34416
rect 18340 33862 18368 34410
rect 18432 34202 18460 34546
rect 18420 34196 18472 34202
rect 18420 34138 18472 34144
rect 18420 33992 18472 33998
rect 19248 33992 19300 33998
rect 18420 33934 18472 33940
rect 18328 33856 18380 33862
rect 18328 33798 18380 33804
rect 17776 33652 17828 33658
rect 17776 33594 17828 33600
rect 17132 33584 17184 33590
rect 17132 33526 17184 33532
rect 17144 33046 17172 33526
rect 18432 33114 18460 33934
rect 18524 33930 18828 33946
rect 19248 33934 19300 33940
rect 18512 33924 18840 33930
rect 18564 33918 18788 33924
rect 18512 33866 18564 33872
rect 18788 33866 18840 33872
rect 18524 33402 18552 33866
rect 18524 33374 18644 33402
rect 18420 33108 18472 33114
rect 18420 33050 18472 33056
rect 17132 33040 17184 33046
rect 17132 32982 17184 32988
rect 17144 32230 17172 32982
rect 18328 32904 18380 32910
rect 18328 32846 18380 32852
rect 18512 32904 18564 32910
rect 18512 32846 18564 32852
rect 17224 32836 17276 32842
rect 17224 32778 17276 32784
rect 18236 32836 18288 32842
rect 18236 32778 18288 32784
rect 17132 32224 17184 32230
rect 17132 32166 17184 32172
rect 17040 32020 17092 32026
rect 17040 31962 17092 31968
rect 16948 30864 17000 30870
rect 16948 30806 17000 30812
rect 16960 30258 16988 30806
rect 16948 30252 17000 30258
rect 16948 30194 17000 30200
rect 17052 29238 17080 31962
rect 17236 31958 17264 32778
rect 17592 32768 17644 32774
rect 17592 32710 17644 32716
rect 17224 31952 17276 31958
rect 17224 31894 17276 31900
rect 17500 30592 17552 30598
rect 17500 30534 17552 30540
rect 17040 29232 17092 29238
rect 17040 29174 17092 29180
rect 17224 29028 17276 29034
rect 17224 28970 17276 28976
rect 17132 28620 17184 28626
rect 17132 28562 17184 28568
rect 17040 28076 17092 28082
rect 17040 28018 17092 28024
rect 17052 27606 17080 28018
rect 17144 27946 17172 28562
rect 17236 28082 17264 28970
rect 17224 28076 17276 28082
rect 17224 28018 17276 28024
rect 17132 27940 17184 27946
rect 17132 27882 17184 27888
rect 17040 27600 17092 27606
rect 17040 27542 17092 27548
rect 16764 27532 16816 27538
rect 16948 27532 17000 27538
rect 16816 27492 16948 27520
rect 16764 27474 16816 27480
rect 16948 27474 17000 27480
rect 17316 27328 17368 27334
rect 17316 27270 17368 27276
rect 17328 26382 17356 27270
rect 16764 26376 16816 26382
rect 16764 26318 16816 26324
rect 17316 26376 17368 26382
rect 17316 26318 17368 26324
rect 16776 25294 16804 26318
rect 17224 25900 17276 25906
rect 17224 25842 17276 25848
rect 16764 25288 16816 25294
rect 16764 25230 16816 25236
rect 17132 25288 17184 25294
rect 17132 25230 17184 25236
rect 16856 25220 16908 25226
rect 16856 25162 16908 25168
rect 16764 24676 16816 24682
rect 16764 24618 16816 24624
rect 16776 24206 16804 24618
rect 16764 24200 16816 24206
rect 16764 24142 16816 24148
rect 16764 23792 16816 23798
rect 16868 23780 16896 25162
rect 17040 24812 17092 24818
rect 17040 24754 17092 24760
rect 17052 24410 17080 24754
rect 17144 24682 17172 25230
rect 17236 24886 17264 25842
rect 17328 25226 17356 26318
rect 17408 26240 17460 26246
rect 17408 26182 17460 26188
rect 17420 25906 17448 26182
rect 17408 25900 17460 25906
rect 17408 25842 17460 25848
rect 17420 25362 17448 25842
rect 17408 25356 17460 25362
rect 17408 25298 17460 25304
rect 17316 25220 17368 25226
rect 17316 25162 17368 25168
rect 17224 24880 17276 24886
rect 17224 24822 17276 24828
rect 17408 24744 17460 24750
rect 17408 24686 17460 24692
rect 17132 24676 17184 24682
rect 17132 24618 17184 24624
rect 17040 24404 17092 24410
rect 17040 24346 17092 24352
rect 16816 23752 16896 23780
rect 16764 23734 16816 23740
rect 16776 23050 16804 23734
rect 17052 23730 17080 24346
rect 17420 24206 17448 24686
rect 17224 24200 17276 24206
rect 17224 24142 17276 24148
rect 17408 24200 17460 24206
rect 17408 24142 17460 24148
rect 17236 23866 17264 24142
rect 17224 23860 17276 23866
rect 17224 23802 17276 23808
rect 16948 23724 17000 23730
rect 16948 23666 17000 23672
rect 17040 23724 17092 23730
rect 17040 23666 17092 23672
rect 16764 23044 16816 23050
rect 16764 22986 16816 22992
rect 16960 22624 16988 23666
rect 17512 22778 17540 30534
rect 17604 29510 17632 32710
rect 18248 32434 18276 32778
rect 18340 32434 18368 32846
rect 18524 32434 18552 32846
rect 18616 32502 18644 33374
rect 19260 33046 19288 33934
rect 20180 33862 20208 34546
rect 20168 33856 20220 33862
rect 20168 33798 20220 33804
rect 19574 33756 19882 33776
rect 19574 33754 19580 33756
rect 19636 33754 19660 33756
rect 19716 33754 19740 33756
rect 19796 33754 19820 33756
rect 19876 33754 19882 33756
rect 19636 33702 19638 33754
rect 19818 33702 19820 33754
rect 19574 33700 19580 33702
rect 19636 33700 19660 33702
rect 19716 33700 19740 33702
rect 19796 33700 19820 33702
rect 19876 33700 19882 33702
rect 19574 33680 19882 33700
rect 19248 33040 19300 33046
rect 19248 32982 19300 32988
rect 18788 32972 18840 32978
rect 18788 32914 18840 32920
rect 18604 32496 18656 32502
rect 18604 32438 18656 32444
rect 18236 32428 18288 32434
rect 18236 32370 18288 32376
rect 18328 32428 18380 32434
rect 18328 32370 18380 32376
rect 18512 32428 18564 32434
rect 18512 32370 18564 32376
rect 18248 32026 18276 32370
rect 18236 32020 18288 32026
rect 18236 31962 18288 31968
rect 17960 31816 18012 31822
rect 17960 31758 18012 31764
rect 18052 31816 18104 31822
rect 18052 31758 18104 31764
rect 17972 31414 18000 31758
rect 17960 31408 18012 31414
rect 17960 31350 18012 31356
rect 18064 31346 18092 31758
rect 18236 31680 18288 31686
rect 18236 31622 18288 31628
rect 18248 31346 18276 31622
rect 18052 31340 18104 31346
rect 18052 31282 18104 31288
rect 18236 31340 18288 31346
rect 18236 31282 18288 31288
rect 18064 30870 18092 31282
rect 18052 30864 18104 30870
rect 18052 30806 18104 30812
rect 17868 30252 17920 30258
rect 17868 30194 17920 30200
rect 17880 29646 17908 30194
rect 18248 30122 18276 31282
rect 18340 31278 18368 32370
rect 18512 31340 18564 31346
rect 18512 31282 18564 31288
rect 18328 31272 18380 31278
rect 18328 31214 18380 31220
rect 18328 31136 18380 31142
rect 18524 31090 18552 31282
rect 18328 31078 18380 31084
rect 18340 30802 18368 31078
rect 18432 31062 18552 31090
rect 18328 30796 18380 30802
rect 18328 30738 18380 30744
rect 18236 30116 18288 30122
rect 18236 30058 18288 30064
rect 18432 30054 18460 31062
rect 18420 30048 18472 30054
rect 18050 30016 18106 30025
rect 18420 29990 18472 29996
rect 18050 29951 18106 29960
rect 17868 29640 17920 29646
rect 17868 29582 17920 29588
rect 17592 29504 17644 29510
rect 17592 29446 17644 29452
rect 17604 29170 17632 29446
rect 17960 29232 18012 29238
rect 17960 29174 18012 29180
rect 17592 29164 17644 29170
rect 17592 29106 17644 29112
rect 17604 27606 17632 29106
rect 17592 27600 17644 27606
rect 17592 27542 17644 27548
rect 17972 27402 18000 29174
rect 18064 29034 18092 29951
rect 18604 29096 18656 29102
rect 18604 29038 18656 29044
rect 18052 29028 18104 29034
rect 18052 28970 18104 28976
rect 18512 29028 18564 29034
rect 18512 28970 18564 28976
rect 18052 27872 18104 27878
rect 18052 27814 18104 27820
rect 17960 27396 18012 27402
rect 17960 27338 18012 27344
rect 17960 26784 18012 26790
rect 17960 26726 18012 26732
rect 17684 26512 17736 26518
rect 17684 26454 17736 26460
rect 17696 26382 17724 26454
rect 17684 26376 17736 26382
rect 17684 26318 17736 26324
rect 17776 26376 17828 26382
rect 17776 26318 17828 26324
rect 17696 25906 17724 26318
rect 17788 26042 17816 26318
rect 17776 26036 17828 26042
rect 17776 25978 17828 25984
rect 17684 25900 17736 25906
rect 17684 25842 17736 25848
rect 17972 25294 18000 26726
rect 18064 25702 18092 27814
rect 18420 27124 18472 27130
rect 18420 27066 18472 27072
rect 18432 26790 18460 27066
rect 18420 26784 18472 26790
rect 18420 26726 18472 26732
rect 18144 26580 18196 26586
rect 18144 26522 18196 26528
rect 18156 26382 18184 26522
rect 18432 26382 18460 26726
rect 18144 26376 18196 26382
rect 18144 26318 18196 26324
rect 18420 26376 18472 26382
rect 18420 26318 18472 26324
rect 18156 25974 18184 26318
rect 18236 26036 18288 26042
rect 18236 25978 18288 25984
rect 18144 25968 18196 25974
rect 18144 25910 18196 25916
rect 18052 25696 18104 25702
rect 18052 25638 18104 25644
rect 17960 25288 18012 25294
rect 17960 25230 18012 25236
rect 17960 24948 18012 24954
rect 17960 24890 18012 24896
rect 17684 24676 17736 24682
rect 17684 24618 17736 24624
rect 17696 23118 17724 24618
rect 17972 24410 18000 24890
rect 17960 24404 18012 24410
rect 17960 24346 18012 24352
rect 17776 24200 17828 24206
rect 17776 24142 17828 24148
rect 17788 23662 17816 24142
rect 17868 24064 17920 24070
rect 17868 24006 17920 24012
rect 17880 23798 17908 24006
rect 17868 23792 17920 23798
rect 17868 23734 17920 23740
rect 17776 23656 17828 23662
rect 17776 23598 17828 23604
rect 18064 23594 18092 25638
rect 18248 25294 18276 25978
rect 18236 25288 18288 25294
rect 18236 25230 18288 25236
rect 18328 25288 18380 25294
rect 18328 25230 18380 25236
rect 18144 25220 18196 25226
rect 18144 25162 18196 25168
rect 18156 23866 18184 25162
rect 18236 25152 18288 25158
rect 18236 25094 18288 25100
rect 18144 23860 18196 23866
rect 18144 23802 18196 23808
rect 18052 23588 18104 23594
rect 18052 23530 18104 23536
rect 17684 23112 17736 23118
rect 17684 23054 17736 23060
rect 17592 23044 17644 23050
rect 17592 22986 17644 22992
rect 17500 22772 17552 22778
rect 17500 22714 17552 22720
rect 17040 22636 17092 22642
rect 16960 22596 17040 22624
rect 17040 22578 17092 22584
rect 17052 22409 17080 22578
rect 17038 22400 17094 22409
rect 17038 22335 17094 22344
rect 17604 22166 17632 22986
rect 17592 22160 17644 22166
rect 17592 22102 17644 22108
rect 16356 21972 16436 21978
rect 16304 21966 16436 21972
rect 16316 21950 16436 21966
rect 16592 22066 16712 22094
rect 16304 21344 16356 21350
rect 16118 21312 16174 21321
rect 16304 21286 16356 21292
rect 16118 21247 16174 21256
rect 16120 21072 16172 21078
rect 16120 21014 16172 21020
rect 16132 20874 16160 21014
rect 16316 20942 16344 21286
rect 16304 20936 16356 20942
rect 16304 20878 16356 20884
rect 16120 20868 16172 20874
rect 16120 20810 16172 20816
rect 15752 20256 15804 20262
rect 15750 20224 15752 20233
rect 15804 20224 15806 20233
rect 15750 20159 15806 20168
rect 16028 19780 16080 19786
rect 16028 19722 16080 19728
rect 15936 19440 15988 19446
rect 15934 19408 15936 19417
rect 15988 19408 15990 19417
rect 16040 19378 16068 19722
rect 15934 19343 15990 19352
rect 16028 19372 16080 19378
rect 16028 19314 16080 19320
rect 15936 18420 15988 18426
rect 15936 18362 15988 18368
rect 15844 16448 15896 16454
rect 15844 16390 15896 16396
rect 15856 16114 15884 16390
rect 15844 16108 15896 16114
rect 15844 16050 15896 16056
rect 15752 15496 15804 15502
rect 15752 15438 15804 15444
rect 15764 14006 15792 15438
rect 15844 15360 15896 15366
rect 15844 15302 15896 15308
rect 15856 15094 15884 15302
rect 15844 15088 15896 15094
rect 15842 15056 15844 15065
rect 15896 15056 15898 15065
rect 15842 14991 15898 15000
rect 15948 14890 15976 18362
rect 16040 18222 16068 19314
rect 16132 19174 16160 20810
rect 16316 20233 16344 20878
rect 16302 20224 16358 20233
rect 16302 20159 16358 20168
rect 16212 19304 16264 19310
rect 16212 19246 16264 19252
rect 16120 19168 16172 19174
rect 16120 19110 16172 19116
rect 16224 18766 16252 19246
rect 16408 19242 16436 21950
rect 16488 21956 16540 21962
rect 16488 21898 16540 21904
rect 16500 21690 16528 21898
rect 16488 21684 16540 21690
rect 16488 21626 16540 21632
rect 16486 20904 16542 20913
rect 16486 20839 16542 20848
rect 16500 20806 16528 20839
rect 16488 20800 16540 20806
rect 16488 20742 16540 20748
rect 16396 19236 16448 19242
rect 16396 19178 16448 19184
rect 16488 19168 16540 19174
rect 16488 19110 16540 19116
rect 16212 18760 16264 18766
rect 16212 18702 16264 18708
rect 16120 18692 16172 18698
rect 16120 18634 16172 18640
rect 16132 18426 16160 18634
rect 16120 18420 16172 18426
rect 16120 18362 16172 18368
rect 16028 18216 16080 18222
rect 16028 18158 16080 18164
rect 16304 16992 16356 16998
rect 16304 16934 16356 16940
rect 16120 16652 16172 16658
rect 16120 16594 16172 16600
rect 16132 16114 16160 16594
rect 16316 16454 16344 16934
rect 16304 16448 16356 16454
rect 16304 16390 16356 16396
rect 16120 16108 16172 16114
rect 16120 16050 16172 16056
rect 16396 15904 16448 15910
rect 16396 15846 16448 15852
rect 16408 15502 16436 15846
rect 16396 15496 16448 15502
rect 16396 15438 16448 15444
rect 16500 15314 16528 19110
rect 16592 17338 16620 22066
rect 17604 21622 17632 22102
rect 17592 21616 17644 21622
rect 17592 21558 17644 21564
rect 18052 21480 18104 21486
rect 18052 21422 18104 21428
rect 17224 21344 17276 21350
rect 17224 21286 17276 21292
rect 17236 21078 17264 21286
rect 17224 21072 17276 21078
rect 17224 21014 17276 21020
rect 18064 21010 18092 21422
rect 18052 21004 18104 21010
rect 18052 20946 18104 20952
rect 16764 20052 16816 20058
rect 16764 19994 16816 20000
rect 16776 19310 16804 19994
rect 17776 19780 17828 19786
rect 17776 19722 17828 19728
rect 17788 19378 17816 19722
rect 18064 19446 18092 20946
rect 18144 20868 18196 20874
rect 18144 20810 18196 20816
rect 18156 20330 18184 20810
rect 18248 20602 18276 25094
rect 18340 24750 18368 25230
rect 18524 25158 18552 28970
rect 18616 28558 18644 29038
rect 18800 28762 18828 32914
rect 19340 32904 19392 32910
rect 19340 32846 19392 32852
rect 19352 30938 19380 32846
rect 19574 32668 19882 32688
rect 19574 32666 19580 32668
rect 19636 32666 19660 32668
rect 19716 32666 19740 32668
rect 19796 32666 19820 32668
rect 19876 32666 19882 32668
rect 19636 32614 19638 32666
rect 19818 32614 19820 32666
rect 19574 32612 19580 32614
rect 19636 32612 19660 32614
rect 19716 32612 19740 32614
rect 19796 32612 19820 32614
rect 19876 32612 19882 32614
rect 19574 32592 19882 32612
rect 20272 31754 20300 37130
rect 22284 37120 22336 37126
rect 22284 37062 22336 37068
rect 24584 37120 24636 37126
rect 24584 37062 24636 37068
rect 26148 37120 26200 37126
rect 26148 37062 26200 37068
rect 21272 36780 21324 36786
rect 21272 36722 21324 36728
rect 21284 36310 21312 36722
rect 21732 36712 21784 36718
rect 21732 36654 21784 36660
rect 21744 36378 21772 36654
rect 21732 36372 21784 36378
rect 21732 36314 21784 36320
rect 21272 36304 21324 36310
rect 21272 36246 21324 36252
rect 21284 36174 21312 36246
rect 21272 36168 21324 36174
rect 21272 36110 21324 36116
rect 22100 36168 22152 36174
rect 22100 36110 22152 36116
rect 21088 35692 21140 35698
rect 21088 35634 21140 35640
rect 20812 35080 20864 35086
rect 20812 35022 20864 35028
rect 20824 34746 20852 35022
rect 21100 34746 21128 35634
rect 21284 35018 21312 36110
rect 22112 35766 22140 36110
rect 22100 35760 22152 35766
rect 22100 35702 22152 35708
rect 22112 35290 22140 35702
rect 22100 35284 22152 35290
rect 22100 35226 22152 35232
rect 21272 35012 21324 35018
rect 21272 34954 21324 34960
rect 22192 34944 22244 34950
rect 22192 34886 22244 34892
rect 22204 34746 22232 34886
rect 20812 34740 20864 34746
rect 20812 34682 20864 34688
rect 21088 34740 21140 34746
rect 21088 34682 21140 34688
rect 22192 34740 22244 34746
rect 22192 34682 22244 34688
rect 22296 34066 22324 37062
rect 24596 36922 24624 37062
rect 24584 36916 24636 36922
rect 24584 36858 24636 36864
rect 23480 36780 23532 36786
rect 23480 36722 23532 36728
rect 23848 36780 23900 36786
rect 23848 36722 23900 36728
rect 23492 36650 23520 36722
rect 23480 36644 23532 36650
rect 23480 36586 23532 36592
rect 23492 35086 23520 36586
rect 23860 36378 23888 36722
rect 24400 36712 24452 36718
rect 24400 36654 24452 36660
rect 25688 36712 25740 36718
rect 25688 36654 25740 36660
rect 23848 36372 23900 36378
rect 23848 36314 23900 36320
rect 24412 36174 24440 36654
rect 25700 36378 25728 36654
rect 25688 36372 25740 36378
rect 25688 36314 25740 36320
rect 23664 36168 23716 36174
rect 23664 36110 23716 36116
rect 23848 36168 23900 36174
rect 23848 36110 23900 36116
rect 24400 36168 24452 36174
rect 24400 36110 24452 36116
rect 24492 36168 24544 36174
rect 24492 36110 24544 36116
rect 23676 36038 23704 36110
rect 23664 36032 23716 36038
rect 23664 35974 23716 35980
rect 23676 35562 23704 35974
rect 23860 35766 23888 36110
rect 24504 36038 24532 36110
rect 24492 36032 24544 36038
rect 24492 35974 24544 35980
rect 23848 35760 23900 35766
rect 23848 35702 23900 35708
rect 23664 35556 23716 35562
rect 23664 35498 23716 35504
rect 24504 35222 24532 35974
rect 24952 35624 25004 35630
rect 24952 35566 25004 35572
rect 24492 35216 24544 35222
rect 24492 35158 24544 35164
rect 23480 35080 23532 35086
rect 23480 35022 23532 35028
rect 22652 35012 22704 35018
rect 22652 34954 22704 34960
rect 22664 34678 22692 34954
rect 24504 34678 24532 35158
rect 24964 34950 24992 35566
rect 25136 35080 25188 35086
rect 25136 35022 25188 35028
rect 24952 34944 25004 34950
rect 24952 34886 25004 34892
rect 22652 34672 22704 34678
rect 22652 34614 22704 34620
rect 24492 34672 24544 34678
rect 24492 34614 24544 34620
rect 22664 34066 22692 34614
rect 24964 34610 24992 34886
rect 25148 34610 25176 35022
rect 24952 34604 25004 34610
rect 24952 34546 25004 34552
rect 25136 34604 25188 34610
rect 25136 34546 25188 34552
rect 25148 34202 25176 34546
rect 25136 34196 25188 34202
rect 25136 34138 25188 34144
rect 24952 34128 25004 34134
rect 24952 34070 25004 34076
rect 22284 34060 22336 34066
rect 22284 34002 22336 34008
rect 22652 34060 22704 34066
rect 22652 34002 22704 34008
rect 23388 34060 23440 34066
rect 23388 34002 23440 34008
rect 23204 33992 23256 33998
rect 23204 33934 23256 33940
rect 23216 33522 23244 33934
rect 23400 33590 23428 34002
rect 24676 33924 24728 33930
rect 24676 33866 24728 33872
rect 23388 33584 23440 33590
rect 23388 33526 23440 33532
rect 24688 33522 24716 33866
rect 22468 33516 22520 33522
rect 22468 33458 22520 33464
rect 23204 33516 23256 33522
rect 23204 33458 23256 33464
rect 24676 33516 24728 33522
rect 24676 33458 24728 33464
rect 22008 32904 22060 32910
rect 22008 32846 22060 32852
rect 22284 32904 22336 32910
rect 22284 32846 22336 32852
rect 22020 32366 22048 32846
rect 22008 32360 22060 32366
rect 22008 32302 22060 32308
rect 21180 32224 21232 32230
rect 21180 32166 21232 32172
rect 20996 31884 21048 31890
rect 20996 31826 21048 31832
rect 20180 31726 20300 31754
rect 19574 31580 19882 31600
rect 19574 31578 19580 31580
rect 19636 31578 19660 31580
rect 19716 31578 19740 31580
rect 19796 31578 19820 31580
rect 19876 31578 19882 31580
rect 19636 31526 19638 31578
rect 19818 31526 19820 31578
rect 19574 31524 19580 31526
rect 19636 31524 19660 31526
rect 19716 31524 19740 31526
rect 19796 31524 19820 31526
rect 19876 31524 19882 31526
rect 19574 31504 19882 31524
rect 19524 31408 19576 31414
rect 19524 31350 19576 31356
rect 19340 30932 19392 30938
rect 19340 30874 19392 30880
rect 19352 30734 19380 30874
rect 19340 30728 19392 30734
rect 19340 30670 19392 30676
rect 19432 30728 19484 30734
rect 19432 30670 19484 30676
rect 19444 30598 19472 30670
rect 19536 30666 19564 31350
rect 19524 30660 19576 30666
rect 19524 30602 19576 30608
rect 19432 30592 19484 30598
rect 19432 30534 19484 30540
rect 19984 30592 20036 30598
rect 19984 30534 20036 30540
rect 19574 30492 19882 30512
rect 19574 30490 19580 30492
rect 19636 30490 19660 30492
rect 19716 30490 19740 30492
rect 19796 30490 19820 30492
rect 19876 30490 19882 30492
rect 19636 30438 19638 30490
rect 19818 30438 19820 30490
rect 19574 30436 19580 30438
rect 19636 30436 19660 30438
rect 19716 30436 19740 30438
rect 19796 30436 19820 30438
rect 19876 30436 19882 30438
rect 19574 30416 19882 30436
rect 19996 30326 20024 30534
rect 19984 30320 20036 30326
rect 19984 30262 20036 30268
rect 19800 30184 19852 30190
rect 19800 30126 19852 30132
rect 19064 29776 19116 29782
rect 19064 29718 19116 29724
rect 19156 29776 19208 29782
rect 19156 29718 19208 29724
rect 18788 28756 18840 28762
rect 18788 28698 18840 28704
rect 18604 28552 18656 28558
rect 18604 28494 18656 28500
rect 18512 25152 18564 25158
rect 18512 25094 18564 25100
rect 18328 24744 18380 24750
rect 18328 24686 18380 24692
rect 18340 23746 18368 24686
rect 18512 24676 18564 24682
rect 18512 24618 18564 24624
rect 18524 24206 18552 24618
rect 18512 24200 18564 24206
rect 18512 24142 18564 24148
rect 18340 23730 18460 23746
rect 18340 23724 18472 23730
rect 18340 23718 18420 23724
rect 18420 23666 18472 23672
rect 18328 23656 18380 23662
rect 18328 23598 18380 23604
rect 18340 23186 18368 23598
rect 18420 23588 18472 23594
rect 18420 23530 18472 23536
rect 18328 23180 18380 23186
rect 18328 23122 18380 23128
rect 18432 21350 18460 23530
rect 18420 21344 18472 21350
rect 18420 21286 18472 21292
rect 18328 20936 18380 20942
rect 18328 20878 18380 20884
rect 18236 20596 18288 20602
rect 18236 20538 18288 20544
rect 18144 20324 18196 20330
rect 18144 20266 18196 20272
rect 18248 19718 18276 20538
rect 18340 20534 18368 20878
rect 18432 20806 18460 21286
rect 18420 20800 18472 20806
rect 18420 20742 18472 20748
rect 18328 20528 18380 20534
rect 18328 20470 18380 20476
rect 18432 20398 18460 20742
rect 18420 20392 18472 20398
rect 18420 20334 18472 20340
rect 18328 20256 18380 20262
rect 18328 20198 18380 20204
rect 18236 19712 18288 19718
rect 18236 19654 18288 19660
rect 18052 19440 18104 19446
rect 18340 19394 18368 20198
rect 18524 19446 18552 24142
rect 18616 22094 18644 28494
rect 18880 27328 18932 27334
rect 18880 27270 18932 27276
rect 18696 27056 18748 27062
rect 18696 26998 18748 27004
rect 18708 26586 18736 26998
rect 18696 26580 18748 26586
rect 18696 26522 18748 26528
rect 18696 26376 18748 26382
rect 18694 26344 18696 26353
rect 18748 26344 18750 26353
rect 18694 26279 18750 26288
rect 18696 25220 18748 25226
rect 18696 25162 18748 25168
rect 18708 23066 18736 25162
rect 18892 23338 18920 27270
rect 19076 27130 19104 29718
rect 19168 29238 19196 29718
rect 19432 29708 19484 29714
rect 19432 29650 19484 29656
rect 19444 29238 19472 29650
rect 19812 29578 19840 30126
rect 19996 29850 20024 30262
rect 19984 29844 20036 29850
rect 19984 29786 20036 29792
rect 19800 29572 19852 29578
rect 19800 29514 19852 29520
rect 19574 29404 19882 29424
rect 19574 29402 19580 29404
rect 19636 29402 19660 29404
rect 19716 29402 19740 29404
rect 19796 29402 19820 29404
rect 19876 29402 19882 29404
rect 19636 29350 19638 29402
rect 19818 29350 19820 29402
rect 19574 29348 19580 29350
rect 19636 29348 19660 29350
rect 19716 29348 19740 29350
rect 19796 29348 19820 29350
rect 19876 29348 19882 29350
rect 19574 29328 19882 29348
rect 19156 29232 19208 29238
rect 19156 29174 19208 29180
rect 19432 29232 19484 29238
rect 19432 29174 19484 29180
rect 19248 29164 19300 29170
rect 19248 29106 19300 29112
rect 19260 28150 19288 29106
rect 19338 29064 19394 29073
rect 19338 28999 19340 29008
rect 19392 28999 19394 29008
rect 19340 28970 19392 28976
rect 19340 28552 19392 28558
rect 19340 28494 19392 28500
rect 19248 28144 19300 28150
rect 19248 28086 19300 28092
rect 19352 27441 19380 28494
rect 19432 28484 19484 28490
rect 19432 28426 19484 28432
rect 19338 27432 19394 27441
rect 19338 27367 19394 27376
rect 19248 27328 19300 27334
rect 19248 27270 19300 27276
rect 19064 27124 19116 27130
rect 19064 27066 19116 27072
rect 19076 26586 19104 27066
rect 19260 26858 19288 27270
rect 19248 26852 19300 26858
rect 19248 26794 19300 26800
rect 19064 26580 19116 26586
rect 19064 26522 19116 26528
rect 19076 26042 19104 26522
rect 19260 26330 19288 26794
rect 19340 26376 19392 26382
rect 19260 26324 19340 26330
rect 19260 26318 19392 26324
rect 19260 26302 19380 26318
rect 19064 26036 19116 26042
rect 19064 25978 19116 25984
rect 19340 24744 19392 24750
rect 19340 24686 19392 24692
rect 19064 24268 19116 24274
rect 19064 24210 19116 24216
rect 18972 23724 19024 23730
rect 18972 23666 19024 23672
rect 18984 23526 19012 23666
rect 18972 23520 19024 23526
rect 18972 23462 19024 23468
rect 18892 23310 19012 23338
rect 18708 23038 18828 23066
rect 18616 22066 18736 22094
rect 18708 21622 18736 22066
rect 18696 21616 18748 21622
rect 18696 21558 18748 21564
rect 18604 21344 18656 21350
rect 18604 21286 18656 21292
rect 18616 21010 18644 21286
rect 18604 21004 18656 21010
rect 18604 20946 18656 20952
rect 18604 20460 18656 20466
rect 18604 20402 18656 20408
rect 18616 19514 18644 20402
rect 18696 19848 18748 19854
rect 18696 19790 18748 19796
rect 18604 19508 18656 19514
rect 18604 19450 18656 19456
rect 18052 19382 18104 19388
rect 17776 19372 17828 19378
rect 17776 19314 17828 19320
rect 16764 19304 16816 19310
rect 16764 19246 16816 19252
rect 17788 18698 17816 19314
rect 18064 18970 18092 19382
rect 18248 19378 18368 19394
rect 18512 19440 18564 19446
rect 18512 19382 18564 19388
rect 18236 19372 18368 19378
rect 18288 19366 18368 19372
rect 18236 19314 18288 19320
rect 18144 19168 18196 19174
rect 18144 19110 18196 19116
rect 17868 18964 17920 18970
rect 17868 18906 17920 18912
rect 18052 18964 18104 18970
rect 18052 18906 18104 18912
rect 17880 18766 17908 18906
rect 17868 18760 17920 18766
rect 17868 18702 17920 18708
rect 16948 18692 17000 18698
rect 16948 18634 17000 18640
rect 17776 18692 17828 18698
rect 17776 18634 17828 18640
rect 16672 17740 16724 17746
rect 16672 17682 16724 17688
rect 16580 17332 16632 17338
rect 16580 17274 16632 17280
rect 16684 16590 16712 17682
rect 16960 17542 16988 18634
rect 17960 18624 18012 18630
rect 17960 18566 18012 18572
rect 17972 18290 18000 18566
rect 18064 18358 18092 18906
rect 18156 18630 18184 19110
rect 18144 18624 18196 18630
rect 18144 18566 18196 18572
rect 18248 18426 18276 19314
rect 18236 18420 18288 18426
rect 18236 18362 18288 18368
rect 18420 18420 18472 18426
rect 18420 18362 18472 18368
rect 18052 18352 18104 18358
rect 18052 18294 18104 18300
rect 17960 18284 18012 18290
rect 17960 18226 18012 18232
rect 18248 17610 18276 18362
rect 18328 18284 18380 18290
rect 18328 18226 18380 18232
rect 18236 17604 18288 17610
rect 18236 17546 18288 17552
rect 18340 17542 18368 18226
rect 16948 17536 17000 17542
rect 16948 17478 17000 17484
rect 18328 17536 18380 17542
rect 18328 17478 18380 17484
rect 16672 16584 16724 16590
rect 16672 16526 16724 16532
rect 16580 15496 16632 15502
rect 16684 15484 16712 16526
rect 16856 15904 16908 15910
rect 16856 15846 16908 15852
rect 16632 15456 16712 15484
rect 16580 15438 16632 15444
rect 16764 15428 16816 15434
rect 16868 15416 16896 15846
rect 16960 15502 16988 17478
rect 17960 17060 18012 17066
rect 17960 17002 18012 17008
rect 17972 16182 18000 17002
rect 17316 16176 17368 16182
rect 17316 16118 17368 16124
rect 17960 16176 18012 16182
rect 17960 16118 18012 16124
rect 16948 15496 17000 15502
rect 16948 15438 17000 15444
rect 16816 15388 16896 15416
rect 16764 15370 16816 15376
rect 16408 15286 16528 15314
rect 15844 14884 15896 14890
rect 15844 14826 15896 14832
rect 15936 14884 15988 14890
rect 15936 14826 15988 14832
rect 15856 14618 15884 14826
rect 15844 14612 15896 14618
rect 15844 14554 15896 14560
rect 15948 14414 15976 14826
rect 16212 14612 16264 14618
rect 16212 14554 16264 14560
rect 15936 14408 15988 14414
rect 15936 14350 15988 14356
rect 15752 14000 15804 14006
rect 15752 13942 15804 13948
rect 15842 13968 15898 13977
rect 15660 13524 15712 13530
rect 15660 13466 15712 13472
rect 15384 13388 15436 13394
rect 15384 13330 15436 13336
rect 15108 12980 15160 12986
rect 15108 12922 15160 12928
rect 15120 12238 15148 12922
rect 15108 12232 15160 12238
rect 15108 12174 15160 12180
rect 15396 11762 15424 13330
rect 15672 12918 15700 13466
rect 15660 12912 15712 12918
rect 15660 12854 15712 12860
rect 15568 12232 15620 12238
rect 15568 12174 15620 12180
rect 15384 11756 15436 11762
rect 15384 11698 15436 11704
rect 15108 11620 15160 11626
rect 15108 11562 15160 11568
rect 15120 11150 15148 11562
rect 15108 11144 15160 11150
rect 15108 11086 15160 11092
rect 15120 10742 15148 11086
rect 15200 11076 15252 11082
rect 15200 11018 15252 11024
rect 15212 10810 15240 11018
rect 15200 10804 15252 10810
rect 15200 10746 15252 10752
rect 15108 10736 15160 10742
rect 15108 10678 15160 10684
rect 15120 10062 15148 10678
rect 15108 10056 15160 10062
rect 15108 9998 15160 10004
rect 15580 8498 15608 12174
rect 15764 12170 15792 13942
rect 15842 13903 15844 13912
rect 15896 13903 15898 13912
rect 15844 13874 15896 13880
rect 15856 12850 15884 13874
rect 15948 13258 15976 14350
rect 16028 14340 16080 14346
rect 16028 14282 16080 14288
rect 16040 13326 16068 14282
rect 16224 14006 16252 14554
rect 16212 14000 16264 14006
rect 16304 14000 16356 14006
rect 16212 13942 16264 13948
rect 16302 13968 16304 13977
rect 16356 13968 16358 13977
rect 16302 13903 16358 13912
rect 16120 13728 16172 13734
rect 16120 13670 16172 13676
rect 16028 13320 16080 13326
rect 16028 13262 16080 13268
rect 15936 13252 15988 13258
rect 15936 13194 15988 13200
rect 15844 12844 15896 12850
rect 15844 12786 15896 12792
rect 16040 12782 16068 13262
rect 16132 12918 16160 13670
rect 16304 13252 16356 13258
rect 16304 13194 16356 13200
rect 16120 12912 16172 12918
rect 16120 12854 16172 12860
rect 16028 12776 16080 12782
rect 16028 12718 16080 12724
rect 15752 12164 15804 12170
rect 15752 12106 15804 12112
rect 16212 12164 16264 12170
rect 16212 12106 16264 12112
rect 15660 12096 15712 12102
rect 15660 12038 15712 12044
rect 15672 11762 15700 12038
rect 15660 11756 15712 11762
rect 15660 11698 15712 11704
rect 16120 11688 16172 11694
rect 16120 11630 16172 11636
rect 15844 11552 15896 11558
rect 15844 11494 15896 11500
rect 15856 11150 15884 11494
rect 16132 11150 16160 11630
rect 15844 11144 15896 11150
rect 15844 11086 15896 11092
rect 16120 11144 16172 11150
rect 16120 11086 16172 11092
rect 16132 10810 16160 11086
rect 16224 11064 16252 12106
rect 16316 11830 16344 13194
rect 16304 11824 16356 11830
rect 16304 11766 16356 11772
rect 16408 11218 16436 15286
rect 16868 14958 16896 15388
rect 16856 14952 16908 14958
rect 16854 14920 16856 14929
rect 16908 14920 16910 14929
rect 16854 14855 16910 14864
rect 16672 14408 16724 14414
rect 16960 14396 16988 15438
rect 17224 14816 17276 14822
rect 17224 14758 17276 14764
rect 17236 14414 17264 14758
rect 16724 14368 16988 14396
rect 17224 14408 17276 14414
rect 16672 14350 16724 14356
rect 17224 14350 17276 14356
rect 16488 14068 16540 14074
rect 16488 14010 16540 14016
rect 16500 12753 16528 14010
rect 16684 13938 16712 14350
rect 16672 13932 16724 13938
rect 16672 13874 16724 13880
rect 16948 13864 17000 13870
rect 16948 13806 17000 13812
rect 16960 13326 16988 13806
rect 16948 13320 17000 13326
rect 16948 13262 17000 13268
rect 16672 13184 16724 13190
rect 16672 13126 16724 13132
rect 16684 12850 16712 13126
rect 16672 12844 16724 12850
rect 16672 12786 16724 12792
rect 17040 12776 17092 12782
rect 16486 12744 16542 12753
rect 17040 12718 17092 12724
rect 16486 12679 16542 12688
rect 17052 12238 17080 12718
rect 17132 12436 17184 12442
rect 17132 12378 17184 12384
rect 17040 12232 17092 12238
rect 17040 12174 17092 12180
rect 17144 12170 17172 12378
rect 17222 12336 17278 12345
rect 17222 12271 17278 12280
rect 16764 12164 16816 12170
rect 16764 12106 16816 12112
rect 17132 12164 17184 12170
rect 17132 12106 17184 12112
rect 16488 12096 16540 12102
rect 16488 12038 16540 12044
rect 16500 11762 16528 12038
rect 16488 11756 16540 11762
rect 16488 11698 16540 11704
rect 16672 11756 16724 11762
rect 16672 11698 16724 11704
rect 16396 11212 16448 11218
rect 16396 11154 16448 11160
rect 16684 11150 16712 11698
rect 16776 11286 16804 12106
rect 17144 11762 17172 12106
rect 16948 11756 17000 11762
rect 16868 11716 16948 11744
rect 16764 11280 16816 11286
rect 16764 11222 16816 11228
rect 16672 11144 16724 11150
rect 16672 11086 16724 11092
rect 16304 11076 16356 11082
rect 16224 11036 16304 11064
rect 16304 11018 16356 11024
rect 16120 10804 16172 10810
rect 16120 10746 16172 10752
rect 15752 10464 15804 10470
rect 15752 10406 15804 10412
rect 15764 9926 15792 10406
rect 16868 9926 16896 11716
rect 16948 11698 17000 11704
rect 17132 11756 17184 11762
rect 17132 11698 17184 11704
rect 16948 11008 17000 11014
rect 16948 10950 17000 10956
rect 16960 10062 16988 10950
rect 17040 10804 17092 10810
rect 17040 10746 17092 10752
rect 17052 10062 17080 10746
rect 16948 10056 17000 10062
rect 16948 9998 17000 10004
rect 17040 10056 17092 10062
rect 17040 9998 17092 10004
rect 15752 9920 15804 9926
rect 15752 9862 15804 9868
rect 16580 9920 16632 9926
rect 16580 9862 16632 9868
rect 16856 9920 16908 9926
rect 16856 9862 16908 9868
rect 15764 9722 15792 9862
rect 15752 9716 15804 9722
rect 15752 9658 15804 9664
rect 15844 9376 15896 9382
rect 15844 9318 15896 9324
rect 15936 9376 15988 9382
rect 15936 9318 15988 9324
rect 15856 8906 15884 9318
rect 15948 9042 15976 9318
rect 15936 9036 15988 9042
rect 15936 8978 15988 8984
rect 15844 8900 15896 8906
rect 15844 8842 15896 8848
rect 15568 8492 15620 8498
rect 15568 8434 15620 8440
rect 15016 8288 15068 8294
rect 15016 8230 15068 8236
rect 14464 7880 14516 7886
rect 14464 7822 14516 7828
rect 14924 7880 14976 7886
rect 14924 7822 14976 7828
rect 14200 7410 14320 7426
rect 14188 7404 14320 7410
rect 14240 7398 14320 7404
rect 14188 7346 14240 7352
rect 14188 7200 14240 7206
rect 14188 7142 14240 7148
rect 14200 6934 14228 7142
rect 14188 6928 14240 6934
rect 14188 6870 14240 6876
rect 14292 6798 14320 7398
rect 14372 7336 14424 7342
rect 14372 7278 14424 7284
rect 14384 7206 14412 7278
rect 14476 7274 14504 7822
rect 14936 7478 14964 7822
rect 14924 7472 14976 7478
rect 14924 7414 14976 7420
rect 14464 7268 14516 7274
rect 14464 7210 14516 7216
rect 14372 7200 14424 7206
rect 14372 7142 14424 7148
rect 14384 6866 14412 7142
rect 16592 6866 16620 9862
rect 16868 9674 16896 9862
rect 16868 9646 16988 9674
rect 17052 9654 17080 9998
rect 16960 9586 16988 9646
rect 17040 9648 17092 9654
rect 17040 9590 17092 9596
rect 16948 9580 17000 9586
rect 16948 9522 17000 9528
rect 17144 8566 17172 11698
rect 17236 8974 17264 12271
rect 17328 11898 17356 16118
rect 17592 15360 17644 15366
rect 17592 15302 17644 15308
rect 17604 15026 17632 15302
rect 17972 15094 18000 16118
rect 17960 15088 18012 15094
rect 17960 15030 18012 15036
rect 17592 15020 17644 15026
rect 17592 14962 17644 14968
rect 17408 14952 17460 14958
rect 17408 14894 17460 14900
rect 17682 14920 17738 14929
rect 17420 13326 17448 14894
rect 17682 14855 17684 14864
rect 17736 14855 17738 14864
rect 17684 14826 17736 14832
rect 17776 14408 17828 14414
rect 17776 14350 17828 14356
rect 17500 14340 17552 14346
rect 17500 14282 17552 14288
rect 17512 13530 17540 14282
rect 17500 13524 17552 13530
rect 17500 13466 17552 13472
rect 17408 13320 17460 13326
rect 17408 13262 17460 13268
rect 17788 13258 17816 14350
rect 17868 13864 17920 13870
rect 17868 13806 17920 13812
rect 17880 13326 17908 13806
rect 17868 13320 17920 13326
rect 17868 13262 17920 13268
rect 17776 13252 17828 13258
rect 17776 13194 17828 13200
rect 17776 12912 17828 12918
rect 17776 12854 17828 12860
rect 17788 12170 17816 12854
rect 17776 12164 17828 12170
rect 17776 12106 17828 12112
rect 17592 12096 17644 12102
rect 17592 12038 17644 12044
rect 17316 11892 17368 11898
rect 17316 11834 17368 11840
rect 17604 11218 17632 12038
rect 17592 11212 17644 11218
rect 17592 11154 17644 11160
rect 17880 11150 17908 13262
rect 17972 12850 18000 15030
rect 18236 13456 18288 13462
rect 18236 13398 18288 13404
rect 17960 12844 18012 12850
rect 17960 12786 18012 12792
rect 17868 11144 17920 11150
rect 17868 11086 17920 11092
rect 17774 9208 17830 9217
rect 17774 9143 17830 9152
rect 17498 9072 17554 9081
rect 17498 9007 17500 9016
rect 17552 9007 17554 9016
rect 17500 8978 17552 8984
rect 17224 8968 17276 8974
rect 17224 8910 17276 8916
rect 17684 8832 17736 8838
rect 17684 8774 17736 8780
rect 17132 8560 17184 8566
rect 17132 8502 17184 8508
rect 17408 7948 17460 7954
rect 17408 7890 17460 7896
rect 17420 7410 17448 7890
rect 17696 7410 17724 8774
rect 17788 8634 17816 9143
rect 18248 8634 18276 13398
rect 17776 8628 17828 8634
rect 17776 8570 17828 8576
rect 18236 8628 18288 8634
rect 18236 8570 18288 8576
rect 17788 7954 17816 8570
rect 17776 7948 17828 7954
rect 17776 7890 17828 7896
rect 18248 7886 18276 8570
rect 18236 7880 18288 7886
rect 18236 7822 18288 7828
rect 18052 7744 18104 7750
rect 18052 7686 18104 7692
rect 17408 7404 17460 7410
rect 17408 7346 17460 7352
rect 17684 7404 17736 7410
rect 17684 7346 17736 7352
rect 16856 7200 16908 7206
rect 16856 7142 16908 7148
rect 14372 6860 14424 6866
rect 14372 6802 14424 6808
rect 16580 6860 16632 6866
rect 16580 6802 16632 6808
rect 16764 6860 16816 6866
rect 16764 6802 16816 6808
rect 14280 6792 14332 6798
rect 11624 6390 11652 6734
rect 14108 6718 14228 6746
rect 14280 6734 14332 6740
rect 12808 6452 12860 6458
rect 12808 6394 12860 6400
rect 11612 6384 11664 6390
rect 11612 6326 11664 6332
rect 12820 5778 12848 6394
rect 14004 6384 14056 6390
rect 14004 6326 14056 6332
rect 13544 6316 13596 6322
rect 13544 6258 13596 6264
rect 13636 6316 13688 6322
rect 13636 6258 13688 6264
rect 13452 6112 13504 6118
rect 13452 6054 13504 6060
rect 10508 5772 10560 5778
rect 10508 5714 10560 5720
rect 12808 5772 12860 5778
rect 12808 5714 12860 5720
rect 10416 5704 10468 5710
rect 10416 5646 10468 5652
rect 10336 5494 10456 5522
rect 10324 5024 10376 5030
rect 10324 4966 10376 4972
rect 10232 4684 10284 4690
rect 10232 4626 10284 4632
rect 10336 4622 10364 4966
rect 10324 4616 10376 4622
rect 10324 4558 10376 4564
rect 10324 4072 10376 4078
rect 10324 4014 10376 4020
rect 9772 3732 9824 3738
rect 9772 3674 9824 3680
rect 10048 3732 10100 3738
rect 10048 3674 10100 3680
rect 10060 3466 10088 3674
rect 10048 3460 10100 3466
rect 10048 3402 10100 3408
rect 10140 3188 10192 3194
rect 10140 3130 10192 3136
rect 10152 3058 10180 3130
rect 10336 3058 10364 4014
rect 10140 3052 10192 3058
rect 10140 2994 10192 3000
rect 10324 3052 10376 3058
rect 10324 2994 10376 3000
rect 9680 2916 9732 2922
rect 9680 2858 9732 2864
rect 8760 2576 8812 2582
rect 8760 2518 8812 2524
rect 10152 2514 10180 2994
rect 10428 2774 10456 5494
rect 13464 5234 13492 6054
rect 13556 5642 13584 6258
rect 13648 5778 13676 6258
rect 13636 5772 13688 5778
rect 13636 5714 13688 5720
rect 14016 5710 14044 6326
rect 14004 5704 14056 5710
rect 14004 5646 14056 5652
rect 13544 5636 13596 5642
rect 13544 5578 13596 5584
rect 13452 5228 13504 5234
rect 13452 5170 13504 5176
rect 11060 4616 11112 4622
rect 11060 4558 11112 4564
rect 11072 4010 11100 4558
rect 11152 4480 11204 4486
rect 11152 4422 11204 4428
rect 12716 4480 12768 4486
rect 12716 4422 12768 4428
rect 11164 4214 11192 4422
rect 12728 4214 12756 4422
rect 11152 4208 11204 4214
rect 11152 4150 11204 4156
rect 12716 4208 12768 4214
rect 12716 4150 12768 4156
rect 11796 4140 11848 4146
rect 11796 4082 11848 4088
rect 11336 4072 11388 4078
rect 11336 4014 11388 4020
rect 11060 4004 11112 4010
rect 11060 3946 11112 3952
rect 10600 3528 10652 3534
rect 10600 3470 10652 3476
rect 10612 2990 10640 3470
rect 11072 3398 11100 3946
rect 11348 3534 11376 4014
rect 11808 3942 11836 4082
rect 11888 4072 11940 4078
rect 11888 4014 11940 4020
rect 11980 4072 12032 4078
rect 11980 4014 12032 4020
rect 12900 4072 12952 4078
rect 12900 4014 12952 4020
rect 11796 3936 11848 3942
rect 11796 3878 11848 3884
rect 11336 3528 11388 3534
rect 11336 3470 11388 3476
rect 11428 3528 11480 3534
rect 11428 3470 11480 3476
rect 11060 3392 11112 3398
rect 11440 3346 11468 3470
rect 11060 3334 11112 3340
rect 11348 3318 11468 3346
rect 11520 3392 11572 3398
rect 11520 3334 11572 3340
rect 11348 3194 11376 3318
rect 11532 3194 11560 3334
rect 11336 3188 11388 3194
rect 11336 3130 11388 3136
rect 11520 3188 11572 3194
rect 11520 3130 11572 3136
rect 11808 2990 11836 3878
rect 11900 3602 11928 4014
rect 11888 3596 11940 3602
rect 11888 3538 11940 3544
rect 11992 3466 12020 4014
rect 12440 3936 12492 3942
rect 12440 3878 12492 3884
rect 12452 3738 12480 3878
rect 12912 3738 12940 4014
rect 13452 3936 13504 3942
rect 13452 3878 13504 3884
rect 12440 3732 12492 3738
rect 12440 3674 12492 3680
rect 12900 3732 12952 3738
rect 12900 3674 12952 3680
rect 13464 3534 13492 3878
rect 13452 3528 13504 3534
rect 13452 3470 13504 3476
rect 11980 3460 12032 3466
rect 11980 3402 12032 3408
rect 11992 3058 12020 3402
rect 14096 3392 14148 3398
rect 14096 3334 14148 3340
rect 14108 3126 14136 3334
rect 14096 3120 14148 3126
rect 14096 3062 14148 3068
rect 11980 3052 12032 3058
rect 11980 2994 12032 3000
rect 10600 2984 10652 2990
rect 10600 2926 10652 2932
rect 11796 2984 11848 2990
rect 11796 2926 11848 2932
rect 13452 2916 13504 2922
rect 13452 2858 13504 2864
rect 10428 2746 10548 2774
rect 10520 2514 10548 2746
rect 10140 2508 10192 2514
rect 10140 2450 10192 2456
rect 10508 2508 10560 2514
rect 10508 2450 10560 2456
rect 13464 2446 13492 2858
rect 7748 2440 7800 2446
rect 7748 2382 7800 2388
rect 8484 2440 8536 2446
rect 8484 2382 8536 2388
rect 9680 2440 9732 2446
rect 9680 2382 9732 2388
rect 13452 2440 13504 2446
rect 13452 2382 13504 2388
rect 5172 2100 5224 2106
rect 5172 2042 5224 2048
rect 7760 800 7788 2382
rect 9692 800 9720 2382
rect 11612 2304 11664 2310
rect 11612 2246 11664 2252
rect 12532 2304 12584 2310
rect 12532 2246 12584 2252
rect 13544 2304 13596 2310
rect 13544 2246 13596 2252
rect 11624 800 11652 2246
rect 12544 2038 12572 2246
rect 12532 2032 12584 2038
rect 12532 1974 12584 1980
rect 13556 800 13584 2246
rect 14200 1902 14228 6718
rect 16592 6322 16620 6802
rect 16580 6316 16632 6322
rect 16580 6258 16632 6264
rect 16776 6118 16804 6802
rect 16868 6798 16896 7142
rect 17420 7002 17448 7346
rect 18064 7274 18092 7686
rect 18052 7268 18104 7274
rect 18052 7210 18104 7216
rect 18340 7002 18368 17478
rect 18432 14550 18460 18362
rect 18524 17678 18552 19382
rect 18616 17678 18644 19450
rect 18708 19378 18736 19790
rect 18800 19496 18828 23038
rect 18880 19508 18932 19514
rect 18800 19468 18880 19496
rect 18880 19450 18932 19456
rect 18696 19372 18748 19378
rect 18696 19314 18748 19320
rect 18880 18692 18932 18698
rect 18880 18634 18932 18640
rect 18892 18222 18920 18634
rect 18880 18216 18932 18222
rect 18880 18158 18932 18164
rect 18512 17672 18564 17678
rect 18512 17614 18564 17620
rect 18604 17672 18656 17678
rect 18604 17614 18656 17620
rect 18880 15904 18932 15910
rect 18880 15846 18932 15852
rect 18420 14544 18472 14550
rect 18420 14486 18472 14492
rect 18892 12850 18920 15846
rect 18880 12844 18932 12850
rect 18880 12786 18932 12792
rect 18512 12776 18564 12782
rect 18512 12718 18564 12724
rect 18524 12102 18552 12718
rect 18892 12646 18920 12786
rect 18880 12640 18932 12646
rect 18880 12582 18932 12588
rect 18788 12164 18840 12170
rect 18788 12106 18840 12112
rect 18512 12096 18564 12102
rect 18512 12038 18564 12044
rect 18524 11626 18552 12038
rect 18800 11898 18828 12106
rect 18788 11892 18840 11898
rect 18788 11834 18840 11840
rect 18512 11620 18564 11626
rect 18512 11562 18564 11568
rect 18696 10464 18748 10470
rect 18696 10406 18748 10412
rect 18708 10130 18736 10406
rect 18696 10124 18748 10130
rect 18696 10066 18748 10072
rect 17408 6996 17460 7002
rect 17408 6938 17460 6944
rect 18328 6996 18380 7002
rect 18328 6938 18380 6944
rect 16856 6792 16908 6798
rect 16856 6734 16908 6740
rect 16868 6322 16896 6734
rect 17224 6656 17276 6662
rect 17224 6598 17276 6604
rect 17236 6322 17264 6598
rect 16856 6316 16908 6322
rect 16856 6258 16908 6264
rect 17224 6316 17276 6322
rect 17224 6258 17276 6264
rect 17960 6316 18012 6322
rect 17960 6258 18012 6264
rect 16764 6112 16816 6118
rect 16764 6054 16816 6060
rect 17236 5778 17264 6258
rect 17592 6112 17644 6118
rect 17592 6054 17644 6060
rect 17684 6112 17736 6118
rect 17684 6054 17736 6060
rect 17224 5772 17276 5778
rect 17224 5714 17276 5720
rect 17604 5710 17632 6054
rect 16580 5704 16632 5710
rect 16580 5646 16632 5652
rect 17592 5704 17644 5710
rect 17592 5646 17644 5652
rect 14464 5568 14516 5574
rect 14464 5510 14516 5516
rect 14476 5234 14504 5510
rect 14464 5228 14516 5234
rect 14464 5170 14516 5176
rect 16592 5098 16620 5646
rect 17696 5098 17724 6054
rect 17972 5846 18000 6258
rect 17960 5840 18012 5846
rect 17960 5782 18012 5788
rect 16580 5092 16632 5098
rect 16580 5034 16632 5040
rect 17684 5092 17736 5098
rect 17684 5034 17736 5040
rect 16672 5024 16724 5030
rect 16672 4966 16724 4972
rect 17592 5024 17644 5030
rect 17592 4966 17644 4972
rect 15844 4820 15896 4826
rect 15844 4762 15896 4768
rect 16028 4820 16080 4826
rect 16028 4762 16080 4768
rect 15856 4214 15884 4762
rect 16040 4282 16068 4762
rect 16684 4554 16712 4966
rect 17604 4622 17632 4966
rect 17972 4826 18000 5782
rect 17960 4820 18012 4826
rect 17960 4762 18012 4768
rect 17592 4616 17644 4622
rect 17592 4558 17644 4564
rect 16672 4548 16724 4554
rect 16672 4490 16724 4496
rect 16028 4276 16080 4282
rect 16028 4218 16080 4224
rect 16212 4276 16264 4282
rect 16212 4218 16264 4224
rect 15752 4208 15804 4214
rect 15752 4150 15804 4156
rect 15844 4208 15896 4214
rect 16224 4162 16252 4218
rect 15844 4150 15896 4156
rect 15764 4060 15792 4150
rect 16132 4134 16252 4162
rect 16684 4146 16712 4490
rect 16948 4480 17000 4486
rect 16948 4422 17000 4428
rect 16672 4140 16724 4146
rect 16132 4060 16160 4134
rect 16672 4082 16724 4088
rect 15764 4032 16160 4060
rect 16672 4004 16724 4010
rect 16672 3946 16724 3952
rect 14924 3936 14976 3942
rect 14924 3878 14976 3884
rect 14936 3738 14964 3878
rect 14924 3732 14976 3738
rect 14924 3674 14976 3680
rect 14280 3664 14332 3670
rect 14280 3606 14332 3612
rect 14292 3398 14320 3606
rect 14936 3534 14964 3674
rect 15016 3664 15068 3670
rect 15016 3606 15068 3612
rect 14924 3528 14976 3534
rect 14924 3470 14976 3476
rect 14280 3392 14332 3398
rect 14280 3334 14332 3340
rect 15028 3126 15056 3606
rect 16684 3534 16712 3946
rect 16960 3942 16988 4422
rect 17684 4072 17736 4078
rect 17684 4014 17736 4020
rect 16948 3936 17000 3942
rect 16948 3878 17000 3884
rect 15108 3528 15160 3534
rect 15108 3470 15160 3476
rect 16672 3528 16724 3534
rect 16672 3470 16724 3476
rect 15120 3194 15148 3470
rect 15108 3188 15160 3194
rect 15108 3130 15160 3136
rect 15016 3120 15068 3126
rect 15016 3062 15068 3068
rect 16960 2990 16988 3878
rect 17696 3534 17724 4014
rect 18052 3596 18104 3602
rect 18052 3538 18104 3544
rect 17316 3528 17368 3534
rect 17316 3470 17368 3476
rect 17408 3528 17460 3534
rect 17408 3470 17460 3476
rect 17684 3528 17736 3534
rect 17684 3470 17736 3476
rect 17328 3058 17356 3470
rect 17316 3052 17368 3058
rect 17316 2994 17368 3000
rect 16948 2984 17000 2990
rect 16948 2926 17000 2932
rect 17420 2854 17448 3470
rect 17960 3392 18012 3398
rect 17960 3334 18012 3340
rect 17972 2990 18000 3334
rect 18064 3097 18092 3538
rect 18050 3088 18106 3097
rect 18050 3023 18052 3032
rect 18104 3023 18106 3032
rect 18052 2994 18104 3000
rect 17960 2984 18012 2990
rect 17960 2926 18012 2932
rect 17408 2848 17460 2854
rect 17408 2790 17460 2796
rect 18984 2774 19012 23310
rect 19076 21672 19104 24210
rect 19352 23866 19380 24686
rect 19248 23860 19300 23866
rect 19248 23802 19300 23808
rect 19340 23860 19392 23866
rect 19340 23802 19392 23808
rect 19156 22976 19208 22982
rect 19156 22918 19208 22924
rect 19168 22642 19196 22918
rect 19260 22778 19288 23802
rect 19444 23730 19472 28426
rect 20076 28416 20128 28422
rect 20076 28358 20128 28364
rect 19574 28316 19882 28336
rect 19574 28314 19580 28316
rect 19636 28314 19660 28316
rect 19716 28314 19740 28316
rect 19796 28314 19820 28316
rect 19876 28314 19882 28316
rect 19636 28262 19638 28314
rect 19818 28262 19820 28314
rect 19574 28260 19580 28262
rect 19636 28260 19660 28262
rect 19716 28260 19740 28262
rect 19796 28260 19820 28262
rect 19876 28260 19882 28262
rect 19574 28240 19882 28260
rect 19574 27228 19882 27248
rect 19574 27226 19580 27228
rect 19636 27226 19660 27228
rect 19716 27226 19740 27228
rect 19796 27226 19820 27228
rect 19876 27226 19882 27228
rect 19636 27174 19638 27226
rect 19818 27174 19820 27226
rect 19574 27172 19580 27174
rect 19636 27172 19660 27174
rect 19716 27172 19740 27174
rect 19796 27172 19820 27174
rect 19876 27172 19882 27174
rect 19574 27152 19882 27172
rect 19984 27124 20036 27130
rect 19984 27066 20036 27072
rect 19996 26586 20024 27066
rect 19616 26580 19668 26586
rect 19616 26522 19668 26528
rect 19984 26580 20036 26586
rect 19984 26522 20036 26528
rect 19628 26314 19656 26522
rect 19708 26376 19760 26382
rect 19706 26344 19708 26353
rect 19760 26344 19762 26353
rect 19616 26308 19668 26314
rect 19706 26279 19762 26288
rect 19616 26250 19668 26256
rect 19574 26140 19882 26160
rect 19574 26138 19580 26140
rect 19636 26138 19660 26140
rect 19716 26138 19740 26140
rect 19796 26138 19820 26140
rect 19876 26138 19882 26140
rect 19636 26086 19638 26138
rect 19818 26086 19820 26138
rect 19574 26084 19580 26086
rect 19636 26084 19660 26086
rect 19716 26084 19740 26086
rect 19796 26084 19820 26086
rect 19876 26084 19882 26086
rect 19574 26064 19882 26084
rect 19574 25052 19882 25072
rect 19574 25050 19580 25052
rect 19636 25050 19660 25052
rect 19716 25050 19740 25052
rect 19796 25050 19820 25052
rect 19876 25050 19882 25052
rect 19636 24998 19638 25050
rect 19818 24998 19820 25050
rect 19574 24996 19580 24998
rect 19636 24996 19660 24998
rect 19716 24996 19740 24998
rect 19796 24996 19820 24998
rect 19876 24996 19882 24998
rect 19574 24976 19882 24996
rect 20088 24936 20116 28358
rect 20180 27470 20208 31726
rect 21008 30122 21036 31826
rect 20996 30116 21048 30122
rect 20996 30058 21048 30064
rect 21192 29306 21220 32166
rect 22020 31890 22048 32302
rect 22296 32298 22324 32846
rect 22480 32366 22508 33458
rect 23216 32978 23244 33458
rect 23204 32972 23256 32978
rect 23204 32914 23256 32920
rect 24688 32502 24716 33458
rect 24964 33454 24992 34070
rect 25320 33584 25372 33590
rect 25320 33526 25372 33532
rect 24952 33448 25004 33454
rect 24952 33390 25004 33396
rect 24768 32768 24820 32774
rect 24768 32710 24820 32716
rect 24780 32502 24808 32710
rect 24400 32496 24452 32502
rect 24400 32438 24452 32444
rect 24676 32496 24728 32502
rect 24676 32438 24728 32444
rect 24768 32496 24820 32502
rect 24768 32438 24820 32444
rect 24216 32428 24268 32434
rect 24216 32370 24268 32376
rect 22468 32360 22520 32366
rect 22468 32302 22520 32308
rect 22100 32292 22152 32298
rect 22100 32234 22152 32240
rect 22284 32292 22336 32298
rect 22284 32234 22336 32240
rect 22008 31884 22060 31890
rect 22008 31826 22060 31832
rect 22112 30938 22140 32234
rect 22296 31210 22324 32234
rect 24228 31890 24256 32370
rect 24216 31884 24268 31890
rect 24216 31826 24268 31832
rect 24412 31822 24440 32438
rect 24400 31816 24452 31822
rect 24400 31758 24452 31764
rect 22836 31408 22888 31414
rect 22836 31350 22888 31356
rect 22284 31204 22336 31210
rect 22284 31146 22336 31152
rect 22100 30932 22152 30938
rect 22100 30874 22152 30880
rect 22848 30870 22876 31350
rect 22836 30864 22888 30870
rect 22836 30806 22888 30812
rect 22836 30728 22888 30734
rect 22836 30670 22888 30676
rect 23112 30728 23164 30734
rect 23112 30670 23164 30676
rect 22192 30592 22244 30598
rect 22192 30534 22244 30540
rect 22204 30054 22232 30534
rect 22848 30394 22876 30670
rect 23020 30592 23072 30598
rect 23020 30534 23072 30540
rect 22836 30388 22888 30394
rect 22836 30330 22888 30336
rect 22928 30252 22980 30258
rect 22928 30194 22980 30200
rect 22940 30054 22968 30194
rect 22192 30048 22244 30054
rect 22192 29990 22244 29996
rect 22928 30048 22980 30054
rect 22928 29990 22980 29996
rect 22940 29850 22968 29990
rect 23032 29850 23060 30534
rect 23124 30258 23152 30670
rect 24412 30394 24440 31758
rect 24768 30592 24820 30598
rect 24768 30534 24820 30540
rect 24400 30388 24452 30394
rect 24400 30330 24452 30336
rect 23112 30252 23164 30258
rect 23112 30194 23164 30200
rect 22928 29844 22980 29850
rect 22928 29786 22980 29792
rect 23020 29844 23072 29850
rect 23020 29786 23072 29792
rect 22940 29646 22968 29786
rect 23124 29714 23152 30194
rect 24308 30184 24360 30190
rect 24308 30126 24360 30132
rect 23112 29708 23164 29714
rect 23112 29650 23164 29656
rect 22928 29640 22980 29646
rect 22928 29582 22980 29588
rect 22376 29504 22428 29510
rect 22376 29446 22428 29452
rect 21180 29300 21232 29306
rect 21180 29242 21232 29248
rect 21192 28994 21220 29242
rect 21100 28966 21220 28994
rect 21100 28626 21128 28966
rect 21088 28620 21140 28626
rect 21088 28562 21140 28568
rect 22284 28620 22336 28626
rect 22284 28562 22336 28568
rect 22008 28484 22060 28490
rect 22008 28426 22060 28432
rect 22100 28484 22152 28490
rect 22100 28426 22152 28432
rect 22020 28014 22048 28426
rect 22008 28008 22060 28014
rect 22006 27976 22008 27985
rect 22060 27976 22062 27985
rect 22006 27911 22062 27920
rect 22112 27554 22140 28426
rect 22296 28082 22324 28562
rect 22284 28076 22336 28082
rect 22284 28018 22336 28024
rect 22020 27538 22140 27554
rect 22296 27538 22324 28018
rect 20352 27532 20404 27538
rect 20352 27474 20404 27480
rect 22008 27532 22140 27538
rect 22060 27526 22140 27532
rect 22284 27532 22336 27538
rect 22008 27474 22060 27480
rect 22284 27474 22336 27480
rect 20168 27464 20220 27470
rect 20168 27406 20220 27412
rect 20364 26926 20392 27474
rect 20812 27464 20864 27470
rect 20812 27406 20864 27412
rect 20536 26988 20588 26994
rect 20824 26976 20852 27406
rect 20588 26948 20852 26976
rect 20536 26930 20588 26936
rect 20168 26920 20220 26926
rect 20168 26862 20220 26868
rect 20352 26920 20404 26926
rect 20352 26862 20404 26868
rect 20180 25430 20208 26862
rect 20720 26852 20772 26858
rect 20720 26794 20772 26800
rect 20628 26784 20680 26790
rect 20628 26726 20680 26732
rect 20640 26450 20668 26726
rect 20628 26444 20680 26450
rect 20628 26386 20680 26392
rect 20628 26240 20680 26246
rect 20628 26182 20680 26188
rect 20640 26042 20668 26182
rect 20628 26036 20680 26042
rect 20628 25978 20680 25984
rect 20168 25424 20220 25430
rect 20168 25366 20220 25372
rect 19996 24908 20116 24936
rect 19996 24857 20024 24908
rect 20180 24886 20208 25366
rect 20640 25294 20668 25978
rect 20732 25498 20760 26794
rect 20824 26790 20852 26948
rect 22192 26988 22244 26994
rect 22192 26930 22244 26936
rect 21180 26920 21232 26926
rect 21180 26862 21232 26868
rect 21640 26920 21692 26926
rect 21640 26862 21692 26868
rect 20812 26784 20864 26790
rect 20812 26726 20864 26732
rect 20824 26625 20852 26726
rect 20810 26616 20866 26625
rect 20810 26551 20866 26560
rect 21088 26512 21140 26518
rect 21088 26454 21140 26460
rect 21100 26246 21128 26454
rect 21088 26240 21140 26246
rect 21088 26182 21140 26188
rect 21100 25974 21128 26182
rect 21088 25968 21140 25974
rect 21088 25910 21140 25916
rect 20904 25764 20956 25770
rect 20904 25706 20956 25712
rect 20720 25492 20772 25498
rect 20720 25434 20772 25440
rect 20628 25288 20680 25294
rect 20628 25230 20680 25236
rect 20168 24880 20220 24886
rect 19982 24848 20038 24857
rect 20168 24822 20220 24828
rect 20350 24848 20406 24857
rect 19982 24783 20038 24792
rect 20076 24812 20128 24818
rect 20350 24783 20406 24792
rect 20076 24754 20128 24760
rect 20088 24614 20116 24754
rect 20260 24676 20312 24682
rect 20260 24618 20312 24624
rect 20076 24608 20128 24614
rect 20076 24550 20128 24556
rect 20088 24206 20116 24550
rect 20076 24200 20128 24206
rect 20076 24142 20128 24148
rect 20168 24200 20220 24206
rect 20168 24142 20220 24148
rect 19984 24132 20036 24138
rect 19984 24074 20036 24080
rect 19574 23964 19882 23984
rect 19574 23962 19580 23964
rect 19636 23962 19660 23964
rect 19716 23962 19740 23964
rect 19796 23962 19820 23964
rect 19876 23962 19882 23964
rect 19636 23910 19638 23962
rect 19818 23910 19820 23962
rect 19574 23908 19580 23910
rect 19636 23908 19660 23910
rect 19716 23908 19740 23910
rect 19796 23908 19820 23910
rect 19876 23908 19882 23910
rect 19574 23888 19882 23908
rect 19432 23724 19484 23730
rect 19432 23666 19484 23672
rect 19996 23662 20024 24074
rect 20180 24041 20208 24142
rect 20272 24070 20300 24618
rect 20260 24064 20312 24070
rect 20166 24032 20222 24041
rect 20088 23990 20166 24018
rect 19984 23656 20036 23662
rect 19984 23598 20036 23604
rect 19340 23520 19392 23526
rect 19340 23462 19392 23468
rect 19248 22772 19300 22778
rect 19248 22714 19300 22720
rect 19352 22642 19380 23462
rect 19984 23180 20036 23186
rect 19984 23122 20036 23128
rect 19574 22876 19882 22896
rect 19574 22874 19580 22876
rect 19636 22874 19660 22876
rect 19716 22874 19740 22876
rect 19796 22874 19820 22876
rect 19876 22874 19882 22876
rect 19636 22822 19638 22874
rect 19818 22822 19820 22874
rect 19574 22820 19580 22822
rect 19636 22820 19660 22822
rect 19716 22820 19740 22822
rect 19796 22820 19820 22822
rect 19876 22820 19882 22822
rect 19574 22800 19882 22820
rect 19996 22778 20024 23122
rect 20088 23118 20116 23990
rect 20260 24006 20312 24012
rect 20166 23967 20222 23976
rect 20168 23860 20220 23866
rect 20168 23802 20220 23808
rect 20180 23730 20208 23802
rect 20168 23724 20220 23730
rect 20168 23666 20220 23672
rect 20272 23254 20300 24006
rect 20364 23866 20392 24783
rect 20812 24744 20864 24750
rect 20812 24686 20864 24692
rect 20536 24608 20588 24614
rect 20536 24550 20588 24556
rect 20444 24132 20496 24138
rect 20444 24074 20496 24080
rect 20352 23860 20404 23866
rect 20352 23802 20404 23808
rect 20260 23248 20312 23254
rect 20260 23190 20312 23196
rect 20076 23112 20128 23118
rect 20076 23054 20128 23060
rect 20168 23044 20220 23050
rect 20168 22986 20220 22992
rect 20076 22976 20128 22982
rect 20076 22918 20128 22924
rect 19984 22772 20036 22778
rect 19984 22714 20036 22720
rect 19156 22636 19208 22642
rect 19156 22578 19208 22584
rect 19340 22636 19392 22642
rect 19340 22578 19392 22584
rect 19352 21894 19380 22578
rect 19432 22160 19484 22166
rect 19432 22102 19484 22108
rect 19340 21888 19392 21894
rect 19340 21830 19392 21836
rect 19076 21644 19196 21672
rect 19064 21548 19116 21554
rect 19064 21490 19116 21496
rect 19076 20602 19104 21490
rect 19168 20602 19196 21644
rect 19338 21312 19394 21321
rect 19338 21247 19394 21256
rect 19064 20596 19116 20602
rect 19064 20538 19116 20544
rect 19156 20596 19208 20602
rect 19156 20538 19208 20544
rect 19168 20482 19196 20538
rect 19076 20454 19196 20482
rect 19076 15910 19104 20454
rect 19156 20324 19208 20330
rect 19156 20266 19208 20272
rect 19168 19446 19196 20266
rect 19248 19780 19300 19786
rect 19248 19722 19300 19728
rect 19156 19440 19208 19446
rect 19156 19382 19208 19388
rect 19260 18766 19288 19722
rect 19248 18760 19300 18766
rect 19248 18702 19300 18708
rect 19352 16114 19380 21247
rect 19444 20942 19472 22102
rect 19892 22024 19944 22030
rect 19892 21966 19944 21972
rect 19904 21876 19932 21966
rect 19904 21865 20024 21876
rect 19904 21856 20038 21865
rect 19904 21848 19982 21856
rect 19574 21788 19882 21808
rect 19982 21791 20038 21800
rect 19574 21786 19580 21788
rect 19636 21786 19660 21788
rect 19716 21786 19740 21788
rect 19796 21786 19820 21788
rect 19876 21786 19882 21788
rect 19636 21734 19638 21786
rect 19818 21734 19820 21786
rect 19574 21732 19580 21734
rect 19636 21732 19660 21734
rect 19716 21732 19740 21734
rect 19796 21732 19820 21734
rect 19876 21732 19882 21734
rect 19574 21712 19882 21732
rect 20088 21690 20116 22918
rect 20180 21894 20208 22986
rect 20352 22568 20404 22574
rect 20352 22510 20404 22516
rect 20168 21888 20220 21894
rect 20168 21830 20220 21836
rect 20076 21684 20128 21690
rect 20076 21626 20128 21632
rect 19984 21616 20036 21622
rect 19984 21558 20036 21564
rect 19616 21548 19668 21554
rect 19668 21508 19932 21536
rect 19616 21490 19668 21496
rect 19800 21140 19852 21146
rect 19800 21082 19852 21088
rect 19524 21072 19576 21078
rect 19524 21014 19576 21020
rect 19432 20936 19484 20942
rect 19432 20878 19484 20884
rect 19536 20890 19564 21014
rect 19812 20890 19840 21082
rect 19904 20942 19932 21508
rect 19536 20862 19840 20890
rect 19892 20936 19944 20942
rect 19892 20878 19944 20884
rect 19432 20800 19484 20806
rect 19432 20742 19484 20748
rect 19444 19122 19472 20742
rect 19574 20700 19882 20720
rect 19574 20698 19580 20700
rect 19636 20698 19660 20700
rect 19716 20698 19740 20700
rect 19796 20698 19820 20700
rect 19876 20698 19882 20700
rect 19636 20646 19638 20698
rect 19818 20646 19820 20698
rect 19574 20644 19580 20646
rect 19636 20644 19660 20646
rect 19716 20644 19740 20646
rect 19796 20644 19820 20646
rect 19876 20644 19882 20646
rect 19574 20624 19882 20644
rect 19996 20466 20024 21558
rect 20076 20936 20128 20942
rect 20076 20878 20128 20884
rect 19984 20460 20036 20466
rect 19984 20402 20036 20408
rect 20088 19990 20116 20878
rect 20076 19984 20128 19990
rect 20076 19926 20128 19932
rect 19984 19916 20036 19922
rect 19984 19858 20036 19864
rect 19574 19612 19882 19632
rect 19574 19610 19580 19612
rect 19636 19610 19660 19612
rect 19716 19610 19740 19612
rect 19796 19610 19820 19612
rect 19876 19610 19882 19612
rect 19636 19558 19638 19610
rect 19818 19558 19820 19610
rect 19574 19556 19580 19558
rect 19636 19556 19660 19558
rect 19716 19556 19740 19558
rect 19796 19556 19820 19558
rect 19876 19556 19882 19558
rect 19574 19536 19882 19556
rect 19996 19514 20024 19858
rect 20076 19712 20128 19718
rect 20076 19654 20128 19660
rect 19984 19508 20036 19514
rect 19984 19450 20036 19456
rect 19524 19372 19576 19378
rect 19524 19314 19576 19320
rect 19708 19372 19760 19378
rect 19708 19314 19760 19320
rect 19536 19122 19564 19314
rect 19444 19094 19564 19122
rect 19444 18154 19472 19094
rect 19720 18970 19748 19314
rect 19984 19304 20036 19310
rect 19984 19246 20036 19252
rect 19708 18964 19760 18970
rect 19708 18906 19760 18912
rect 19574 18524 19882 18544
rect 19574 18522 19580 18524
rect 19636 18522 19660 18524
rect 19716 18522 19740 18524
rect 19796 18522 19820 18524
rect 19876 18522 19882 18524
rect 19636 18470 19638 18522
rect 19818 18470 19820 18522
rect 19574 18468 19580 18470
rect 19636 18468 19660 18470
rect 19716 18468 19740 18470
rect 19796 18468 19820 18470
rect 19876 18468 19882 18470
rect 19574 18448 19882 18468
rect 19892 18284 19944 18290
rect 19892 18226 19944 18232
rect 19432 18148 19484 18154
rect 19432 18090 19484 18096
rect 19432 17740 19484 17746
rect 19432 17682 19484 17688
rect 19444 17218 19472 17682
rect 19904 17524 19932 18226
rect 19996 17814 20024 19246
rect 19984 17808 20036 17814
rect 19984 17750 20036 17756
rect 20088 17762 20116 19654
rect 20180 18358 20208 21830
rect 20364 21622 20392 22510
rect 20352 21616 20404 21622
rect 20352 21558 20404 21564
rect 20352 21412 20404 21418
rect 20352 21354 20404 21360
rect 20364 21321 20392 21354
rect 20350 21312 20406 21321
rect 20350 21247 20406 21256
rect 20258 21176 20314 21185
rect 20258 21111 20314 21120
rect 20272 20806 20300 21111
rect 20364 20942 20392 21247
rect 20352 20936 20404 20942
rect 20352 20878 20404 20884
rect 20456 20874 20484 24074
rect 20548 23866 20576 24550
rect 20720 24404 20772 24410
rect 20720 24346 20772 24352
rect 20732 23866 20760 24346
rect 20536 23860 20588 23866
rect 20536 23802 20588 23808
rect 20720 23860 20772 23866
rect 20720 23802 20772 23808
rect 20536 23588 20588 23594
rect 20536 23530 20588 23536
rect 20548 21690 20576 23530
rect 20732 22778 20760 23802
rect 20824 23322 20852 24686
rect 20916 24206 20944 25706
rect 20904 24200 20956 24206
rect 20904 24142 20956 24148
rect 21192 24138 21220 26862
rect 21456 26580 21508 26586
rect 21456 26522 21508 26528
rect 21364 25152 21416 25158
rect 21364 25094 21416 25100
rect 21376 24886 21404 25094
rect 21272 24880 21324 24886
rect 21272 24822 21324 24828
rect 21364 24880 21416 24886
rect 21364 24822 21416 24828
rect 21180 24132 21232 24138
rect 21180 24074 21232 24080
rect 20996 24064 21048 24070
rect 20996 24006 21048 24012
rect 20904 23792 20956 23798
rect 20904 23734 20956 23740
rect 20812 23316 20864 23322
rect 20812 23258 20864 23264
rect 20720 22772 20772 22778
rect 20720 22714 20772 22720
rect 20824 22710 20852 23258
rect 20916 22982 20944 23734
rect 21008 23730 21036 24006
rect 21192 23866 21220 24074
rect 21180 23860 21232 23866
rect 21180 23802 21232 23808
rect 20996 23724 21048 23730
rect 20996 23666 21048 23672
rect 21008 23118 21036 23666
rect 21284 23474 21312 24822
rect 21468 24410 21496 26522
rect 21548 25764 21600 25770
rect 21548 25706 21600 25712
rect 21560 25430 21588 25706
rect 21548 25424 21600 25430
rect 21548 25366 21600 25372
rect 21456 24404 21508 24410
rect 21456 24346 21508 24352
rect 21456 24200 21508 24206
rect 21456 24142 21508 24148
rect 21364 24064 21416 24070
rect 21364 24006 21416 24012
rect 21376 23866 21404 24006
rect 21364 23860 21416 23866
rect 21364 23802 21416 23808
rect 21192 23446 21312 23474
rect 20996 23112 21048 23118
rect 20996 23054 21048 23060
rect 20904 22976 20956 22982
rect 20904 22918 20956 22924
rect 20812 22704 20864 22710
rect 20812 22646 20864 22652
rect 21008 22642 21036 23054
rect 20996 22636 21048 22642
rect 20996 22578 21048 22584
rect 20628 22568 20680 22574
rect 20628 22510 20680 22516
rect 20640 22234 20668 22510
rect 21192 22386 21220 23446
rect 21376 23338 21404 23802
rect 20732 22358 21220 22386
rect 21284 23310 21404 23338
rect 20628 22228 20680 22234
rect 20628 22170 20680 22176
rect 20732 22114 20760 22358
rect 20640 22086 20760 22114
rect 20640 22030 20668 22086
rect 20628 22024 20680 22030
rect 20628 21966 20680 21972
rect 20720 22024 20772 22030
rect 20720 21966 20772 21972
rect 20536 21684 20588 21690
rect 20536 21626 20588 21632
rect 20640 21570 20668 21966
rect 20548 21542 20668 21570
rect 20444 20868 20496 20874
rect 20444 20810 20496 20816
rect 20260 20800 20312 20806
rect 20260 20742 20312 20748
rect 20456 20466 20484 20810
rect 20444 20460 20496 20466
rect 20444 20402 20496 20408
rect 20548 20346 20576 21542
rect 20732 21350 20760 21966
rect 21088 21888 21140 21894
rect 21088 21830 21140 21836
rect 20904 21684 20956 21690
rect 20904 21626 20956 21632
rect 20628 21344 20680 21350
rect 20628 21286 20680 21292
rect 20720 21344 20772 21350
rect 20720 21286 20772 21292
rect 20640 20874 20668 21286
rect 20916 20942 20944 21626
rect 21100 21622 21128 21830
rect 21088 21616 21140 21622
rect 21088 21558 21140 21564
rect 20904 20936 20956 20942
rect 20904 20878 20956 20884
rect 20628 20868 20680 20874
rect 20628 20810 20680 20816
rect 20812 20868 20864 20874
rect 20812 20810 20864 20816
rect 20364 20318 20576 20346
rect 20168 18352 20220 18358
rect 20168 18294 20220 18300
rect 20088 17734 20208 17762
rect 20076 17672 20128 17678
rect 20076 17614 20128 17620
rect 19904 17496 20024 17524
rect 19574 17436 19882 17456
rect 19574 17434 19580 17436
rect 19636 17434 19660 17436
rect 19716 17434 19740 17436
rect 19796 17434 19820 17436
rect 19876 17434 19882 17436
rect 19636 17382 19638 17434
rect 19818 17382 19820 17434
rect 19574 17380 19580 17382
rect 19636 17380 19660 17382
rect 19716 17380 19740 17382
rect 19796 17380 19820 17382
rect 19876 17380 19882 17382
rect 19574 17360 19882 17380
rect 19996 17320 20024 17496
rect 20088 17338 20116 17614
rect 19720 17292 20024 17320
rect 20076 17332 20128 17338
rect 19444 17202 19564 17218
rect 19720 17202 19748 17292
rect 19444 17196 19576 17202
rect 19444 17190 19524 17196
rect 19524 17138 19576 17144
rect 19708 17196 19760 17202
rect 19708 17138 19760 17144
rect 19432 17128 19484 17134
rect 19432 17070 19484 17076
rect 19340 16108 19392 16114
rect 19340 16050 19392 16056
rect 19064 15904 19116 15910
rect 19064 15846 19116 15852
rect 19352 15502 19380 16050
rect 19444 15978 19472 17070
rect 19536 16726 19564 17138
rect 19524 16720 19576 16726
rect 19524 16662 19576 16668
rect 19706 16688 19762 16697
rect 19706 16623 19708 16632
rect 19760 16623 19762 16632
rect 19904 16640 19932 17292
rect 20076 17274 20128 17280
rect 20180 17202 20208 17734
rect 20364 17338 20392 20318
rect 20628 18964 20680 18970
rect 20628 18906 20680 18912
rect 20444 18216 20496 18222
rect 20444 18158 20496 18164
rect 20456 17610 20484 18158
rect 20536 17740 20588 17746
rect 20536 17682 20588 17688
rect 20444 17604 20496 17610
rect 20444 17546 20496 17552
rect 20352 17332 20404 17338
rect 20272 17292 20352 17320
rect 20168 17196 20220 17202
rect 20168 17138 20220 17144
rect 20272 17082 20300 17292
rect 20352 17274 20404 17280
rect 20352 17196 20404 17202
rect 20352 17138 20404 17144
rect 20088 17054 20300 17082
rect 20088 16998 20116 17054
rect 20076 16992 20128 16998
rect 20076 16934 20128 16940
rect 20168 16992 20220 16998
rect 20168 16934 20220 16940
rect 19904 16612 20116 16640
rect 19708 16594 19760 16600
rect 19800 16584 19852 16590
rect 19852 16532 20024 16538
rect 19800 16526 20024 16532
rect 19812 16510 20024 16526
rect 19574 16348 19882 16368
rect 19574 16346 19580 16348
rect 19636 16346 19660 16348
rect 19716 16346 19740 16348
rect 19796 16346 19820 16348
rect 19876 16346 19882 16348
rect 19636 16294 19638 16346
rect 19818 16294 19820 16346
rect 19574 16292 19580 16294
rect 19636 16292 19660 16294
rect 19716 16292 19740 16294
rect 19796 16292 19820 16294
rect 19876 16292 19882 16294
rect 19574 16272 19882 16292
rect 19616 16108 19668 16114
rect 19616 16050 19668 16056
rect 19432 15972 19484 15978
rect 19432 15914 19484 15920
rect 19628 15706 19656 16050
rect 19616 15700 19668 15706
rect 19616 15642 19668 15648
rect 19432 15632 19484 15638
rect 19432 15574 19484 15580
rect 19444 15502 19472 15574
rect 19340 15496 19392 15502
rect 19340 15438 19392 15444
rect 19432 15496 19484 15502
rect 19432 15438 19484 15444
rect 19340 15156 19392 15162
rect 19340 15098 19392 15104
rect 19352 14385 19380 15098
rect 19338 14376 19394 14385
rect 19444 14346 19472 15438
rect 19574 15260 19882 15280
rect 19574 15258 19580 15260
rect 19636 15258 19660 15260
rect 19716 15258 19740 15260
rect 19796 15258 19820 15260
rect 19876 15258 19882 15260
rect 19636 15206 19638 15258
rect 19818 15206 19820 15258
rect 19574 15204 19580 15206
rect 19636 15204 19660 15206
rect 19716 15204 19740 15206
rect 19796 15204 19820 15206
rect 19876 15204 19882 15206
rect 19574 15184 19882 15204
rect 19522 15056 19578 15065
rect 19522 14991 19578 15000
rect 19536 14890 19564 14991
rect 19524 14884 19576 14890
rect 19524 14826 19576 14832
rect 19338 14311 19394 14320
rect 19432 14340 19484 14346
rect 19432 14282 19484 14288
rect 19574 14172 19882 14192
rect 19574 14170 19580 14172
rect 19636 14170 19660 14172
rect 19716 14170 19740 14172
rect 19796 14170 19820 14172
rect 19876 14170 19882 14172
rect 19636 14118 19638 14170
rect 19818 14118 19820 14170
rect 19574 14116 19580 14118
rect 19636 14116 19660 14118
rect 19716 14116 19740 14118
rect 19796 14116 19820 14118
rect 19876 14116 19882 14118
rect 19574 14096 19882 14116
rect 19996 13410 20024 16510
rect 20088 16454 20116 16612
rect 20180 16590 20208 16934
rect 20364 16590 20392 17138
rect 20168 16584 20220 16590
rect 20168 16526 20220 16532
rect 20352 16584 20404 16590
rect 20352 16526 20404 16532
rect 20076 16448 20128 16454
rect 20076 16390 20128 16396
rect 20088 15638 20116 16390
rect 20364 16130 20392 16526
rect 20456 16522 20484 17546
rect 20548 17202 20576 17682
rect 20640 17678 20668 18906
rect 20720 18896 20772 18902
rect 20720 18838 20772 18844
rect 20732 17882 20760 18838
rect 20824 18766 20852 20810
rect 20916 19786 20944 20878
rect 20904 19780 20956 19786
rect 20904 19722 20956 19728
rect 20996 19712 21048 19718
rect 20996 19654 21048 19660
rect 21008 19334 21036 19654
rect 20916 19306 21036 19334
rect 20812 18760 20864 18766
rect 20812 18702 20864 18708
rect 20720 17876 20772 17882
rect 20720 17818 20772 17824
rect 20628 17672 20680 17678
rect 20628 17614 20680 17620
rect 20536 17196 20588 17202
rect 20536 17138 20588 17144
rect 20444 16516 20496 16522
rect 20444 16458 20496 16464
rect 20456 16182 20484 16458
rect 20168 16108 20220 16114
rect 20168 16050 20220 16056
rect 20272 16102 20392 16130
rect 20444 16176 20496 16182
rect 20444 16118 20496 16124
rect 20076 15632 20128 15638
rect 20076 15574 20128 15580
rect 20076 15020 20128 15026
rect 20076 14962 20128 14968
rect 20088 14618 20116 14962
rect 20180 14822 20208 16050
rect 20272 15502 20300 16102
rect 20352 15972 20404 15978
rect 20352 15914 20404 15920
rect 20364 15570 20392 15914
rect 20444 15632 20496 15638
rect 20444 15574 20496 15580
rect 20352 15564 20404 15570
rect 20352 15506 20404 15512
rect 20260 15496 20312 15502
rect 20260 15438 20312 15444
rect 20456 15416 20484 15574
rect 20364 15388 20484 15416
rect 20260 15360 20312 15366
rect 20260 15302 20312 15308
rect 20168 14816 20220 14822
rect 20168 14758 20220 14764
rect 20076 14612 20128 14618
rect 20076 14554 20128 14560
rect 20180 13938 20208 14758
rect 20272 14414 20300 15302
rect 20364 14958 20392 15388
rect 20548 15314 20576 17138
rect 20640 16114 20668 17614
rect 20732 17610 20760 17818
rect 20720 17604 20772 17610
rect 20720 17546 20772 17552
rect 20812 17536 20864 17542
rect 20810 17504 20812 17513
rect 20864 17504 20866 17513
rect 20810 17439 20866 17448
rect 20720 16516 20772 16522
rect 20720 16458 20772 16464
rect 20628 16108 20680 16114
rect 20628 16050 20680 16056
rect 20626 16008 20682 16017
rect 20626 15943 20682 15952
rect 20640 15910 20668 15943
rect 20628 15904 20680 15910
rect 20628 15846 20680 15852
rect 20732 15314 20760 16458
rect 20916 15638 20944 19306
rect 21284 18902 21312 23310
rect 21468 23050 21496 24142
rect 21456 23044 21508 23050
rect 21456 22986 21508 22992
rect 21560 22030 21588 25366
rect 21652 23594 21680 26862
rect 22204 26382 22232 26930
rect 22192 26376 22244 26382
rect 22244 26324 22324 26330
rect 22192 26318 22324 26324
rect 22204 26302 22324 26318
rect 21916 26240 21968 26246
rect 21916 26182 21968 26188
rect 21732 25968 21784 25974
rect 21732 25910 21784 25916
rect 21744 25498 21772 25910
rect 21732 25492 21784 25498
rect 21732 25434 21784 25440
rect 21732 25220 21784 25226
rect 21732 25162 21784 25168
rect 21640 23588 21692 23594
rect 21640 23530 21692 23536
rect 21640 23248 21692 23254
rect 21640 23190 21692 23196
rect 21456 22024 21508 22030
rect 21456 21966 21508 21972
rect 21548 22024 21600 22030
rect 21548 21966 21600 21972
rect 21364 21956 21416 21962
rect 21364 21898 21416 21904
rect 21376 21010 21404 21898
rect 21468 21418 21496 21966
rect 21560 21690 21588 21966
rect 21652 21894 21680 23190
rect 21744 21962 21772 25162
rect 21824 22636 21876 22642
rect 21824 22578 21876 22584
rect 21836 22234 21864 22578
rect 21824 22228 21876 22234
rect 21824 22170 21876 22176
rect 21824 22092 21876 22098
rect 21824 22034 21876 22040
rect 21732 21956 21784 21962
rect 21732 21898 21784 21904
rect 21640 21888 21692 21894
rect 21640 21830 21692 21836
rect 21548 21684 21600 21690
rect 21548 21626 21600 21632
rect 21456 21412 21508 21418
rect 21456 21354 21508 21360
rect 21364 21004 21416 21010
rect 21364 20946 21416 20952
rect 21272 18896 21324 18902
rect 21272 18838 21324 18844
rect 21376 18698 21404 20946
rect 21468 19446 21496 21354
rect 21652 20942 21680 21830
rect 21836 21418 21864 22034
rect 21824 21412 21876 21418
rect 21824 21354 21876 21360
rect 21822 21312 21878 21321
rect 21822 21247 21878 21256
rect 21836 20942 21864 21247
rect 21640 20936 21692 20942
rect 21640 20878 21692 20884
rect 21824 20936 21876 20942
rect 21824 20878 21876 20884
rect 21456 19440 21508 19446
rect 21456 19382 21508 19388
rect 21456 19304 21508 19310
rect 21456 19246 21508 19252
rect 21468 18834 21496 19246
rect 21456 18828 21508 18834
rect 21456 18770 21508 18776
rect 21364 18692 21416 18698
rect 21364 18634 21416 18640
rect 21652 17066 21680 20878
rect 21732 20800 21784 20806
rect 21732 20742 21784 20748
rect 21744 20602 21772 20742
rect 21928 20602 21956 26182
rect 22296 25906 22324 26302
rect 22284 25900 22336 25906
rect 22284 25842 22336 25848
rect 22192 25492 22244 25498
rect 22192 25434 22244 25440
rect 22204 22642 22232 25434
rect 22192 22636 22244 22642
rect 22192 22578 22244 22584
rect 22008 22432 22060 22438
rect 22008 22374 22060 22380
rect 21732 20596 21784 20602
rect 21732 20538 21784 20544
rect 21916 20596 21968 20602
rect 21916 20538 21968 20544
rect 21928 19242 21956 20538
rect 21916 19236 21968 19242
rect 21916 19178 21968 19184
rect 21732 18760 21784 18766
rect 21732 18702 21784 18708
rect 21640 17060 21692 17066
rect 21640 17002 21692 17008
rect 21272 16584 21324 16590
rect 21272 16526 21324 16532
rect 21284 16250 21312 16526
rect 21272 16244 21324 16250
rect 21272 16186 21324 16192
rect 20996 16176 21048 16182
rect 20996 16118 21048 16124
rect 20904 15632 20956 15638
rect 20904 15574 20956 15580
rect 20456 15286 20576 15314
rect 20640 15286 20760 15314
rect 20352 14952 20404 14958
rect 20352 14894 20404 14900
rect 20260 14408 20312 14414
rect 20260 14350 20312 14356
rect 20168 13932 20220 13938
rect 20168 13874 20220 13880
rect 20272 13870 20300 14350
rect 20352 13932 20404 13938
rect 20352 13874 20404 13880
rect 20260 13864 20312 13870
rect 20260 13806 20312 13812
rect 20168 13796 20220 13802
rect 20168 13738 20220 13744
rect 20180 13462 20208 13738
rect 20168 13456 20220 13462
rect 19996 13382 20116 13410
rect 20168 13398 20220 13404
rect 19340 13320 19392 13326
rect 19340 13262 19392 13268
rect 19982 13288 20038 13297
rect 19352 12986 19380 13262
rect 19982 13223 19984 13232
rect 20036 13223 20038 13232
rect 19984 13194 20036 13200
rect 19574 13084 19882 13104
rect 19574 13082 19580 13084
rect 19636 13082 19660 13084
rect 19716 13082 19740 13084
rect 19796 13082 19820 13084
rect 19876 13082 19882 13084
rect 19636 13030 19638 13082
rect 19818 13030 19820 13082
rect 19574 13028 19580 13030
rect 19636 13028 19660 13030
rect 19716 13028 19740 13030
rect 19796 13028 19820 13030
rect 19876 13028 19882 13030
rect 19574 13008 19882 13028
rect 20088 12986 20116 13382
rect 19340 12980 19392 12986
rect 19340 12922 19392 12928
rect 19432 12980 19484 12986
rect 19432 12922 19484 12928
rect 20076 12980 20128 12986
rect 20076 12922 20128 12928
rect 19340 12368 19392 12374
rect 19340 12310 19392 12316
rect 19248 12096 19300 12102
rect 19248 12038 19300 12044
rect 19156 10192 19208 10198
rect 19156 10134 19208 10140
rect 19168 9586 19196 10134
rect 19260 10062 19288 12038
rect 19352 11898 19380 12310
rect 19444 12238 19472 12922
rect 20088 12850 20116 12922
rect 20076 12844 20128 12850
rect 20076 12786 20128 12792
rect 20180 12322 20208 13398
rect 20364 13258 20392 13874
rect 20352 13252 20404 13258
rect 20352 13194 20404 13200
rect 20364 12782 20392 13194
rect 20352 12776 20404 12782
rect 20352 12718 20404 12724
rect 20088 12294 20208 12322
rect 19432 12232 19484 12238
rect 19432 12174 19484 12180
rect 19574 11996 19882 12016
rect 19574 11994 19580 11996
rect 19636 11994 19660 11996
rect 19716 11994 19740 11996
rect 19796 11994 19820 11996
rect 19876 11994 19882 11996
rect 19636 11942 19638 11994
rect 19818 11942 19820 11994
rect 19574 11940 19580 11942
rect 19636 11940 19660 11942
rect 19716 11940 19740 11942
rect 19796 11940 19820 11942
rect 19876 11940 19882 11942
rect 19574 11920 19882 11940
rect 19340 11892 19392 11898
rect 19340 11834 19392 11840
rect 19352 11762 19380 11834
rect 19340 11756 19392 11762
rect 19340 11698 19392 11704
rect 19340 11212 19392 11218
rect 19340 11154 19392 11160
rect 19248 10056 19300 10062
rect 19248 9998 19300 10004
rect 19156 9580 19208 9586
rect 19156 9522 19208 9528
rect 19260 8974 19288 9998
rect 19352 9625 19380 11154
rect 19984 11144 20036 11150
rect 19984 11086 20036 11092
rect 19574 10908 19882 10928
rect 19574 10906 19580 10908
rect 19636 10906 19660 10908
rect 19716 10906 19740 10908
rect 19796 10906 19820 10908
rect 19876 10906 19882 10908
rect 19636 10854 19638 10906
rect 19818 10854 19820 10906
rect 19574 10852 19580 10854
rect 19636 10852 19660 10854
rect 19716 10852 19740 10854
rect 19796 10852 19820 10854
rect 19876 10852 19882 10854
rect 19574 10832 19882 10852
rect 19708 10668 19760 10674
rect 19996 10656 20024 11086
rect 20088 10742 20116 12294
rect 20364 12238 20392 12718
rect 20168 12232 20220 12238
rect 20168 12174 20220 12180
rect 20352 12232 20404 12238
rect 20352 12174 20404 12180
rect 20180 11898 20208 12174
rect 20168 11892 20220 11898
rect 20168 11834 20220 11840
rect 20456 11762 20484 15286
rect 20536 15156 20588 15162
rect 20640 15144 20668 15286
rect 20588 15116 20668 15144
rect 20718 15192 20774 15201
rect 20718 15127 20720 15136
rect 20536 15098 20588 15104
rect 20772 15127 20774 15136
rect 20720 15098 20772 15104
rect 21008 15094 21036 16118
rect 21744 16046 21772 18702
rect 21824 18692 21876 18698
rect 21824 18634 21876 18640
rect 21836 18290 21864 18634
rect 21824 18284 21876 18290
rect 21824 18226 21876 18232
rect 21928 17678 21956 19178
rect 22020 18714 22048 22374
rect 22100 21888 22152 21894
rect 22098 21856 22100 21865
rect 22152 21856 22154 21865
rect 22098 21791 22154 21800
rect 22204 21321 22232 22578
rect 22388 22094 22416 29446
rect 23124 29306 23152 29650
rect 23848 29640 23900 29646
rect 23848 29582 23900 29588
rect 23112 29300 23164 29306
rect 23112 29242 23164 29248
rect 22744 29164 22796 29170
rect 22744 29106 22796 29112
rect 22468 28960 22520 28966
rect 22468 28902 22520 28908
rect 22480 28558 22508 28902
rect 22756 28694 22784 29106
rect 23294 29064 23350 29073
rect 23294 28999 23350 29008
rect 22744 28688 22796 28694
rect 22744 28630 22796 28636
rect 22468 28552 22520 28558
rect 22468 28494 22520 28500
rect 22296 22066 22416 22094
rect 22190 21312 22246 21321
rect 22112 21270 22190 21298
rect 22112 19446 22140 21270
rect 22190 21247 22246 21256
rect 22192 19712 22244 19718
rect 22192 19654 22244 19660
rect 22100 19440 22152 19446
rect 22100 19382 22152 19388
rect 22204 19378 22232 19654
rect 22192 19372 22244 19378
rect 22192 19314 22244 19320
rect 22100 18828 22152 18834
rect 22100 18770 22152 18776
rect 22112 18714 22140 18770
rect 22020 18686 22140 18714
rect 22020 18426 22048 18686
rect 22008 18420 22060 18426
rect 22008 18362 22060 18368
rect 22100 18420 22152 18426
rect 22100 18362 22152 18368
rect 22112 17882 22140 18362
rect 22100 17876 22152 17882
rect 22100 17818 22152 17824
rect 21916 17672 21968 17678
rect 21916 17614 21968 17620
rect 22296 17218 22324 22066
rect 22376 20868 22428 20874
rect 22376 20810 22428 20816
rect 22388 20602 22416 20810
rect 22376 20596 22428 20602
rect 22376 20538 22428 20544
rect 22376 19508 22428 19514
rect 22376 19450 22428 19456
rect 22388 18970 22416 19450
rect 22480 19334 22508 28494
rect 22560 28484 22612 28490
rect 22560 28426 22612 28432
rect 22572 22094 22600 28426
rect 22836 28416 22888 28422
rect 22836 28358 22888 28364
rect 22848 27606 22876 28358
rect 22836 27600 22888 27606
rect 22836 27542 22888 27548
rect 22744 27328 22796 27334
rect 22744 27270 22796 27276
rect 22928 27328 22980 27334
rect 22928 27270 22980 27276
rect 22756 26518 22784 27270
rect 22836 26988 22888 26994
rect 22836 26930 22888 26936
rect 22744 26512 22796 26518
rect 22744 26454 22796 26460
rect 22848 26450 22876 26930
rect 22836 26444 22888 26450
rect 22836 26386 22888 26392
rect 22940 25838 22968 27270
rect 23308 26382 23336 28999
rect 23860 28694 23888 29582
rect 24124 29504 24176 29510
rect 24124 29446 24176 29452
rect 24136 29102 24164 29446
rect 24124 29096 24176 29102
rect 24124 29038 24176 29044
rect 23848 28688 23900 28694
rect 23848 28630 23900 28636
rect 23664 28552 23716 28558
rect 23664 28494 23716 28500
rect 23676 28014 23704 28494
rect 24136 28082 24164 29038
rect 24320 29034 24348 30126
rect 24412 29646 24440 30330
rect 24780 30054 24808 30534
rect 24860 30252 24912 30258
rect 24860 30194 24912 30200
rect 24768 30048 24820 30054
rect 24768 29990 24820 29996
rect 24780 29646 24808 29990
rect 24872 29782 24900 30194
rect 24860 29776 24912 29782
rect 24860 29718 24912 29724
rect 24400 29640 24452 29646
rect 24400 29582 24452 29588
rect 24768 29640 24820 29646
rect 24768 29582 24820 29588
rect 24860 29300 24912 29306
rect 24860 29242 24912 29248
rect 24584 29096 24636 29102
rect 24584 29038 24636 29044
rect 24308 29028 24360 29034
rect 24308 28970 24360 28976
rect 24320 28558 24348 28970
rect 24596 28558 24624 29038
rect 24872 28762 24900 29242
rect 24860 28756 24912 28762
rect 24860 28698 24912 28704
rect 24768 28688 24820 28694
rect 24768 28630 24820 28636
rect 24308 28552 24360 28558
rect 24308 28494 24360 28500
rect 24584 28552 24636 28558
rect 24584 28494 24636 28500
rect 24124 28076 24176 28082
rect 24124 28018 24176 28024
rect 23664 28008 23716 28014
rect 23664 27950 23716 27956
rect 24216 28008 24268 28014
rect 24216 27950 24268 27956
rect 23676 27470 23704 27950
rect 24228 27878 24256 27950
rect 24216 27872 24268 27878
rect 24216 27814 24268 27820
rect 23664 27464 23716 27470
rect 23664 27406 23716 27412
rect 23388 27328 23440 27334
rect 23388 27270 23440 27276
rect 23400 26450 23428 27270
rect 23676 26994 23704 27406
rect 23664 26988 23716 26994
rect 23664 26930 23716 26936
rect 23572 26784 23624 26790
rect 23572 26726 23624 26732
rect 23388 26444 23440 26450
rect 23388 26386 23440 26392
rect 23296 26376 23348 26382
rect 23296 26318 23348 26324
rect 22928 25832 22980 25838
rect 22928 25774 22980 25780
rect 22744 24064 22796 24070
rect 22744 24006 22796 24012
rect 22572 22066 22692 22094
rect 22480 19306 22600 19334
rect 22376 18964 22428 18970
rect 22376 18906 22428 18912
rect 22204 17190 22324 17218
rect 21732 16040 21784 16046
rect 21732 15982 21784 15988
rect 21086 15736 21142 15745
rect 21086 15671 21142 15680
rect 20996 15088 21048 15094
rect 20996 15030 21048 15036
rect 20536 15020 20588 15026
rect 20536 14962 20588 14968
rect 20548 14822 20576 14962
rect 20720 14884 20772 14890
rect 20720 14826 20772 14832
rect 20536 14816 20588 14822
rect 20732 14793 20760 14826
rect 20536 14758 20588 14764
rect 20718 14784 20774 14793
rect 20718 14719 20774 14728
rect 20536 14612 20588 14618
rect 20536 14554 20588 14560
rect 20548 14482 20576 14554
rect 20536 14476 20588 14482
rect 20536 14418 20588 14424
rect 20812 14476 20864 14482
rect 20812 14418 20864 14424
rect 20548 13326 20576 14418
rect 20824 14006 20852 14418
rect 21008 14414 21036 15030
rect 20996 14408 21048 14414
rect 20996 14350 21048 14356
rect 20812 14000 20864 14006
rect 20812 13942 20864 13948
rect 20904 13932 20956 13938
rect 20904 13874 20956 13880
rect 20916 13841 20944 13874
rect 20902 13832 20958 13841
rect 20902 13767 20958 13776
rect 20996 13796 21048 13802
rect 20996 13738 21048 13744
rect 20536 13320 20588 13326
rect 20536 13262 20588 13268
rect 20626 12200 20682 12209
rect 21008 12170 21036 13738
rect 21100 12374 21128 15671
rect 21744 15502 21772 15982
rect 21732 15496 21784 15502
rect 21732 15438 21784 15444
rect 21916 15360 21968 15366
rect 21916 15302 21968 15308
rect 21824 14544 21876 14550
rect 21928 14532 21956 15302
rect 22100 15088 22152 15094
rect 22100 15030 22152 15036
rect 21876 14504 21956 14532
rect 21824 14486 21876 14492
rect 21180 14408 21232 14414
rect 21180 14350 21232 14356
rect 21640 14408 21692 14414
rect 21640 14350 21692 14356
rect 21192 12442 21220 14350
rect 21652 14006 21680 14350
rect 21824 14272 21876 14278
rect 21824 14214 21876 14220
rect 21640 14000 21692 14006
rect 21640 13942 21692 13948
rect 21836 13841 21864 14214
rect 21928 13938 21956 14504
rect 22008 14408 22060 14414
rect 22008 14350 22060 14356
rect 21916 13932 21968 13938
rect 21916 13874 21968 13880
rect 21822 13832 21878 13841
rect 21364 13796 21416 13802
rect 21822 13767 21878 13776
rect 21364 13738 21416 13744
rect 21376 13394 21404 13738
rect 21364 13388 21416 13394
rect 21364 13330 21416 13336
rect 21180 12436 21232 12442
rect 21180 12378 21232 12384
rect 21088 12368 21140 12374
rect 21088 12310 21140 12316
rect 21192 12238 21220 12378
rect 21454 12336 21510 12345
rect 21454 12271 21510 12280
rect 21180 12232 21232 12238
rect 21180 12174 21232 12180
rect 21468 12170 21496 12271
rect 20626 12135 20628 12144
rect 20680 12135 20682 12144
rect 20996 12164 21048 12170
rect 20628 12106 20680 12112
rect 20996 12106 21048 12112
rect 21456 12164 21508 12170
rect 21836 12152 21864 13767
rect 21916 12164 21968 12170
rect 21836 12124 21916 12152
rect 21456 12106 21508 12112
rect 21916 12106 21968 12112
rect 20444 11756 20496 11762
rect 20444 11698 20496 11704
rect 20076 10736 20128 10742
rect 20076 10678 20128 10684
rect 19760 10628 20024 10656
rect 19708 10610 19760 10616
rect 20352 10600 20404 10606
rect 20352 10542 20404 10548
rect 20364 10198 20392 10542
rect 20352 10192 20404 10198
rect 20352 10134 20404 10140
rect 20260 10056 20312 10062
rect 20260 9998 20312 10004
rect 19574 9820 19882 9840
rect 19574 9818 19580 9820
rect 19636 9818 19660 9820
rect 19716 9818 19740 9820
rect 19796 9818 19820 9820
rect 19876 9818 19882 9820
rect 19636 9766 19638 9818
rect 19818 9766 19820 9818
rect 19574 9764 19580 9766
rect 19636 9764 19660 9766
rect 19716 9764 19740 9766
rect 19796 9764 19820 9766
rect 19876 9764 19882 9766
rect 19574 9744 19882 9764
rect 19338 9616 19394 9625
rect 19338 9551 19394 9560
rect 20168 9376 20220 9382
rect 20168 9318 20220 9324
rect 19248 8968 19300 8974
rect 19524 8968 19576 8974
rect 19248 8910 19300 8916
rect 19444 8928 19524 8956
rect 19444 8498 19472 8928
rect 19524 8910 19576 8916
rect 19574 8732 19882 8752
rect 19574 8730 19580 8732
rect 19636 8730 19660 8732
rect 19716 8730 19740 8732
rect 19796 8730 19820 8732
rect 19876 8730 19882 8732
rect 19636 8678 19638 8730
rect 19818 8678 19820 8730
rect 19574 8676 19580 8678
rect 19636 8676 19660 8678
rect 19716 8676 19740 8678
rect 19796 8676 19820 8678
rect 19876 8676 19882 8678
rect 19574 8656 19882 8676
rect 19432 8492 19484 8498
rect 19432 8434 19484 8440
rect 20180 7954 20208 9318
rect 20272 8974 20300 9998
rect 20364 9586 20392 10134
rect 20456 10062 20484 11698
rect 21008 11218 21036 12106
rect 21272 12096 21324 12102
rect 21272 12038 21324 12044
rect 21284 11898 21312 12038
rect 21272 11892 21324 11898
rect 21272 11834 21324 11840
rect 21468 11830 21496 12106
rect 21456 11824 21508 11830
rect 21456 11766 21508 11772
rect 21088 11552 21140 11558
rect 21088 11494 21140 11500
rect 20996 11212 21048 11218
rect 20996 11154 21048 11160
rect 21100 11150 21128 11494
rect 21088 11144 21140 11150
rect 21088 11086 21140 11092
rect 21928 11082 21956 12106
rect 20536 11076 20588 11082
rect 20536 11018 20588 11024
rect 21916 11076 21968 11082
rect 21916 11018 21968 11024
rect 20444 10056 20496 10062
rect 20444 9998 20496 10004
rect 20548 9654 20576 11018
rect 21928 10985 21956 11018
rect 21914 10976 21970 10985
rect 21914 10911 21970 10920
rect 21824 10260 21876 10266
rect 21824 10202 21876 10208
rect 21836 10062 21864 10202
rect 21824 10056 21876 10062
rect 21824 9998 21876 10004
rect 20536 9648 20588 9654
rect 20536 9590 20588 9596
rect 20352 9580 20404 9586
rect 20352 9522 20404 9528
rect 20548 9058 20576 9590
rect 20628 9580 20680 9586
rect 20628 9522 20680 9528
rect 20720 9580 20772 9586
rect 20720 9522 20772 9528
rect 20640 9178 20668 9522
rect 20732 9353 20760 9522
rect 20718 9344 20774 9353
rect 20718 9279 20774 9288
rect 20628 9172 20680 9178
rect 20628 9114 20680 9120
rect 20548 9042 20944 9058
rect 20548 9036 20956 9042
rect 20548 9030 20904 9036
rect 20904 8978 20956 8984
rect 20260 8968 20312 8974
rect 20260 8910 20312 8916
rect 20260 8832 20312 8838
rect 20260 8774 20312 8780
rect 20168 7948 20220 7954
rect 20168 7890 20220 7896
rect 20272 7886 20300 8774
rect 22020 8634 22048 14350
rect 22112 14074 22140 15030
rect 22100 14068 22152 14074
rect 22100 14010 22152 14016
rect 22112 13326 22140 14010
rect 22100 13320 22152 13326
rect 22100 13262 22152 13268
rect 22100 13184 22152 13190
rect 22100 13126 22152 13132
rect 22112 12238 22140 13126
rect 22100 12232 22152 12238
rect 22100 12174 22152 12180
rect 22112 11694 22140 12174
rect 22100 11688 22152 11694
rect 22100 11630 22152 11636
rect 21180 8628 21232 8634
rect 21180 8570 21232 8576
rect 22008 8628 22060 8634
rect 22008 8570 22060 8576
rect 21192 7886 21220 8570
rect 21364 8288 21416 8294
rect 21364 8230 21416 8236
rect 21376 7954 21404 8230
rect 21364 7948 21416 7954
rect 21364 7890 21416 7896
rect 20260 7880 20312 7886
rect 20260 7822 20312 7828
rect 21180 7880 21232 7886
rect 21180 7822 21232 7828
rect 20628 7812 20680 7818
rect 20628 7754 20680 7760
rect 19984 7744 20036 7750
rect 19984 7686 20036 7692
rect 19574 7644 19882 7664
rect 19574 7642 19580 7644
rect 19636 7642 19660 7644
rect 19716 7642 19740 7644
rect 19796 7642 19820 7644
rect 19876 7642 19882 7644
rect 19636 7590 19638 7642
rect 19818 7590 19820 7642
rect 19574 7588 19580 7590
rect 19636 7588 19660 7590
rect 19716 7588 19740 7590
rect 19796 7588 19820 7590
rect 19876 7588 19882 7590
rect 19574 7568 19882 7588
rect 19996 6934 20024 7686
rect 20640 7546 20668 7754
rect 20628 7540 20680 7546
rect 20628 7482 20680 7488
rect 20260 7268 20312 7274
rect 20260 7210 20312 7216
rect 19984 6928 20036 6934
rect 19984 6870 20036 6876
rect 19574 6556 19882 6576
rect 19574 6554 19580 6556
rect 19636 6554 19660 6556
rect 19716 6554 19740 6556
rect 19796 6554 19820 6556
rect 19876 6554 19882 6556
rect 19636 6502 19638 6554
rect 19818 6502 19820 6554
rect 19574 6500 19580 6502
rect 19636 6500 19660 6502
rect 19716 6500 19740 6502
rect 19796 6500 19820 6502
rect 19876 6500 19882 6502
rect 19574 6480 19882 6500
rect 19996 6254 20024 6870
rect 20272 6866 20300 7210
rect 20260 6860 20312 6866
rect 20260 6802 20312 6808
rect 20272 6322 20300 6802
rect 20444 6724 20496 6730
rect 20444 6666 20496 6672
rect 21088 6724 21140 6730
rect 21088 6666 21140 6672
rect 20456 6322 20484 6666
rect 20996 6452 21048 6458
rect 20996 6394 21048 6400
rect 20260 6316 20312 6322
rect 20260 6258 20312 6264
rect 20444 6316 20496 6322
rect 20444 6258 20496 6264
rect 19984 6248 20036 6254
rect 19984 6190 20036 6196
rect 20352 6248 20404 6254
rect 20352 6190 20404 6196
rect 20168 5840 20220 5846
rect 20168 5782 20220 5788
rect 19984 5772 20036 5778
rect 19984 5714 20036 5720
rect 19432 5636 19484 5642
rect 19432 5578 19484 5584
rect 19340 5568 19392 5574
rect 19340 5510 19392 5516
rect 19352 5302 19380 5510
rect 19340 5296 19392 5302
rect 19340 5238 19392 5244
rect 19444 5030 19472 5578
rect 19574 5468 19882 5488
rect 19574 5466 19580 5468
rect 19636 5466 19660 5468
rect 19716 5466 19740 5468
rect 19796 5466 19820 5468
rect 19876 5466 19882 5468
rect 19636 5414 19638 5466
rect 19818 5414 19820 5466
rect 19574 5412 19580 5414
rect 19636 5412 19660 5414
rect 19716 5412 19740 5414
rect 19796 5412 19820 5414
rect 19876 5412 19882 5414
rect 19574 5392 19882 5412
rect 19996 5302 20024 5714
rect 19984 5296 20036 5302
rect 19984 5238 20036 5244
rect 20180 5166 20208 5782
rect 20364 5710 20392 6190
rect 21008 5914 21036 6394
rect 21100 6390 21128 6666
rect 21088 6384 21140 6390
rect 21088 6326 21140 6332
rect 20996 5908 21048 5914
rect 20996 5850 21048 5856
rect 21008 5710 21036 5850
rect 21100 5710 21128 6326
rect 20352 5704 20404 5710
rect 20352 5646 20404 5652
rect 20996 5704 21048 5710
rect 20996 5646 21048 5652
rect 21088 5704 21140 5710
rect 21088 5646 21140 5652
rect 20168 5160 20220 5166
rect 20168 5102 20220 5108
rect 19432 5024 19484 5030
rect 19432 4966 19484 4972
rect 19892 5024 19944 5030
rect 19892 4966 19944 4972
rect 20076 5024 20128 5030
rect 20076 4966 20128 4972
rect 19904 4826 19932 4966
rect 19892 4820 19944 4826
rect 19892 4762 19944 4768
rect 20088 4622 20116 4966
rect 20076 4616 20128 4622
rect 20076 4558 20128 4564
rect 20180 4554 20208 5102
rect 20168 4548 20220 4554
rect 20168 4490 20220 4496
rect 19574 4380 19882 4400
rect 19574 4378 19580 4380
rect 19636 4378 19660 4380
rect 19716 4378 19740 4380
rect 19796 4378 19820 4380
rect 19876 4378 19882 4380
rect 19636 4326 19638 4378
rect 19818 4326 19820 4378
rect 19574 4324 19580 4326
rect 19636 4324 19660 4326
rect 19716 4324 19740 4326
rect 19796 4324 19820 4326
rect 19876 4324 19882 4326
rect 19574 4304 19882 4324
rect 20536 4276 20588 4282
rect 20536 4218 20588 4224
rect 20260 4140 20312 4146
rect 20260 4082 20312 4088
rect 20272 3534 20300 4082
rect 19248 3528 19300 3534
rect 19432 3528 19484 3534
rect 19248 3470 19300 3476
rect 19352 3488 19432 3516
rect 19260 3194 19288 3470
rect 19352 3398 19380 3488
rect 19432 3470 19484 3476
rect 20260 3528 20312 3534
rect 20260 3470 20312 3476
rect 19340 3392 19392 3398
rect 19340 3334 19392 3340
rect 19352 3194 19380 3334
rect 19574 3292 19882 3312
rect 19574 3290 19580 3292
rect 19636 3290 19660 3292
rect 19716 3290 19740 3292
rect 19796 3290 19820 3292
rect 19876 3290 19882 3292
rect 19636 3238 19638 3290
rect 19818 3238 19820 3290
rect 19574 3236 19580 3238
rect 19636 3236 19660 3238
rect 19716 3236 19740 3238
rect 19796 3236 19820 3238
rect 19876 3236 19882 3238
rect 19574 3216 19882 3236
rect 19248 3188 19300 3194
rect 19248 3130 19300 3136
rect 19340 3188 19392 3194
rect 19340 3130 19392 3136
rect 20548 2922 20576 4218
rect 20628 4140 20680 4146
rect 20628 4082 20680 4088
rect 20640 3398 20668 4082
rect 20904 3664 20956 3670
rect 20904 3606 20956 3612
rect 20628 3392 20680 3398
rect 20628 3334 20680 3340
rect 20640 3058 20668 3334
rect 20628 3052 20680 3058
rect 20628 2994 20680 3000
rect 20916 2990 20944 3606
rect 21088 3528 21140 3534
rect 21088 3470 21140 3476
rect 20904 2984 20956 2990
rect 20904 2926 20956 2932
rect 20536 2916 20588 2922
rect 20536 2858 20588 2864
rect 20548 2774 20576 2858
rect 20916 2774 20944 2926
rect 18984 2746 19196 2774
rect 20548 2746 20668 2774
rect 19168 2446 19196 2746
rect 20640 2514 20668 2746
rect 20824 2746 20944 2774
rect 20628 2508 20680 2514
rect 20628 2450 20680 2456
rect 20824 2446 20852 2746
rect 21100 2514 21128 3470
rect 21192 2774 21220 7822
rect 21376 6662 21404 7890
rect 21364 6656 21416 6662
rect 21364 6598 21416 6604
rect 22204 4078 22232 17190
rect 22376 16176 22428 16182
rect 22376 16118 22428 16124
rect 22388 15978 22416 16118
rect 22376 15972 22428 15978
rect 22376 15914 22428 15920
rect 22284 15360 22336 15366
rect 22284 15302 22336 15308
rect 22296 14618 22324 15302
rect 22284 14612 22336 14618
rect 22284 14554 22336 14560
rect 22388 14346 22416 15914
rect 22376 14340 22428 14346
rect 22376 14282 22428 14288
rect 22388 14074 22416 14282
rect 22376 14068 22428 14074
rect 22376 14010 22428 14016
rect 22284 13728 22336 13734
rect 22284 13670 22336 13676
rect 22468 13728 22520 13734
rect 22468 13670 22520 13676
rect 22296 12322 22324 13670
rect 22480 13161 22508 13670
rect 22466 13152 22522 13161
rect 22466 13087 22522 13096
rect 22296 12294 22508 12322
rect 22480 12238 22508 12294
rect 22376 12232 22428 12238
rect 22376 12174 22428 12180
rect 22468 12232 22520 12238
rect 22468 12174 22520 12180
rect 22284 11756 22336 11762
rect 22284 11698 22336 11704
rect 22296 11354 22324 11698
rect 22388 11354 22416 12174
rect 22284 11348 22336 11354
rect 22284 11290 22336 11296
rect 22376 11348 22428 11354
rect 22376 11290 22428 11296
rect 22480 10266 22508 12174
rect 22468 10260 22520 10266
rect 22468 10202 22520 10208
rect 22376 9920 22428 9926
rect 22376 9862 22428 9868
rect 22284 9444 22336 9450
rect 22284 9386 22336 9392
rect 22296 8838 22324 9386
rect 22284 8832 22336 8838
rect 22284 8774 22336 8780
rect 22388 7954 22416 9862
rect 22468 9376 22520 9382
rect 22468 9318 22520 9324
rect 22480 8974 22508 9318
rect 22468 8968 22520 8974
rect 22468 8910 22520 8916
rect 22376 7948 22428 7954
rect 22376 7890 22428 7896
rect 21640 4072 21692 4078
rect 21640 4014 21692 4020
rect 22192 4072 22244 4078
rect 22192 4014 22244 4020
rect 21652 3534 21680 4014
rect 21640 3528 21692 3534
rect 21640 3470 21692 3476
rect 21652 3126 21680 3470
rect 21640 3120 21692 3126
rect 21640 3062 21692 3068
rect 21732 3052 21784 3058
rect 21732 2994 21784 3000
rect 21744 2854 21772 2994
rect 21732 2848 21784 2854
rect 21732 2790 21784 2796
rect 21916 2848 21968 2854
rect 21916 2790 21968 2796
rect 21192 2746 21312 2774
rect 21284 2650 21312 2746
rect 21272 2644 21324 2650
rect 21272 2586 21324 2592
rect 21088 2508 21140 2514
rect 21088 2450 21140 2456
rect 21928 2446 21956 2790
rect 22572 2650 22600 19306
rect 22664 13258 22692 22066
rect 22756 21350 22784 24006
rect 22836 21548 22888 21554
rect 22836 21490 22888 21496
rect 22744 21344 22796 21350
rect 22744 21286 22796 21292
rect 22848 21078 22876 21490
rect 22836 21072 22888 21078
rect 22836 21014 22888 21020
rect 22744 19440 22796 19446
rect 22744 19382 22796 19388
rect 22756 17270 22784 19382
rect 22744 17264 22796 17270
rect 22744 17206 22796 17212
rect 22836 16108 22888 16114
rect 22836 16050 22888 16056
rect 22848 15706 22876 16050
rect 22836 15700 22888 15706
rect 22836 15642 22888 15648
rect 22940 13938 22968 25774
rect 23400 25294 23428 26386
rect 23584 26382 23612 26726
rect 23572 26376 23624 26382
rect 23572 26318 23624 26324
rect 23940 26376 23992 26382
rect 23940 26318 23992 26324
rect 23584 25294 23612 26318
rect 23952 25702 23980 26318
rect 24124 26308 24176 26314
rect 24124 26250 24176 26256
rect 24032 26240 24084 26246
rect 24032 26182 24084 26188
rect 24044 25906 24072 26182
rect 24032 25900 24084 25906
rect 24032 25842 24084 25848
rect 23940 25696 23992 25702
rect 23940 25638 23992 25644
rect 23388 25288 23440 25294
rect 23388 25230 23440 25236
rect 23572 25288 23624 25294
rect 23572 25230 23624 25236
rect 23756 25288 23808 25294
rect 23756 25230 23808 25236
rect 23480 24812 23532 24818
rect 23480 24754 23532 24760
rect 23388 24336 23440 24342
rect 23388 24278 23440 24284
rect 23020 24132 23072 24138
rect 23020 24074 23072 24080
rect 23032 23866 23060 24074
rect 23020 23860 23072 23866
rect 23020 23802 23072 23808
rect 23020 23248 23072 23254
rect 23020 23190 23072 23196
rect 23032 19378 23060 23190
rect 23400 23089 23428 24278
rect 23492 23118 23520 24754
rect 23584 24206 23612 25230
rect 23768 24818 23796 25230
rect 23756 24812 23808 24818
rect 23756 24754 23808 24760
rect 23664 24676 23716 24682
rect 23664 24618 23716 24624
rect 23676 24274 23704 24618
rect 23664 24268 23716 24274
rect 23664 24210 23716 24216
rect 23572 24200 23624 24206
rect 23572 24142 23624 24148
rect 23572 23792 23624 23798
rect 23572 23734 23624 23740
rect 23584 23526 23612 23734
rect 23676 23662 23704 24210
rect 23952 24138 23980 25638
rect 23940 24132 23992 24138
rect 23940 24074 23992 24080
rect 23952 23730 23980 24074
rect 23756 23724 23808 23730
rect 23756 23666 23808 23672
rect 23940 23724 23992 23730
rect 23940 23666 23992 23672
rect 23664 23656 23716 23662
rect 23664 23598 23716 23604
rect 23572 23520 23624 23526
rect 23572 23462 23624 23468
rect 23768 23322 23796 23666
rect 23756 23316 23808 23322
rect 23756 23258 23808 23264
rect 23768 23118 23796 23258
rect 23480 23112 23532 23118
rect 23386 23080 23442 23089
rect 23480 23054 23532 23060
rect 23756 23112 23808 23118
rect 23756 23054 23808 23060
rect 23386 23015 23442 23024
rect 23492 22778 23520 23054
rect 23480 22772 23532 22778
rect 23480 22714 23532 22720
rect 23572 22636 23624 22642
rect 23572 22578 23624 22584
rect 24032 22636 24084 22642
rect 24032 22578 24084 22584
rect 23112 22228 23164 22234
rect 23112 22170 23164 22176
rect 23124 22137 23152 22170
rect 23110 22128 23166 22137
rect 23110 22063 23166 22072
rect 23124 21690 23152 22063
rect 23584 21894 23612 22578
rect 23664 22500 23716 22506
rect 23664 22442 23716 22448
rect 23676 22030 23704 22442
rect 23664 22024 23716 22030
rect 23664 21966 23716 21972
rect 23572 21888 23624 21894
rect 23572 21830 23624 21836
rect 23112 21684 23164 21690
rect 23112 21626 23164 21632
rect 23584 20942 23612 21830
rect 23676 21690 23704 21966
rect 23664 21684 23716 21690
rect 23664 21626 23716 21632
rect 24044 21604 24072 22578
rect 24136 21962 24164 26250
rect 24228 22642 24256 27814
rect 24320 23594 24348 28494
rect 24400 26376 24452 26382
rect 24400 26318 24452 26324
rect 24412 24818 24440 26318
rect 24492 25900 24544 25906
rect 24492 25842 24544 25848
rect 24504 25430 24532 25842
rect 24596 25838 24624 28494
rect 24780 28150 24808 28630
rect 24768 28144 24820 28150
rect 24768 28086 24820 28092
rect 25136 28076 25188 28082
rect 25136 28018 25188 28024
rect 25044 27872 25096 27878
rect 25044 27814 25096 27820
rect 25056 27538 25084 27814
rect 25044 27532 25096 27538
rect 25044 27474 25096 27480
rect 25148 27470 25176 28018
rect 25136 27464 25188 27470
rect 25136 27406 25188 27412
rect 24768 27056 24820 27062
rect 24768 26998 24820 27004
rect 24780 25974 24808 26998
rect 25148 26586 25176 27406
rect 25136 26580 25188 26586
rect 25136 26522 25188 26528
rect 24768 25968 24820 25974
rect 24768 25910 24820 25916
rect 24952 25900 25004 25906
rect 24952 25842 25004 25848
rect 24584 25832 24636 25838
rect 24584 25774 24636 25780
rect 24492 25424 24544 25430
rect 24492 25366 24544 25372
rect 24596 25294 24624 25774
rect 24584 25288 24636 25294
rect 24584 25230 24636 25236
rect 24400 24812 24452 24818
rect 24400 24754 24452 24760
rect 24596 24206 24624 25230
rect 24768 25220 24820 25226
rect 24768 25162 24820 25168
rect 24780 24274 24808 25162
rect 24964 24410 24992 25842
rect 25136 24812 25188 24818
rect 25136 24754 25188 24760
rect 25148 24410 25176 24754
rect 25332 24750 25360 33526
rect 25412 29776 25464 29782
rect 25412 29718 25464 29724
rect 25424 28218 25452 29718
rect 25412 28212 25464 28218
rect 25412 28154 25464 28160
rect 26160 27470 26188 37062
rect 26516 36848 26568 36854
rect 28080 36848 28132 36854
rect 26516 36790 26568 36796
rect 28078 36816 28080 36825
rect 28132 36816 28134 36825
rect 26424 36712 26476 36718
rect 26424 36654 26476 36660
rect 26436 36378 26464 36654
rect 26424 36372 26476 36378
rect 26424 36314 26476 36320
rect 26528 36174 26556 36790
rect 27896 36780 27948 36786
rect 28078 36751 28134 36760
rect 27896 36722 27948 36728
rect 27908 36310 27936 36722
rect 28644 36378 28672 37130
rect 28632 36372 28684 36378
rect 28632 36314 28684 36320
rect 27896 36304 27948 36310
rect 27896 36246 27948 36252
rect 26516 36168 26568 36174
rect 26516 36110 26568 36116
rect 27908 35290 27936 36246
rect 28448 36168 28500 36174
rect 28448 36110 28500 36116
rect 28632 36168 28684 36174
rect 28632 36110 28684 36116
rect 27988 35760 28040 35766
rect 27988 35702 28040 35708
rect 27896 35284 27948 35290
rect 27896 35226 27948 35232
rect 27908 34678 27936 35226
rect 28000 34950 28028 35702
rect 28356 35488 28408 35494
rect 28356 35430 28408 35436
rect 28368 35086 28396 35430
rect 28460 35290 28488 36110
rect 28644 35562 28672 36110
rect 28724 35828 28776 35834
rect 28724 35770 28776 35776
rect 28632 35556 28684 35562
rect 28632 35498 28684 35504
rect 28448 35284 28500 35290
rect 28448 35226 28500 35232
rect 28736 35086 28764 35770
rect 28356 35080 28408 35086
rect 28356 35022 28408 35028
rect 28724 35080 28776 35086
rect 28724 35022 28776 35028
rect 27988 34944 28040 34950
rect 27988 34886 28040 34892
rect 27896 34672 27948 34678
rect 27896 34614 27948 34620
rect 27804 34604 27856 34610
rect 27804 34546 27856 34552
rect 27620 34196 27672 34202
rect 27620 34138 27672 34144
rect 27632 33658 27660 34138
rect 27816 33930 27844 34546
rect 27908 34202 27936 34614
rect 28000 34474 28028 34886
rect 27988 34468 28040 34474
rect 27988 34410 28040 34416
rect 27896 34196 27948 34202
rect 27896 34138 27948 34144
rect 28368 34134 28396 35022
rect 28920 35018 28948 37266
rect 32232 37126 32260 39200
rect 34164 37262 34192 39200
rect 34934 37564 35242 37584
rect 34934 37562 34940 37564
rect 34996 37562 35020 37564
rect 35076 37562 35100 37564
rect 35156 37562 35180 37564
rect 35236 37562 35242 37564
rect 34996 37510 34998 37562
rect 35178 37510 35180 37562
rect 34934 37508 34940 37510
rect 34996 37508 35020 37510
rect 35076 37508 35100 37510
rect 35156 37508 35180 37510
rect 35236 37508 35242 37510
rect 34934 37488 35242 37508
rect 36096 37346 36124 39200
rect 37556 37664 37608 37670
rect 37556 37606 37608 37612
rect 37568 37466 37596 37606
rect 37556 37460 37608 37466
rect 37556 37402 37608 37408
rect 37648 37460 37700 37466
rect 37648 37402 37700 37408
rect 36096 37318 36216 37346
rect 36188 37262 36216 37318
rect 32588 37256 32640 37262
rect 32588 37198 32640 37204
rect 34152 37256 34204 37262
rect 34152 37198 34204 37204
rect 35808 37256 35860 37262
rect 35808 37198 35860 37204
rect 36176 37256 36228 37262
rect 36176 37198 36228 37204
rect 37188 37256 37240 37262
rect 37188 37198 37240 37204
rect 32220 37120 32272 37126
rect 32220 37062 32272 37068
rect 32404 36916 32456 36922
rect 32404 36858 32456 36864
rect 31300 36780 31352 36786
rect 31300 36722 31352 36728
rect 30840 36644 30892 36650
rect 30840 36586 30892 36592
rect 29092 36576 29144 36582
rect 29092 36518 29144 36524
rect 30196 36576 30248 36582
rect 30196 36518 30248 36524
rect 29104 36174 29132 36518
rect 29092 36168 29144 36174
rect 29092 36110 29144 36116
rect 29104 35630 29132 36110
rect 29644 36032 29696 36038
rect 29644 35974 29696 35980
rect 29656 35698 29684 35974
rect 30208 35698 30236 36518
rect 30852 36174 30880 36586
rect 31312 36174 31340 36722
rect 31576 36712 31628 36718
rect 31576 36654 31628 36660
rect 31588 36378 31616 36654
rect 31576 36372 31628 36378
rect 31576 36314 31628 36320
rect 32416 36174 32444 36858
rect 32496 36576 32548 36582
rect 32496 36518 32548 36524
rect 32508 36242 32536 36518
rect 32496 36236 32548 36242
rect 32496 36178 32548 36184
rect 30840 36168 30892 36174
rect 30840 36110 30892 36116
rect 31300 36168 31352 36174
rect 31300 36110 31352 36116
rect 32404 36168 32456 36174
rect 32404 36110 32456 36116
rect 31760 36032 31812 36038
rect 31760 35974 31812 35980
rect 31772 35698 31800 35974
rect 32416 35698 32444 36110
rect 29644 35692 29696 35698
rect 29644 35634 29696 35640
rect 30196 35692 30248 35698
rect 30196 35634 30248 35640
rect 31760 35692 31812 35698
rect 31760 35634 31812 35640
rect 32404 35692 32456 35698
rect 32404 35634 32456 35640
rect 29092 35624 29144 35630
rect 29092 35566 29144 35572
rect 30208 35494 30236 35634
rect 30196 35488 30248 35494
rect 30196 35430 30248 35436
rect 28908 35012 28960 35018
rect 28908 34954 28960 34960
rect 28448 34604 28500 34610
rect 28448 34546 28500 34552
rect 28460 34406 28488 34546
rect 28448 34400 28500 34406
rect 28448 34342 28500 34348
rect 28356 34128 28408 34134
rect 28356 34070 28408 34076
rect 28264 33992 28316 33998
rect 28264 33934 28316 33940
rect 27712 33924 27764 33930
rect 27712 33866 27764 33872
rect 27804 33924 27856 33930
rect 27804 33866 27856 33872
rect 27620 33652 27672 33658
rect 27620 33594 27672 33600
rect 27724 33522 27752 33866
rect 27816 33658 27844 33866
rect 28080 33856 28132 33862
rect 28080 33798 28132 33804
rect 27804 33652 27856 33658
rect 27804 33594 27856 33600
rect 27712 33516 27764 33522
rect 27712 33458 27764 33464
rect 26332 33380 26384 33386
rect 26332 33322 26384 33328
rect 26344 32978 26372 33322
rect 27988 33312 28040 33318
rect 27988 33254 28040 33260
rect 28000 33114 28028 33254
rect 27988 33108 28040 33114
rect 27988 33050 28040 33056
rect 26332 32972 26384 32978
rect 26332 32914 26384 32920
rect 27988 32904 28040 32910
rect 28092 32892 28120 33798
rect 28276 32978 28304 33934
rect 28368 33454 28396 34070
rect 28460 33590 28488 34342
rect 28540 34196 28592 34202
rect 28540 34138 28592 34144
rect 28448 33584 28500 33590
rect 28448 33526 28500 33532
rect 28356 33448 28408 33454
rect 28356 33390 28408 33396
rect 28552 33318 28580 34138
rect 28908 33584 28960 33590
rect 28908 33526 28960 33532
rect 28632 33516 28684 33522
rect 28632 33458 28684 33464
rect 28540 33312 28592 33318
rect 28540 33254 28592 33260
rect 28644 33114 28672 33458
rect 28632 33108 28684 33114
rect 28632 33050 28684 33056
rect 28264 32972 28316 32978
rect 28264 32914 28316 32920
rect 28040 32864 28120 32892
rect 27988 32846 28040 32852
rect 27528 32836 27580 32842
rect 27528 32778 27580 32784
rect 26976 32768 27028 32774
rect 26976 32710 27028 32716
rect 26884 31884 26936 31890
rect 26884 31826 26936 31832
rect 26700 31272 26752 31278
rect 26700 31214 26752 31220
rect 26148 27464 26200 27470
rect 26148 27406 26200 27412
rect 26240 27328 26292 27334
rect 26240 27270 26292 27276
rect 26252 27062 26280 27270
rect 26240 27056 26292 27062
rect 26240 26998 26292 27004
rect 26608 25152 26660 25158
rect 26608 25094 26660 25100
rect 26240 24812 26292 24818
rect 26240 24754 26292 24760
rect 25320 24744 25372 24750
rect 25320 24686 25372 24692
rect 25412 24744 25464 24750
rect 25412 24686 25464 24692
rect 24952 24404 25004 24410
rect 24952 24346 25004 24352
rect 25136 24404 25188 24410
rect 25136 24346 25188 24352
rect 24768 24268 24820 24274
rect 24768 24210 24820 24216
rect 24492 24200 24544 24206
rect 24492 24142 24544 24148
rect 24584 24200 24636 24206
rect 24584 24142 24636 24148
rect 24308 23588 24360 23594
rect 24308 23530 24360 23536
rect 24504 23322 24532 24142
rect 24584 24064 24636 24070
rect 24584 24006 24636 24012
rect 24858 24032 24914 24041
rect 24492 23316 24544 23322
rect 24492 23258 24544 23264
rect 24216 22636 24268 22642
rect 24216 22578 24268 22584
rect 24492 22636 24544 22642
rect 24492 22578 24544 22584
rect 24400 22432 24452 22438
rect 24400 22374 24452 22380
rect 24412 22030 24440 22374
rect 24400 22024 24452 22030
rect 24400 21966 24452 21972
rect 24124 21956 24176 21962
rect 24124 21898 24176 21904
rect 24216 21616 24268 21622
rect 24044 21576 24216 21604
rect 24504 21570 24532 22578
rect 24216 21558 24268 21564
rect 23756 21344 23808 21350
rect 23756 21286 23808 21292
rect 23572 20936 23624 20942
rect 23572 20878 23624 20884
rect 23204 19712 23256 19718
rect 23204 19654 23256 19660
rect 23020 19372 23072 19378
rect 23072 19320 23152 19334
rect 23020 19314 23152 19320
rect 23032 19310 23152 19314
rect 23032 19306 23164 19310
rect 23112 19304 23164 19306
rect 23112 19246 23164 19252
rect 23216 18766 23244 19654
rect 23388 19508 23440 19514
rect 23388 19450 23440 19456
rect 23296 19372 23348 19378
rect 23296 19314 23348 19320
rect 23308 19156 23336 19314
rect 23400 19281 23428 19450
rect 23480 19372 23532 19378
rect 23480 19314 23532 19320
rect 23386 19272 23442 19281
rect 23386 19207 23442 19216
rect 23388 19168 23440 19174
rect 23308 19128 23388 19156
rect 23388 19110 23440 19116
rect 23204 18760 23256 18766
rect 23204 18702 23256 18708
rect 23112 18420 23164 18426
rect 23112 18362 23164 18368
rect 23124 15434 23152 18362
rect 23216 17882 23244 18702
rect 23204 17876 23256 17882
rect 23204 17818 23256 17824
rect 23204 17536 23256 17542
rect 23204 17478 23256 17484
rect 23216 16046 23244 17478
rect 23296 17060 23348 17066
rect 23296 17002 23348 17008
rect 23308 16590 23336 17002
rect 23296 16584 23348 16590
rect 23296 16526 23348 16532
rect 23308 16114 23336 16526
rect 23400 16454 23428 19110
rect 23492 18970 23520 19314
rect 23480 18964 23532 18970
rect 23480 18906 23532 18912
rect 23480 18080 23532 18086
rect 23480 18022 23532 18028
rect 23768 18034 23796 21286
rect 24228 21078 24256 21558
rect 24320 21554 24532 21570
rect 24308 21548 24532 21554
rect 24360 21542 24532 21548
rect 24308 21490 24360 21496
rect 24320 21350 24348 21490
rect 24308 21344 24360 21350
rect 24308 21286 24360 21292
rect 24216 21072 24268 21078
rect 24216 21014 24268 21020
rect 24228 20534 24256 21014
rect 24320 20602 24348 21286
rect 24308 20596 24360 20602
rect 24308 20538 24360 20544
rect 24216 20528 24268 20534
rect 24216 20470 24268 20476
rect 24492 19372 24544 19378
rect 24596 19360 24624 24006
rect 24858 23967 24914 23976
rect 24768 23656 24820 23662
rect 24768 23598 24820 23604
rect 24780 23254 24808 23598
rect 24768 23248 24820 23254
rect 24768 23190 24820 23196
rect 24872 23118 24900 23967
rect 24964 23798 24992 24346
rect 25044 24200 25096 24206
rect 25044 24142 25096 24148
rect 24952 23792 25004 23798
rect 24952 23734 25004 23740
rect 25056 23730 25084 24142
rect 25044 23724 25096 23730
rect 25044 23666 25096 23672
rect 24860 23112 24912 23118
rect 24860 23054 24912 23060
rect 24952 22976 25004 22982
rect 25056 22964 25084 23666
rect 25424 23526 25452 24686
rect 26252 24682 26280 24754
rect 26240 24676 26292 24682
rect 26240 24618 26292 24624
rect 25596 24404 25648 24410
rect 25596 24346 25648 24352
rect 25412 23520 25464 23526
rect 25412 23462 25464 23468
rect 25004 22936 25084 22964
rect 24952 22918 25004 22924
rect 24768 22024 24820 22030
rect 24768 21966 24820 21972
rect 24780 21146 24808 21966
rect 24768 21140 24820 21146
rect 24768 21082 24820 21088
rect 24676 20936 24728 20942
rect 24676 20878 24728 20884
rect 24688 19446 24716 20878
rect 24676 19440 24728 19446
rect 24676 19382 24728 19388
rect 24544 19332 24624 19360
rect 24492 19314 24544 19320
rect 24308 19304 24360 19310
rect 24308 19246 24360 19252
rect 24216 18692 24268 18698
rect 24216 18634 24268 18640
rect 24124 18352 24176 18358
rect 24122 18320 24124 18329
rect 24176 18320 24178 18329
rect 24122 18255 24178 18264
rect 24228 18222 24256 18634
rect 24320 18290 24348 19246
rect 24492 18624 24544 18630
rect 24492 18566 24544 18572
rect 24308 18284 24360 18290
rect 24308 18226 24360 18232
rect 24216 18216 24268 18222
rect 24216 18158 24268 18164
rect 23492 17610 23520 18022
rect 23768 18006 24164 18034
rect 23756 17876 23808 17882
rect 23756 17818 23808 17824
rect 23768 17678 23796 17818
rect 23756 17672 23808 17678
rect 23756 17614 23808 17620
rect 23480 17604 23532 17610
rect 23480 17546 23532 17552
rect 23388 16448 23440 16454
rect 23388 16390 23440 16396
rect 23296 16108 23348 16114
rect 23296 16050 23348 16056
rect 23204 16040 23256 16046
rect 23204 15982 23256 15988
rect 23112 15428 23164 15434
rect 23112 15370 23164 15376
rect 23124 15094 23152 15370
rect 23112 15088 23164 15094
rect 23112 15030 23164 15036
rect 23308 15026 23336 16050
rect 23400 15502 23428 16390
rect 23492 15570 23520 17546
rect 23768 15638 23796 17614
rect 23848 17536 23900 17542
rect 23848 17478 23900 17484
rect 23860 16590 23888 17478
rect 24136 16590 24164 18006
rect 23848 16584 23900 16590
rect 23848 16526 23900 16532
rect 24124 16584 24176 16590
rect 24124 16526 24176 16532
rect 24136 16114 24164 16526
rect 24124 16108 24176 16114
rect 24124 16050 24176 16056
rect 23756 15632 23808 15638
rect 23756 15574 23808 15580
rect 23480 15564 23532 15570
rect 23480 15506 23532 15512
rect 23388 15496 23440 15502
rect 23388 15438 23440 15444
rect 23386 15328 23442 15337
rect 23386 15263 23442 15272
rect 23296 15020 23348 15026
rect 23296 14962 23348 14968
rect 23400 14074 23428 15263
rect 23572 15156 23624 15162
rect 23572 15098 23624 15104
rect 23584 14822 23612 15098
rect 24136 15042 24164 16050
rect 24228 15162 24256 18158
rect 24320 17202 24348 18226
rect 24308 17196 24360 17202
rect 24308 17138 24360 17144
rect 24504 16590 24532 18566
rect 24596 17610 24624 19332
rect 24688 17746 24716 19382
rect 24780 19378 24808 21082
rect 24964 19514 24992 22918
rect 25320 21888 25372 21894
rect 25320 21830 25372 21836
rect 25332 21554 25360 21830
rect 25608 21690 25636 24346
rect 25964 24064 26016 24070
rect 25964 24006 26016 24012
rect 25976 23798 26004 24006
rect 25964 23792 26016 23798
rect 25964 23734 26016 23740
rect 26424 23112 26476 23118
rect 26424 23054 26476 23060
rect 25596 21684 25648 21690
rect 25596 21626 25648 21632
rect 25044 21548 25096 21554
rect 25044 21490 25096 21496
rect 25136 21548 25188 21554
rect 25136 21490 25188 21496
rect 25320 21548 25372 21554
rect 25320 21490 25372 21496
rect 25412 21548 25464 21554
rect 25412 21490 25464 21496
rect 26332 21548 26384 21554
rect 26332 21490 26384 21496
rect 25056 21146 25084 21490
rect 25148 21350 25176 21490
rect 25136 21344 25188 21350
rect 25136 21286 25188 21292
rect 25044 21140 25096 21146
rect 25044 21082 25096 21088
rect 25424 20942 25452 21490
rect 25688 21480 25740 21486
rect 25688 21422 25740 21428
rect 25700 20942 25728 21422
rect 25964 21344 26016 21350
rect 25964 21286 26016 21292
rect 25412 20936 25464 20942
rect 25412 20878 25464 20884
rect 25688 20936 25740 20942
rect 25688 20878 25740 20884
rect 25320 20800 25372 20806
rect 25320 20742 25372 20748
rect 25332 20534 25360 20742
rect 25700 20534 25728 20878
rect 25976 20874 26004 21286
rect 25964 20868 26016 20874
rect 25964 20810 26016 20816
rect 26240 20800 26292 20806
rect 26240 20742 26292 20748
rect 25320 20528 25372 20534
rect 25320 20470 25372 20476
rect 25688 20528 25740 20534
rect 25688 20470 25740 20476
rect 25964 20256 26016 20262
rect 25964 20198 26016 20204
rect 26056 20256 26108 20262
rect 26056 20198 26108 20204
rect 25976 19786 26004 20198
rect 26068 20058 26096 20198
rect 26056 20052 26108 20058
rect 26056 19994 26108 20000
rect 25964 19780 26016 19786
rect 25964 19722 26016 19728
rect 24952 19508 25004 19514
rect 24952 19450 25004 19456
rect 24768 19372 24820 19378
rect 24768 19314 24820 19320
rect 24780 17814 24808 19314
rect 24964 18408 24992 19450
rect 25688 18760 25740 18766
rect 25688 18702 25740 18708
rect 24872 18380 24992 18408
rect 24768 17808 24820 17814
rect 24768 17750 24820 17756
rect 24676 17740 24728 17746
rect 24676 17682 24728 17688
rect 24584 17604 24636 17610
rect 24584 17546 24636 17552
rect 24596 17338 24624 17546
rect 24584 17332 24636 17338
rect 24584 17274 24636 17280
rect 24688 17270 24716 17682
rect 24872 17678 24900 18380
rect 25044 18352 25096 18358
rect 25042 18320 25044 18329
rect 25096 18320 25098 18329
rect 24952 18284 25004 18290
rect 25042 18255 25098 18264
rect 24952 18226 25004 18232
rect 24964 17882 24992 18226
rect 24952 17876 25004 17882
rect 24952 17818 25004 17824
rect 24860 17672 24912 17678
rect 24860 17614 24912 17620
rect 24872 17270 24900 17614
rect 24952 17604 25004 17610
rect 24952 17546 25004 17552
rect 24676 17264 24728 17270
rect 24676 17206 24728 17212
rect 24860 17264 24912 17270
rect 24860 17206 24912 17212
rect 24492 16584 24544 16590
rect 24492 16526 24544 16532
rect 24504 15910 24532 16526
rect 24964 16114 24992 17546
rect 25056 16182 25084 18255
rect 25700 18086 25728 18702
rect 25688 18080 25740 18086
rect 25688 18022 25740 18028
rect 25976 17610 26004 19722
rect 26252 19310 26280 20742
rect 26344 19854 26372 21490
rect 26332 19848 26384 19854
rect 26332 19790 26384 19796
rect 26240 19304 26292 19310
rect 26240 19246 26292 19252
rect 26252 18426 26280 19246
rect 26436 18766 26464 23054
rect 26516 21412 26568 21418
rect 26516 21354 26568 21360
rect 26528 20942 26556 21354
rect 26516 20936 26568 20942
rect 26516 20878 26568 20884
rect 26528 20602 26556 20878
rect 26516 20596 26568 20602
rect 26516 20538 26568 20544
rect 26514 20224 26570 20233
rect 26514 20159 26570 20168
rect 26528 20058 26556 20159
rect 26516 20052 26568 20058
rect 26516 19994 26568 20000
rect 26528 19854 26556 19994
rect 26516 19848 26568 19854
rect 26516 19790 26568 19796
rect 26424 18760 26476 18766
rect 26424 18702 26476 18708
rect 26240 18420 26292 18426
rect 26240 18362 26292 18368
rect 26252 17746 26280 18362
rect 26240 17740 26292 17746
rect 26240 17682 26292 17688
rect 26424 17672 26476 17678
rect 26424 17614 26476 17620
rect 25964 17604 26016 17610
rect 25964 17546 26016 17552
rect 26332 17536 26384 17542
rect 26332 17478 26384 17484
rect 26344 17134 26372 17478
rect 26332 17128 26384 17134
rect 26238 17096 26294 17105
rect 26332 17070 26384 17076
rect 26238 17031 26294 17040
rect 25228 16992 25280 16998
rect 25228 16934 25280 16940
rect 25136 16448 25188 16454
rect 25136 16390 25188 16396
rect 25044 16176 25096 16182
rect 25044 16118 25096 16124
rect 24952 16108 25004 16114
rect 24952 16050 25004 16056
rect 24492 15904 24544 15910
rect 24492 15846 24544 15852
rect 24768 15904 24820 15910
rect 24768 15846 24820 15852
rect 24780 15745 24808 15846
rect 24766 15736 24822 15745
rect 24766 15671 24822 15680
rect 24308 15632 24360 15638
rect 24768 15632 24820 15638
rect 24360 15580 24440 15586
rect 24308 15574 24440 15580
rect 24768 15574 24820 15580
rect 24320 15558 24440 15574
rect 24412 15502 24440 15558
rect 24676 15564 24728 15570
rect 24676 15506 24728 15512
rect 24400 15496 24452 15502
rect 24400 15438 24452 15444
rect 24216 15156 24268 15162
rect 24216 15098 24268 15104
rect 24136 15014 24256 15042
rect 23572 14816 23624 14822
rect 23572 14758 23624 14764
rect 24124 14816 24176 14822
rect 24124 14758 24176 14764
rect 23388 14068 23440 14074
rect 23388 14010 23440 14016
rect 22836 13932 22888 13938
rect 22836 13874 22888 13880
rect 22928 13932 22980 13938
rect 22928 13874 22980 13880
rect 22848 13462 22876 13874
rect 23112 13728 23164 13734
rect 23112 13670 23164 13676
rect 22836 13456 22888 13462
rect 22836 13398 22888 13404
rect 22652 13252 22704 13258
rect 22652 13194 22704 13200
rect 22652 12436 22704 12442
rect 22652 12378 22704 12384
rect 22664 11762 22692 12378
rect 22848 11762 22876 13398
rect 23124 13394 23152 13670
rect 23112 13388 23164 13394
rect 23112 13330 23164 13336
rect 23020 13320 23072 13326
rect 23020 13262 23072 13268
rect 23032 12646 23060 13262
rect 23296 13252 23348 13258
rect 23296 13194 23348 13200
rect 23308 12986 23336 13194
rect 23296 12980 23348 12986
rect 23296 12922 23348 12928
rect 23020 12640 23072 12646
rect 23020 12582 23072 12588
rect 23478 12608 23534 12617
rect 23032 12481 23060 12582
rect 23478 12543 23534 12552
rect 23018 12472 23074 12481
rect 23018 12407 23074 12416
rect 23492 11801 23520 12543
rect 23584 11830 23612 14758
rect 23664 14272 23716 14278
rect 23664 14214 23716 14220
rect 23676 14006 23704 14214
rect 23664 14000 23716 14006
rect 23664 13942 23716 13948
rect 24136 13530 24164 14758
rect 24124 13524 24176 13530
rect 24124 13466 24176 13472
rect 23756 13456 23808 13462
rect 23756 13398 23808 13404
rect 23572 11824 23624 11830
rect 23478 11792 23534 11801
rect 22652 11756 22704 11762
rect 22652 11698 22704 11704
rect 22836 11756 22888 11762
rect 23572 11766 23624 11772
rect 23478 11727 23534 11736
rect 23664 11756 23716 11762
rect 22836 11698 22888 11704
rect 23664 11698 23716 11704
rect 22664 9926 22692 11698
rect 23296 11620 23348 11626
rect 23296 11562 23348 11568
rect 23020 11552 23072 11558
rect 23020 11494 23072 11500
rect 23032 11257 23060 11494
rect 23018 11248 23074 11257
rect 23018 11183 23074 11192
rect 22928 11008 22980 11014
rect 22928 10950 22980 10956
rect 22940 10674 22968 10950
rect 23308 10674 23336 11562
rect 23676 11082 23704 11698
rect 23664 11076 23716 11082
rect 23664 11018 23716 11024
rect 22928 10668 22980 10674
rect 22928 10610 22980 10616
rect 23296 10668 23348 10674
rect 23296 10610 23348 10616
rect 22652 9920 22704 9926
rect 22652 9862 22704 9868
rect 23308 9722 23336 10610
rect 23664 10600 23716 10606
rect 23664 10542 23716 10548
rect 23676 9994 23704 10542
rect 23388 9988 23440 9994
rect 23388 9930 23440 9936
rect 23664 9988 23716 9994
rect 23664 9930 23716 9936
rect 23296 9716 23348 9722
rect 23296 9658 23348 9664
rect 22928 9648 22980 9654
rect 22650 9616 22706 9625
rect 22928 9590 22980 9596
rect 22650 9551 22652 9560
rect 22704 9551 22706 9560
rect 22652 9522 22704 9528
rect 22940 8956 22968 9590
rect 23308 9586 23336 9658
rect 23400 9654 23428 9930
rect 23388 9648 23440 9654
rect 23388 9590 23440 9596
rect 23296 9580 23348 9586
rect 23296 9522 23348 9528
rect 23020 8968 23072 8974
rect 22940 8928 23020 8956
rect 22940 8566 22968 8928
rect 23020 8910 23072 8916
rect 23020 8832 23072 8838
rect 23020 8774 23072 8780
rect 22928 8560 22980 8566
rect 22928 8502 22980 8508
rect 23032 5778 23060 8774
rect 23400 8362 23428 9590
rect 23676 9586 23704 9930
rect 23664 9580 23716 9586
rect 23664 9522 23716 9528
rect 23388 8356 23440 8362
rect 23388 8298 23440 8304
rect 23572 7744 23624 7750
rect 23572 7686 23624 7692
rect 23584 7478 23612 7686
rect 23572 7472 23624 7478
rect 23572 7414 23624 7420
rect 23768 7410 23796 13398
rect 24124 13252 24176 13258
rect 24124 13194 24176 13200
rect 24032 12912 24084 12918
rect 24032 12854 24084 12860
rect 23940 11688 23992 11694
rect 23940 11630 23992 11636
rect 23952 10538 23980 11630
rect 23940 10532 23992 10538
rect 23940 10474 23992 10480
rect 24044 9897 24072 12854
rect 24136 10470 24164 13194
rect 24228 12238 24256 15014
rect 24412 13938 24440 15438
rect 24492 14340 24544 14346
rect 24492 14282 24544 14288
rect 24400 13932 24452 13938
rect 24400 13874 24452 13880
rect 24504 12850 24532 14282
rect 24688 12918 24716 15506
rect 24780 15026 24808 15574
rect 24860 15428 24912 15434
rect 24964 15416 24992 16050
rect 25044 16040 25096 16046
rect 25044 15982 25096 15988
rect 24912 15388 24992 15416
rect 24860 15370 24912 15376
rect 24768 15020 24820 15026
rect 24768 14962 24820 14968
rect 24964 14414 24992 15388
rect 25056 15094 25084 15982
rect 25044 15088 25096 15094
rect 25044 15030 25096 15036
rect 24952 14408 25004 14414
rect 24952 14350 25004 14356
rect 24768 13932 24820 13938
rect 24768 13874 24820 13880
rect 24676 12912 24728 12918
rect 24676 12854 24728 12860
rect 24492 12844 24544 12850
rect 24492 12786 24544 12792
rect 24216 12232 24268 12238
rect 24216 12174 24268 12180
rect 24228 11286 24256 12174
rect 24504 11762 24532 12786
rect 24688 12238 24716 12854
rect 24780 12850 24808 13874
rect 24952 13864 25004 13870
rect 24952 13806 25004 13812
rect 24860 13320 24912 13326
rect 24860 13262 24912 13268
rect 24872 12986 24900 13262
rect 24860 12980 24912 12986
rect 24860 12922 24912 12928
rect 24964 12850 24992 13806
rect 25056 13326 25084 15030
rect 25148 13734 25176 16390
rect 25240 15502 25268 16934
rect 26252 16250 26280 17031
rect 26436 16946 26464 17614
rect 26344 16918 26464 16946
rect 26240 16244 26292 16250
rect 26240 16186 26292 16192
rect 26344 16130 26372 16918
rect 26424 16584 26476 16590
rect 26424 16526 26476 16532
rect 26516 16584 26568 16590
rect 26516 16526 26568 16532
rect 26436 16250 26464 16526
rect 26424 16244 26476 16250
rect 26424 16186 26476 16192
rect 26528 16182 26556 16526
rect 26252 16102 26372 16130
rect 26516 16176 26568 16182
rect 26516 16118 26568 16124
rect 26252 15910 26280 16102
rect 26240 15904 26292 15910
rect 26240 15846 26292 15852
rect 26252 15570 26280 15846
rect 26240 15564 26292 15570
rect 26240 15506 26292 15512
rect 25228 15496 25280 15502
rect 25228 15438 25280 15444
rect 25136 13728 25188 13734
rect 25136 13670 25188 13676
rect 25044 13320 25096 13326
rect 25044 13262 25096 13268
rect 24768 12844 24820 12850
rect 24768 12786 24820 12792
rect 24952 12844 25004 12850
rect 24952 12786 25004 12792
rect 24676 12232 24728 12238
rect 24676 12174 24728 12180
rect 24492 11756 24544 11762
rect 24492 11698 24544 11704
rect 24216 11280 24268 11286
rect 24216 11222 24268 11228
rect 24398 10976 24454 10985
rect 24398 10911 24454 10920
rect 24412 10742 24440 10911
rect 24780 10810 24808 12786
rect 24964 11762 24992 12786
rect 25056 12782 25084 13262
rect 25148 13258 25176 13670
rect 25240 13326 25268 15438
rect 25872 15360 25924 15366
rect 25872 15302 25924 15308
rect 25884 15026 25912 15302
rect 26252 15094 26280 15506
rect 26240 15088 26292 15094
rect 26240 15030 26292 15036
rect 25872 15020 25924 15026
rect 25872 14962 25924 14968
rect 25596 14952 25648 14958
rect 25596 14894 25648 14900
rect 25608 13326 25636 14894
rect 26332 14340 26384 14346
rect 26332 14282 26384 14288
rect 26344 14074 26372 14282
rect 26240 14068 26292 14074
rect 26240 14010 26292 14016
rect 26332 14068 26384 14074
rect 26332 14010 26384 14016
rect 26252 13326 26280 14010
rect 25228 13320 25280 13326
rect 25228 13262 25280 13268
rect 25596 13320 25648 13326
rect 25596 13262 25648 13268
rect 26240 13320 26292 13326
rect 26240 13262 26292 13268
rect 25136 13252 25188 13258
rect 25136 13194 25188 13200
rect 25044 12776 25096 12782
rect 25044 12718 25096 12724
rect 25240 12345 25268 13262
rect 25608 12850 25636 13262
rect 25596 12844 25648 12850
rect 25596 12786 25648 12792
rect 25780 12708 25832 12714
rect 25780 12650 25832 12656
rect 25792 12434 25820 12650
rect 25700 12406 25820 12434
rect 25226 12336 25282 12345
rect 25226 12271 25282 12280
rect 25700 12238 25728 12406
rect 25688 12232 25740 12238
rect 25688 12174 25740 12180
rect 24952 11756 25004 11762
rect 24952 11698 25004 11704
rect 25228 11688 25280 11694
rect 25228 11630 25280 11636
rect 24768 10804 24820 10810
rect 24768 10746 24820 10752
rect 24308 10736 24360 10742
rect 24308 10678 24360 10684
rect 24400 10736 24452 10742
rect 24400 10678 24452 10684
rect 24320 10470 24348 10678
rect 25240 10674 25268 11630
rect 25596 11620 25648 11626
rect 25596 11562 25648 11568
rect 25320 11552 25372 11558
rect 25320 11494 25372 11500
rect 25332 11150 25360 11494
rect 25608 11354 25636 11562
rect 25596 11348 25648 11354
rect 25596 11290 25648 11296
rect 25700 11150 25728 12174
rect 25780 12096 25832 12102
rect 25780 12038 25832 12044
rect 25792 11830 25820 12038
rect 25780 11824 25832 11830
rect 25780 11766 25832 11772
rect 25964 11756 26016 11762
rect 25964 11698 26016 11704
rect 25320 11144 25372 11150
rect 25320 11086 25372 11092
rect 25688 11144 25740 11150
rect 25688 11086 25740 11092
rect 25976 10674 26004 11698
rect 26516 11212 26568 11218
rect 26516 11154 26568 11160
rect 25228 10668 25280 10674
rect 25228 10610 25280 10616
rect 25964 10668 26016 10674
rect 25964 10610 26016 10616
rect 25412 10600 25464 10606
rect 25464 10548 25544 10554
rect 25412 10542 25544 10548
rect 25424 10526 25544 10542
rect 24124 10464 24176 10470
rect 24124 10406 24176 10412
rect 24308 10464 24360 10470
rect 24308 10406 24360 10412
rect 24952 10464 25004 10470
rect 24952 10406 25004 10412
rect 24030 9888 24086 9897
rect 24030 9823 24086 9832
rect 24032 9648 24084 9654
rect 24032 9590 24084 9596
rect 24044 9353 24072 9590
rect 24216 9512 24268 9518
rect 24216 9454 24268 9460
rect 24030 9344 24086 9353
rect 24030 9279 24086 9288
rect 24228 9042 24256 9454
rect 24320 9450 24348 10406
rect 24964 10062 24992 10406
rect 25320 10260 25372 10266
rect 25320 10202 25372 10208
rect 24952 10056 25004 10062
rect 24952 9998 25004 10004
rect 24768 9920 24820 9926
rect 24768 9862 24820 9868
rect 24780 9586 24808 9862
rect 24676 9580 24728 9586
rect 24676 9522 24728 9528
rect 24768 9580 24820 9586
rect 24768 9522 24820 9528
rect 24308 9444 24360 9450
rect 24308 9386 24360 9392
rect 24688 9110 24716 9522
rect 24676 9104 24728 9110
rect 24676 9046 24728 9052
rect 24216 9036 24268 9042
rect 24216 8978 24268 8984
rect 24780 8498 24808 9522
rect 24860 9376 24912 9382
rect 24860 9318 24912 9324
rect 24872 9042 24900 9318
rect 24860 9036 24912 9042
rect 24860 8978 24912 8984
rect 25044 8968 25096 8974
rect 25044 8910 25096 8916
rect 25056 8566 25084 8910
rect 25044 8560 25096 8566
rect 25044 8502 25096 8508
rect 25332 8498 25360 10202
rect 25516 9994 25544 10526
rect 25976 9994 26004 10610
rect 26056 10464 26108 10470
rect 26056 10406 26108 10412
rect 25504 9988 25556 9994
rect 25504 9930 25556 9936
rect 25596 9988 25648 9994
rect 25596 9930 25648 9936
rect 25964 9988 26016 9994
rect 25964 9930 26016 9936
rect 25516 9586 25544 9930
rect 25608 9654 25636 9930
rect 25596 9648 25648 9654
rect 25596 9590 25648 9596
rect 25504 9580 25556 9586
rect 25504 9522 25556 9528
rect 25688 9580 25740 9586
rect 25688 9522 25740 9528
rect 25516 9178 25544 9522
rect 25700 9450 25728 9522
rect 26068 9518 26096 10406
rect 26528 10062 26556 11154
rect 26516 10056 26568 10062
rect 26516 9998 26568 10004
rect 26330 9616 26386 9625
rect 26528 9586 26556 9998
rect 26330 9551 26386 9560
rect 26516 9580 26568 9586
rect 26056 9512 26108 9518
rect 26056 9454 26108 9460
rect 25688 9444 25740 9450
rect 25688 9386 25740 9392
rect 25504 9172 25556 9178
rect 25504 9114 25556 9120
rect 25596 9104 25648 9110
rect 25596 9046 25648 9052
rect 24768 8492 24820 8498
rect 24768 8434 24820 8440
rect 25320 8492 25372 8498
rect 25320 8434 25372 8440
rect 25608 8430 25636 9046
rect 26068 8974 26096 9454
rect 26344 8974 26372 9551
rect 26516 9522 26568 9528
rect 26056 8968 26108 8974
rect 26056 8910 26108 8916
rect 26332 8968 26384 8974
rect 26332 8910 26384 8916
rect 25596 8424 25648 8430
rect 25596 8366 25648 8372
rect 23848 7948 23900 7954
rect 23848 7890 23900 7896
rect 23860 7750 23888 7890
rect 24216 7812 24268 7818
rect 24216 7754 24268 7760
rect 23848 7744 23900 7750
rect 23848 7686 23900 7692
rect 23664 7404 23716 7410
rect 23664 7346 23716 7352
rect 23756 7404 23808 7410
rect 23756 7346 23808 7352
rect 23296 7200 23348 7206
rect 23296 7142 23348 7148
rect 23020 5772 23072 5778
rect 23020 5714 23072 5720
rect 23308 5710 23336 7142
rect 23676 6458 23704 7346
rect 24228 6798 24256 7754
rect 26344 7478 26372 8910
rect 26516 8900 26568 8906
rect 26516 8842 26568 8848
rect 26528 8090 26556 8842
rect 26516 8084 26568 8090
rect 26516 8026 26568 8032
rect 26332 7472 26384 7478
rect 26332 7414 26384 7420
rect 25228 7200 25280 7206
rect 25228 7142 25280 7148
rect 25240 6798 25268 7142
rect 24216 6792 24268 6798
rect 24216 6734 24268 6740
rect 25228 6792 25280 6798
rect 25228 6734 25280 6740
rect 23664 6452 23716 6458
rect 23664 6394 23716 6400
rect 24228 6186 24256 6734
rect 25240 6390 25268 6734
rect 25228 6384 25280 6390
rect 25228 6326 25280 6332
rect 26240 6316 26292 6322
rect 26240 6258 26292 6264
rect 24216 6180 24268 6186
rect 24216 6122 24268 6128
rect 23296 5704 23348 5710
rect 24032 5704 24084 5710
rect 23348 5652 23520 5658
rect 23296 5646 23520 5652
rect 24032 5646 24084 5652
rect 23308 5630 23520 5646
rect 23388 5568 23440 5574
rect 23388 5510 23440 5516
rect 23400 5234 23428 5510
rect 23492 5302 23520 5630
rect 23480 5296 23532 5302
rect 23480 5238 23532 5244
rect 24044 5234 24072 5646
rect 24584 5636 24636 5642
rect 24584 5578 24636 5584
rect 24596 5302 24624 5578
rect 24768 5568 24820 5574
rect 24768 5510 24820 5516
rect 25320 5568 25372 5574
rect 25320 5510 25372 5516
rect 24584 5296 24636 5302
rect 24584 5238 24636 5244
rect 23388 5228 23440 5234
rect 23388 5170 23440 5176
rect 24032 5228 24084 5234
rect 24032 5170 24084 5176
rect 23400 4690 23428 5170
rect 23756 5024 23808 5030
rect 23756 4966 23808 4972
rect 23388 4684 23440 4690
rect 23388 4626 23440 4632
rect 23768 4214 23796 4966
rect 24780 4622 24808 5510
rect 25332 5166 25360 5510
rect 26148 5296 26200 5302
rect 26148 5238 26200 5244
rect 25320 5160 25372 5166
rect 25320 5102 25372 5108
rect 24768 4616 24820 4622
rect 24768 4558 24820 4564
rect 23756 4208 23808 4214
rect 23756 4150 23808 4156
rect 23388 4004 23440 4010
rect 23388 3946 23440 3952
rect 23400 3194 23428 3946
rect 23572 3936 23624 3942
rect 23572 3878 23624 3884
rect 23388 3188 23440 3194
rect 23388 3130 23440 3136
rect 23584 2922 23612 3878
rect 23768 3534 23796 4150
rect 24768 4140 24820 4146
rect 24768 4082 24820 4088
rect 24780 3602 24808 4082
rect 25872 4004 25924 4010
rect 25872 3946 25924 3952
rect 23940 3596 23992 3602
rect 23940 3538 23992 3544
rect 24768 3596 24820 3602
rect 24768 3538 24820 3544
rect 23756 3528 23808 3534
rect 23756 3470 23808 3476
rect 23756 3392 23808 3398
rect 23756 3334 23808 3340
rect 23664 2984 23716 2990
rect 23664 2926 23716 2932
rect 23572 2916 23624 2922
rect 23572 2858 23624 2864
rect 22560 2644 22612 2650
rect 22560 2586 22612 2592
rect 23676 2514 23704 2926
rect 23664 2508 23716 2514
rect 23664 2450 23716 2456
rect 23768 2446 23796 3334
rect 23952 3097 23980 3538
rect 24216 3392 24268 3398
rect 24216 3334 24268 3340
rect 24400 3392 24452 3398
rect 24400 3334 24452 3340
rect 24228 3126 24256 3334
rect 24216 3120 24268 3126
rect 23938 3088 23994 3097
rect 24216 3062 24268 3068
rect 24306 3088 24362 3097
rect 23938 3023 23994 3032
rect 23952 2774 23980 3023
rect 23860 2746 23980 2774
rect 23860 2650 23888 2746
rect 24228 2650 24256 3062
rect 24306 3023 24308 3032
rect 24360 3023 24362 3032
rect 24308 2994 24360 3000
rect 24412 2990 24440 3334
rect 24400 2984 24452 2990
rect 24400 2926 24452 2932
rect 23848 2644 23900 2650
rect 23848 2586 23900 2592
rect 24216 2644 24268 2650
rect 24216 2586 24268 2592
rect 25780 2508 25832 2514
rect 25780 2450 25832 2456
rect 15476 2440 15528 2446
rect 15476 2382 15528 2388
rect 18420 2440 18472 2446
rect 18420 2382 18472 2388
rect 19156 2440 19208 2446
rect 19156 2382 19208 2388
rect 20812 2440 20864 2446
rect 20812 2382 20864 2388
rect 21916 2440 21968 2446
rect 21916 2382 21968 2388
rect 23756 2440 23808 2446
rect 23756 2382 23808 2388
rect 14188 1896 14240 1902
rect 14188 1838 14240 1844
rect 15488 800 15516 2382
rect 18052 2304 18104 2310
rect 18052 2246 18104 2252
rect 18064 800 18092 2246
rect 18432 1970 18460 2382
rect 19984 2372 20036 2378
rect 19984 2314 20036 2320
rect 19574 2204 19882 2224
rect 19574 2202 19580 2204
rect 19636 2202 19660 2204
rect 19716 2202 19740 2204
rect 19796 2202 19820 2204
rect 19876 2202 19882 2204
rect 19636 2150 19638 2202
rect 19818 2150 19820 2202
rect 19574 2148 19580 2150
rect 19636 2148 19660 2150
rect 19716 2148 19740 2150
rect 19796 2148 19820 2150
rect 19876 2148 19882 2150
rect 19574 2128 19882 2148
rect 18420 1964 18472 1970
rect 18420 1906 18472 1912
rect 19996 800 20024 2314
rect 20168 2304 20220 2310
rect 20168 2246 20220 2252
rect 20180 1834 20208 2246
rect 20168 1828 20220 1834
rect 20168 1770 20220 1776
rect 21928 800 21956 2382
rect 23848 2372 23900 2378
rect 23848 2314 23900 2320
rect 23860 800 23888 2314
rect 25792 2258 25820 2450
rect 25884 2446 25912 3946
rect 26160 3738 26188 5238
rect 26148 3732 26200 3738
rect 26148 3674 26200 3680
rect 25964 3392 26016 3398
rect 25964 3334 26016 3340
rect 25976 2514 26004 3334
rect 26252 3074 26280 6258
rect 26424 4072 26476 4078
rect 26424 4014 26476 4020
rect 26436 3534 26464 4014
rect 26424 3528 26476 3534
rect 26424 3470 26476 3476
rect 26332 3392 26384 3398
rect 26332 3334 26384 3340
rect 26068 3046 26280 3074
rect 25964 2508 26016 2514
rect 25964 2450 26016 2456
rect 25872 2440 25924 2446
rect 25872 2382 25924 2388
rect 26068 2258 26096 3046
rect 26344 2990 26372 3334
rect 26148 2984 26200 2990
rect 26332 2984 26384 2990
rect 26200 2932 26280 2938
rect 26148 2926 26280 2932
rect 26332 2926 26384 2932
rect 26160 2910 26280 2926
rect 26252 2836 26280 2910
rect 26436 2836 26464 3470
rect 26252 2808 26464 2836
rect 26516 2848 26568 2854
rect 26344 2514 26372 2808
rect 26516 2790 26568 2796
rect 26332 2508 26384 2514
rect 26332 2450 26384 2456
rect 26528 2446 26556 2790
rect 26516 2440 26568 2446
rect 26516 2382 26568 2388
rect 25792 2230 26096 2258
rect 26620 1970 26648 25094
rect 26712 4690 26740 31214
rect 26896 30802 26924 31826
rect 26988 31822 27016 32710
rect 27540 32026 27568 32778
rect 27896 32768 27948 32774
rect 27896 32710 27948 32716
rect 27908 32230 27936 32710
rect 27896 32224 27948 32230
rect 27896 32166 27948 32172
rect 27068 32020 27120 32026
rect 27068 31962 27120 31968
rect 27528 32020 27580 32026
rect 27528 31962 27580 31968
rect 26976 31816 27028 31822
rect 26976 31758 27028 31764
rect 27080 31414 27108 31962
rect 27804 31816 27856 31822
rect 27804 31758 27856 31764
rect 27816 31414 27844 31758
rect 27908 31754 27936 32166
rect 28632 31884 28684 31890
rect 28632 31826 28684 31832
rect 27908 31726 28028 31754
rect 27068 31408 27120 31414
rect 27068 31350 27120 31356
rect 27804 31408 27856 31414
rect 27804 31350 27856 31356
rect 27816 30938 27844 31350
rect 27804 30932 27856 30938
rect 27804 30874 27856 30880
rect 26884 30796 26936 30802
rect 26884 30738 26936 30744
rect 26976 30728 27028 30734
rect 26976 30670 27028 30676
rect 26988 30394 27016 30670
rect 27712 30592 27764 30598
rect 27712 30534 27764 30540
rect 26976 30388 27028 30394
rect 26976 30330 27028 30336
rect 27068 30116 27120 30122
rect 27068 30058 27120 30064
rect 27080 29238 27108 30058
rect 27724 29646 27752 30534
rect 27804 29844 27856 29850
rect 27804 29786 27856 29792
rect 27712 29640 27764 29646
rect 27712 29582 27764 29588
rect 27160 29504 27212 29510
rect 27160 29446 27212 29452
rect 27068 29232 27120 29238
rect 27068 29174 27120 29180
rect 27172 29170 27200 29446
rect 27160 29164 27212 29170
rect 27160 29106 27212 29112
rect 27712 29028 27764 29034
rect 27712 28970 27764 28976
rect 27620 28960 27672 28966
rect 27620 28902 27672 28908
rect 27632 28694 27660 28902
rect 27620 28688 27672 28694
rect 27620 28630 27672 28636
rect 27724 28422 27752 28970
rect 27816 28626 27844 29786
rect 27896 29640 27948 29646
rect 27896 29582 27948 29588
rect 27908 28966 27936 29582
rect 27896 28960 27948 28966
rect 27896 28902 27948 28908
rect 27804 28620 27856 28626
rect 27804 28562 27856 28568
rect 27252 28416 27304 28422
rect 27252 28358 27304 28364
rect 27712 28416 27764 28422
rect 27712 28358 27764 28364
rect 27264 27674 27292 28358
rect 27804 28144 27856 28150
rect 27804 28086 27856 28092
rect 27252 27668 27304 27674
rect 27252 27610 27304 27616
rect 27436 27464 27488 27470
rect 27436 27406 27488 27412
rect 26884 27396 26936 27402
rect 26884 27338 26936 27344
rect 26896 26926 26924 27338
rect 27448 27062 27476 27406
rect 27436 27056 27488 27062
rect 27436 26998 27488 27004
rect 26884 26920 26936 26926
rect 26884 26862 26936 26868
rect 27712 25356 27764 25362
rect 27712 25298 27764 25304
rect 27620 25288 27672 25294
rect 27620 25230 27672 25236
rect 27632 24954 27660 25230
rect 27620 24948 27672 24954
rect 27620 24890 27672 24896
rect 27724 24818 27752 25298
rect 27712 24812 27764 24818
rect 27712 24754 27764 24760
rect 26792 24676 26844 24682
rect 26792 24618 26844 24624
rect 26804 23118 26832 24618
rect 27724 24410 27752 24754
rect 27816 24410 27844 28086
rect 27896 26784 27948 26790
rect 27896 26726 27948 26732
rect 27908 26382 27936 26726
rect 27896 26376 27948 26382
rect 27896 26318 27948 26324
rect 27712 24404 27764 24410
rect 27712 24346 27764 24352
rect 27804 24404 27856 24410
rect 27804 24346 27856 24352
rect 27712 23520 27764 23526
rect 27712 23462 27764 23468
rect 26792 23112 26844 23118
rect 26792 23054 26844 23060
rect 27724 22982 27752 23462
rect 27816 23118 27844 24346
rect 27804 23112 27856 23118
rect 27804 23054 27856 23060
rect 27712 22976 27764 22982
rect 27712 22918 27764 22924
rect 26792 21888 26844 21894
rect 26792 21830 26844 21836
rect 26804 21622 26832 21830
rect 26792 21616 26844 21622
rect 26792 21558 26844 21564
rect 27618 21584 27674 21593
rect 27618 21519 27674 21528
rect 27632 21078 27660 21519
rect 27620 21072 27672 21078
rect 27342 21040 27398 21049
rect 27620 21014 27672 21020
rect 27342 20975 27398 20984
rect 27356 20874 27384 20975
rect 27528 20936 27580 20942
rect 27632 20924 27660 21014
rect 27580 20896 27660 20924
rect 27528 20878 27580 20884
rect 27344 20868 27396 20874
rect 27344 20810 27396 20816
rect 27356 20534 27384 20810
rect 27344 20528 27396 20534
rect 27344 20470 27396 20476
rect 27160 19848 27212 19854
rect 27160 19790 27212 19796
rect 27172 18970 27200 19790
rect 27160 18964 27212 18970
rect 27160 18906 27212 18912
rect 27632 18902 27660 20896
rect 27724 20262 27752 22918
rect 27816 22166 27844 23054
rect 27804 22160 27856 22166
rect 27804 22102 27856 22108
rect 27816 21554 27844 22102
rect 28000 22094 28028 31726
rect 28356 31748 28408 31754
rect 28356 31690 28408 31696
rect 28368 31142 28396 31690
rect 28644 31346 28672 31826
rect 28632 31340 28684 31346
rect 28632 31282 28684 31288
rect 28356 31136 28408 31142
rect 28356 31078 28408 31084
rect 28368 29850 28396 31078
rect 28724 30728 28776 30734
rect 28724 30670 28776 30676
rect 28736 30598 28764 30670
rect 28724 30592 28776 30598
rect 28724 30534 28776 30540
rect 28736 30394 28764 30534
rect 28724 30388 28776 30394
rect 28724 30330 28776 30336
rect 28356 29844 28408 29850
rect 28356 29786 28408 29792
rect 28080 29640 28132 29646
rect 28080 29582 28132 29588
rect 28092 29170 28120 29582
rect 28172 29504 28224 29510
rect 28172 29446 28224 29452
rect 28184 29170 28212 29446
rect 28080 29164 28132 29170
rect 28080 29106 28132 29112
rect 28172 29164 28224 29170
rect 28172 29106 28224 29112
rect 28092 29050 28120 29106
rect 28264 29096 28316 29102
rect 28092 29044 28264 29050
rect 28092 29038 28316 29044
rect 28092 29022 28304 29038
rect 28276 28558 28304 29022
rect 28632 28960 28684 28966
rect 28632 28902 28684 28908
rect 28264 28552 28316 28558
rect 28264 28494 28316 28500
rect 28540 28416 28592 28422
rect 28540 28358 28592 28364
rect 28552 27470 28580 28358
rect 28080 27464 28132 27470
rect 28080 27406 28132 27412
rect 28540 27464 28592 27470
rect 28540 27406 28592 27412
rect 28092 26790 28120 27406
rect 28552 26994 28580 27406
rect 28644 27334 28672 28902
rect 28736 27334 28764 30330
rect 28632 27328 28684 27334
rect 28632 27270 28684 27276
rect 28724 27328 28776 27334
rect 28724 27270 28776 27276
rect 28644 27062 28672 27270
rect 28632 27056 28684 27062
rect 28632 26998 28684 27004
rect 28540 26988 28592 26994
rect 28540 26930 28592 26936
rect 28080 26784 28132 26790
rect 28080 26726 28132 26732
rect 28092 26330 28120 26726
rect 28092 26302 28212 26330
rect 28080 26240 28132 26246
rect 28080 26182 28132 26188
rect 28092 25906 28120 26182
rect 28184 26042 28212 26302
rect 28172 26036 28224 26042
rect 28172 25978 28224 25984
rect 28080 25900 28132 25906
rect 28080 25842 28132 25848
rect 28092 24818 28120 25842
rect 28184 25294 28212 25978
rect 28264 25832 28316 25838
rect 28264 25774 28316 25780
rect 28276 25362 28304 25774
rect 28264 25356 28316 25362
rect 28264 25298 28316 25304
rect 28172 25288 28224 25294
rect 28172 25230 28224 25236
rect 28724 25288 28776 25294
rect 28724 25230 28776 25236
rect 28080 24812 28132 24818
rect 28080 24754 28132 24760
rect 28540 24608 28592 24614
rect 28540 24550 28592 24556
rect 28552 24206 28580 24550
rect 28736 24410 28764 25230
rect 28724 24404 28776 24410
rect 28724 24346 28776 24352
rect 28540 24200 28592 24206
rect 28540 24142 28592 24148
rect 28816 24200 28868 24206
rect 28816 24142 28868 24148
rect 28828 23526 28856 24142
rect 28816 23520 28868 23526
rect 28816 23462 28868 23468
rect 28816 23112 28868 23118
rect 28816 23054 28868 23060
rect 28828 22778 28856 23054
rect 28816 22772 28868 22778
rect 28816 22714 28868 22720
rect 27908 22066 28028 22094
rect 27804 21548 27856 21554
rect 27804 21490 27856 21496
rect 27712 20256 27764 20262
rect 27712 20198 27764 20204
rect 27620 18896 27672 18902
rect 27620 18838 27672 18844
rect 27712 18896 27764 18902
rect 27712 18838 27764 18844
rect 27632 18698 27660 18838
rect 27724 18766 27752 18838
rect 27804 18828 27856 18834
rect 27804 18770 27856 18776
rect 27712 18760 27764 18766
rect 27712 18702 27764 18708
rect 27528 18692 27580 18698
rect 27528 18634 27580 18640
rect 27620 18692 27672 18698
rect 27620 18634 27672 18640
rect 27540 18578 27568 18634
rect 27816 18578 27844 18770
rect 27540 18550 27844 18578
rect 26976 18216 27028 18222
rect 26976 18158 27028 18164
rect 26988 18086 27016 18158
rect 26976 18080 27028 18086
rect 26976 18022 27028 18028
rect 26988 17610 27016 18022
rect 26976 17604 27028 17610
rect 26976 17546 27028 17552
rect 27620 17060 27672 17066
rect 27620 17002 27672 17008
rect 26792 16992 26844 16998
rect 26792 16934 26844 16940
rect 26804 16590 26832 16934
rect 26792 16584 26844 16590
rect 26792 16526 26844 16532
rect 26884 16448 26936 16454
rect 26884 16390 26936 16396
rect 26896 15706 26924 16390
rect 27632 16250 27660 17002
rect 27712 16652 27764 16658
rect 27712 16594 27764 16600
rect 27724 16250 27752 16594
rect 27620 16244 27672 16250
rect 27620 16186 27672 16192
rect 27712 16244 27764 16250
rect 27712 16186 27764 16192
rect 27252 16176 27304 16182
rect 27252 16118 27304 16124
rect 26884 15700 26936 15706
rect 26884 15642 26936 15648
rect 26896 15434 26924 15642
rect 26884 15428 26936 15434
rect 26884 15370 26936 15376
rect 26896 15026 26924 15370
rect 26884 15020 26936 15026
rect 26884 14962 26936 14968
rect 26896 14618 26924 14962
rect 26884 14612 26936 14618
rect 26936 14572 27016 14600
rect 26884 14554 26936 14560
rect 26988 12434 27016 14572
rect 27264 13190 27292 16118
rect 27436 16108 27488 16114
rect 27436 16050 27488 16056
rect 27448 15706 27476 16050
rect 27436 15700 27488 15706
rect 27436 15642 27488 15648
rect 27632 15162 27660 16186
rect 27620 15156 27672 15162
rect 27620 15098 27672 15104
rect 27344 14000 27396 14006
rect 27344 13942 27396 13948
rect 27068 13184 27120 13190
rect 27068 13126 27120 13132
rect 27252 13184 27304 13190
rect 27252 13126 27304 13132
rect 27080 12986 27108 13126
rect 27068 12980 27120 12986
rect 27068 12922 27120 12928
rect 26988 12406 27108 12434
rect 26882 10568 26938 10577
rect 26882 10503 26938 10512
rect 26896 9382 26924 10503
rect 26884 9376 26936 9382
rect 26884 9318 26936 9324
rect 26976 5704 27028 5710
rect 26976 5646 27028 5652
rect 26884 5636 26936 5642
rect 26884 5578 26936 5584
rect 26700 4684 26752 4690
rect 26700 4626 26752 4632
rect 26896 4554 26924 5578
rect 26988 5370 27016 5646
rect 26976 5364 27028 5370
rect 26976 5306 27028 5312
rect 26988 4690 27016 5306
rect 26976 4684 27028 4690
rect 26976 4626 27028 4632
rect 26884 4548 26936 4554
rect 26884 4490 26936 4496
rect 26976 3392 27028 3398
rect 26976 3334 27028 3340
rect 26884 3120 26936 3126
rect 26882 3088 26884 3097
rect 26936 3088 26938 3097
rect 26882 3023 26938 3032
rect 26884 2644 26936 2650
rect 26884 2586 26936 2592
rect 26896 2514 26924 2586
rect 26700 2508 26752 2514
rect 26700 2450 26752 2456
rect 26884 2508 26936 2514
rect 26884 2450 26936 2456
rect 26712 2378 26740 2450
rect 26988 2446 27016 3334
rect 27080 2650 27108 12406
rect 27356 9654 27384 13942
rect 27804 13796 27856 13802
rect 27804 13738 27856 13744
rect 27816 13326 27844 13738
rect 27804 13320 27856 13326
rect 27804 13262 27856 13268
rect 27436 12776 27488 12782
rect 27436 12718 27488 12724
rect 27448 10810 27476 12718
rect 27816 12434 27844 13262
rect 27724 12406 27844 12434
rect 27620 11756 27672 11762
rect 27620 11698 27672 11704
rect 27632 11558 27660 11698
rect 27620 11552 27672 11558
rect 27620 11494 27672 11500
rect 27632 11150 27660 11494
rect 27620 11144 27672 11150
rect 27620 11086 27672 11092
rect 27436 10804 27488 10810
rect 27436 10746 27488 10752
rect 27436 10192 27488 10198
rect 27436 10134 27488 10140
rect 27344 9648 27396 9654
rect 27344 9590 27396 9596
rect 27448 9518 27476 10134
rect 27632 10130 27660 11086
rect 27724 10606 27752 12406
rect 27804 11824 27856 11830
rect 27804 11766 27856 11772
rect 27816 11150 27844 11766
rect 27804 11144 27856 11150
rect 27804 11086 27856 11092
rect 27712 10600 27764 10606
rect 27712 10542 27764 10548
rect 27528 10124 27580 10130
rect 27528 10066 27580 10072
rect 27620 10124 27672 10130
rect 27620 10066 27672 10072
rect 27436 9512 27488 9518
rect 27436 9454 27488 9460
rect 27540 8974 27568 10066
rect 27724 9926 27752 10542
rect 27804 10532 27856 10538
rect 27804 10474 27856 10480
rect 27712 9920 27764 9926
rect 27712 9862 27764 9868
rect 27816 9081 27844 10474
rect 27802 9072 27858 9081
rect 27802 9007 27858 9016
rect 27252 8968 27304 8974
rect 27252 8910 27304 8916
rect 27528 8968 27580 8974
rect 27528 8910 27580 8916
rect 27264 8838 27292 8910
rect 27252 8832 27304 8838
rect 27252 8774 27304 8780
rect 27344 8832 27396 8838
rect 27344 8774 27396 8780
rect 27356 7886 27384 8774
rect 27540 8362 27568 8910
rect 27528 8356 27580 8362
rect 27528 8298 27580 8304
rect 27344 7880 27396 7886
rect 27344 7822 27396 7828
rect 27804 7880 27856 7886
rect 27804 7822 27856 7828
rect 27344 7744 27396 7750
rect 27396 7704 27476 7732
rect 27344 7686 27396 7692
rect 27160 7404 27212 7410
rect 27160 7346 27212 7352
rect 27172 7002 27200 7346
rect 27448 7274 27476 7704
rect 27816 7546 27844 7822
rect 27804 7540 27856 7546
rect 27804 7482 27856 7488
rect 27344 7268 27396 7274
rect 27344 7210 27396 7216
rect 27436 7268 27488 7274
rect 27436 7210 27488 7216
rect 27356 7002 27384 7210
rect 27620 7200 27672 7206
rect 27620 7142 27672 7148
rect 27160 6996 27212 7002
rect 27160 6938 27212 6944
rect 27344 6996 27396 7002
rect 27344 6938 27396 6944
rect 27344 6724 27396 6730
rect 27344 6666 27396 6672
rect 27356 5710 27384 6666
rect 27632 6390 27660 7142
rect 27804 6656 27856 6662
rect 27804 6598 27856 6604
rect 27620 6384 27672 6390
rect 27620 6326 27672 6332
rect 27816 6254 27844 6598
rect 27804 6248 27856 6254
rect 27804 6190 27856 6196
rect 27620 5840 27672 5846
rect 27620 5782 27672 5788
rect 27344 5704 27396 5710
rect 27344 5646 27396 5652
rect 27436 5228 27488 5234
rect 27436 5170 27488 5176
rect 27448 4690 27476 5170
rect 27632 5166 27660 5782
rect 27620 5160 27672 5166
rect 27620 5102 27672 5108
rect 27436 4684 27488 4690
rect 27436 4626 27488 4632
rect 27528 4004 27580 4010
rect 27528 3946 27580 3952
rect 27344 3120 27396 3126
rect 27344 3062 27396 3068
rect 27252 3052 27304 3058
rect 27252 2994 27304 3000
rect 27068 2644 27120 2650
rect 27068 2586 27120 2592
rect 26976 2440 27028 2446
rect 26976 2382 27028 2388
rect 26700 2372 26752 2378
rect 26700 2314 26752 2320
rect 26608 1964 26660 1970
rect 26608 1906 26660 1912
rect 26988 1766 27016 2382
rect 27264 2378 27292 2994
rect 27356 2922 27384 3062
rect 27344 2916 27396 2922
rect 27344 2858 27396 2864
rect 27252 2372 27304 2378
rect 27252 2314 27304 2320
rect 27540 1766 27568 3946
rect 27712 3392 27764 3398
rect 27712 3334 27764 3340
rect 27724 2446 27752 3334
rect 27908 2774 27936 22066
rect 27988 21616 28040 21622
rect 27988 21558 28040 21564
rect 28000 14482 28028 21558
rect 28816 21072 28868 21078
rect 28816 21014 28868 21020
rect 28080 20936 28132 20942
rect 28080 20878 28132 20884
rect 28092 19854 28120 20878
rect 28828 20874 28856 21014
rect 28816 20868 28868 20874
rect 28816 20810 28868 20816
rect 28264 20256 28316 20262
rect 28264 20198 28316 20204
rect 28276 19854 28304 20198
rect 28828 19854 28856 20810
rect 28080 19848 28132 19854
rect 28080 19790 28132 19796
rect 28264 19848 28316 19854
rect 28264 19790 28316 19796
rect 28816 19848 28868 19854
rect 28816 19790 28868 19796
rect 28092 19514 28120 19790
rect 28172 19780 28224 19786
rect 28172 19722 28224 19728
rect 28080 19508 28132 19514
rect 28080 19450 28132 19456
rect 28184 18290 28212 19722
rect 28172 18284 28224 18290
rect 28172 18226 28224 18232
rect 28632 17604 28684 17610
rect 28632 17546 28684 17552
rect 28356 17332 28408 17338
rect 28356 17274 28408 17280
rect 28172 17196 28224 17202
rect 28172 17138 28224 17144
rect 28080 16584 28132 16590
rect 28080 16526 28132 16532
rect 28092 16182 28120 16526
rect 28080 16176 28132 16182
rect 28080 16118 28132 16124
rect 28092 15094 28120 16118
rect 28184 16114 28212 17138
rect 28368 16658 28396 17274
rect 28448 17196 28500 17202
rect 28448 17138 28500 17144
rect 28460 17082 28488 17138
rect 28644 17082 28672 17546
rect 28724 17536 28776 17542
rect 28724 17478 28776 17484
rect 28736 17338 28764 17478
rect 28724 17332 28776 17338
rect 28724 17274 28776 17280
rect 28460 17054 28672 17082
rect 28356 16652 28408 16658
rect 28356 16594 28408 16600
rect 28644 16590 28672 17054
rect 28632 16584 28684 16590
rect 28632 16526 28684 16532
rect 28448 16516 28500 16522
rect 28448 16458 28500 16464
rect 28460 16182 28488 16458
rect 28448 16176 28500 16182
rect 28448 16118 28500 16124
rect 28172 16108 28224 16114
rect 28172 16050 28224 16056
rect 28080 15088 28132 15094
rect 28080 15030 28132 15036
rect 27988 14476 28040 14482
rect 27988 14418 28040 14424
rect 28092 14414 28120 15030
rect 28460 14618 28488 16118
rect 28540 15564 28592 15570
rect 28540 15506 28592 15512
rect 28448 14612 28500 14618
rect 28368 14572 28448 14600
rect 28080 14408 28132 14414
rect 28080 14350 28132 14356
rect 28368 14346 28396 14572
rect 28448 14554 28500 14560
rect 28460 14489 28488 14554
rect 28552 14414 28580 15506
rect 28644 15026 28672 16526
rect 28816 15156 28868 15162
rect 28816 15098 28868 15104
rect 28632 15020 28684 15026
rect 28632 14962 28684 14968
rect 28540 14408 28592 14414
rect 28540 14350 28592 14356
rect 28264 14340 28316 14346
rect 28264 14282 28316 14288
rect 28356 14340 28408 14346
rect 28356 14282 28408 14288
rect 27988 14272 28040 14278
rect 27988 14214 28040 14220
rect 28000 13326 28028 14214
rect 28276 13870 28304 14282
rect 28264 13864 28316 13870
rect 28264 13806 28316 13812
rect 27988 13320 28040 13326
rect 27988 13262 28040 13268
rect 28172 12776 28224 12782
rect 28172 12718 28224 12724
rect 28184 11762 28212 12718
rect 28276 11830 28304 13806
rect 28552 12850 28580 14350
rect 28644 14260 28672 14962
rect 28828 14414 28856 15098
rect 28816 14408 28868 14414
rect 28816 14350 28868 14356
rect 28644 14232 28856 14260
rect 28632 14068 28684 14074
rect 28632 14010 28684 14016
rect 28540 12844 28592 12850
rect 28540 12786 28592 12792
rect 28644 12306 28672 14010
rect 28724 13252 28776 13258
rect 28724 13194 28776 13200
rect 28632 12300 28684 12306
rect 28632 12242 28684 12248
rect 28264 11824 28316 11830
rect 28264 11766 28316 11772
rect 28172 11756 28224 11762
rect 28172 11698 28224 11704
rect 27988 11688 28040 11694
rect 27988 11630 28040 11636
rect 28000 11150 28028 11630
rect 27988 11144 28040 11150
rect 27988 11086 28040 11092
rect 28080 11008 28132 11014
rect 28080 10950 28132 10956
rect 28092 10674 28120 10950
rect 28080 10668 28132 10674
rect 28080 10610 28132 10616
rect 28736 10606 28764 13194
rect 28828 12782 28856 14232
rect 28816 12776 28868 12782
rect 28816 12718 28868 12724
rect 28828 12374 28856 12718
rect 28816 12368 28868 12374
rect 28816 12310 28868 12316
rect 28724 10600 28776 10606
rect 28724 10542 28776 10548
rect 28448 10056 28500 10062
rect 28448 9998 28500 10004
rect 28460 9674 28488 9998
rect 28460 9646 28580 9674
rect 28354 9344 28410 9353
rect 28354 9279 28410 9288
rect 28368 8820 28396 9279
rect 28552 8906 28580 9646
rect 28724 9648 28776 9654
rect 28724 9590 28776 9596
rect 28632 9580 28684 9586
rect 28632 9522 28684 9528
rect 28644 8974 28672 9522
rect 28632 8968 28684 8974
rect 28736 8952 28764 9590
rect 28920 9353 28948 33526
rect 30208 33318 30236 35430
rect 32600 35290 32628 37198
rect 34796 37188 34848 37194
rect 34796 37130 34848 37136
rect 35624 37188 35676 37194
rect 35624 37130 35676 37136
rect 34704 37120 34756 37126
rect 34704 37062 34756 37068
rect 34716 36786 34744 37062
rect 34808 36786 34836 37130
rect 35532 37120 35584 37126
rect 35532 37062 35584 37068
rect 35544 36786 35572 37062
rect 34704 36780 34756 36786
rect 34704 36722 34756 36728
rect 34796 36780 34848 36786
rect 34796 36722 34848 36728
rect 35532 36780 35584 36786
rect 35532 36722 35584 36728
rect 33416 36712 33468 36718
rect 33416 36654 33468 36660
rect 33428 36174 33456 36654
rect 33600 36644 33652 36650
rect 33600 36586 33652 36592
rect 33416 36168 33468 36174
rect 33416 36110 33468 36116
rect 33612 36106 33640 36586
rect 34808 36310 34836 36722
rect 34934 36476 35242 36496
rect 34934 36474 34940 36476
rect 34996 36474 35020 36476
rect 35076 36474 35100 36476
rect 35156 36474 35180 36476
rect 35236 36474 35242 36476
rect 34996 36422 34998 36474
rect 35178 36422 35180 36474
rect 34934 36420 34940 36422
rect 34996 36420 35020 36422
rect 35076 36420 35100 36422
rect 35156 36420 35180 36422
rect 35236 36420 35242 36422
rect 34934 36400 35242 36420
rect 35636 36310 35664 37130
rect 35820 36582 35848 37198
rect 37200 36922 37228 37198
rect 37188 36916 37240 36922
rect 37188 36858 37240 36864
rect 35808 36576 35860 36582
rect 35808 36518 35860 36524
rect 36452 36576 36504 36582
rect 36452 36518 36504 36524
rect 34796 36304 34848 36310
rect 34796 36246 34848 36252
rect 35624 36304 35676 36310
rect 35624 36246 35676 36252
rect 36464 36174 36492 36518
rect 34704 36168 34756 36174
rect 34704 36110 34756 36116
rect 36452 36168 36504 36174
rect 36452 36110 36504 36116
rect 33600 36100 33652 36106
rect 33600 36042 33652 36048
rect 33232 36032 33284 36038
rect 33232 35974 33284 35980
rect 33244 35698 33272 35974
rect 33232 35692 33284 35698
rect 33232 35634 33284 35640
rect 32588 35284 32640 35290
rect 32588 35226 32640 35232
rect 32404 34604 32456 34610
rect 32404 34546 32456 34552
rect 32772 34604 32824 34610
rect 32772 34546 32824 34552
rect 32416 33998 32444 34546
rect 32784 34202 32812 34546
rect 33612 34474 33640 36042
rect 34716 35222 34744 36110
rect 35532 36100 35584 36106
rect 35532 36042 35584 36048
rect 34934 35388 35242 35408
rect 34934 35386 34940 35388
rect 34996 35386 35020 35388
rect 35076 35386 35100 35388
rect 35156 35386 35180 35388
rect 35236 35386 35242 35388
rect 34996 35334 34998 35386
rect 35178 35334 35180 35386
rect 34934 35332 34940 35334
rect 34996 35332 35020 35334
rect 35076 35332 35100 35334
rect 35156 35332 35180 35334
rect 35236 35332 35242 35334
rect 34934 35312 35242 35332
rect 34704 35216 34756 35222
rect 34704 35158 34756 35164
rect 35348 35080 35400 35086
rect 35348 35022 35400 35028
rect 34796 34672 34848 34678
rect 34796 34614 34848 34620
rect 33600 34468 33652 34474
rect 33600 34410 33652 34416
rect 34808 34202 34836 34614
rect 35360 34542 35388 35022
rect 35348 34536 35400 34542
rect 35348 34478 35400 34484
rect 34934 34300 35242 34320
rect 34934 34298 34940 34300
rect 34996 34298 35020 34300
rect 35076 34298 35100 34300
rect 35156 34298 35180 34300
rect 35236 34298 35242 34300
rect 34996 34246 34998 34298
rect 35178 34246 35180 34298
rect 34934 34244 34940 34246
rect 34996 34244 35020 34246
rect 35076 34244 35100 34246
rect 35156 34244 35180 34246
rect 35236 34244 35242 34246
rect 34934 34224 35242 34244
rect 32772 34196 32824 34202
rect 32772 34138 32824 34144
rect 34796 34196 34848 34202
rect 34796 34138 34848 34144
rect 31116 33992 31168 33998
rect 31116 33934 31168 33940
rect 31392 33992 31444 33998
rect 31392 33934 31444 33940
rect 32404 33992 32456 33998
rect 32404 33934 32456 33940
rect 31128 33454 31156 33934
rect 31404 33658 31432 33934
rect 31392 33652 31444 33658
rect 31392 33594 31444 33600
rect 31208 33516 31260 33522
rect 31208 33458 31260 33464
rect 31116 33448 31168 33454
rect 31116 33390 31168 33396
rect 30196 33312 30248 33318
rect 30196 33254 30248 33260
rect 30472 32972 30524 32978
rect 30472 32914 30524 32920
rect 30484 32434 30512 32914
rect 30656 32904 30708 32910
rect 30656 32846 30708 32852
rect 30668 32434 30696 32846
rect 30472 32428 30524 32434
rect 30472 32370 30524 32376
rect 30656 32428 30708 32434
rect 30656 32370 30708 32376
rect 30484 31958 30512 32370
rect 30472 31952 30524 31958
rect 30472 31894 30524 31900
rect 30668 31890 30696 32370
rect 30656 31884 30708 31890
rect 30656 31826 30708 31832
rect 29736 31816 29788 31822
rect 29736 31758 29788 31764
rect 29092 31680 29144 31686
rect 29092 31622 29144 31628
rect 29104 31142 29132 31622
rect 29748 31346 29776 31758
rect 29736 31340 29788 31346
rect 29736 31282 29788 31288
rect 29092 31136 29144 31142
rect 29092 31078 29144 31084
rect 29104 30666 29132 31078
rect 30472 30796 30524 30802
rect 30472 30738 30524 30744
rect 29092 30660 29144 30666
rect 29092 30602 29144 30608
rect 30380 30320 30432 30326
rect 30380 30262 30432 30268
rect 30392 29850 30420 30262
rect 30380 29844 30432 29850
rect 30380 29786 30432 29792
rect 30392 29646 30420 29786
rect 30380 29640 30432 29646
rect 30380 29582 30432 29588
rect 29276 29028 29328 29034
rect 29276 28970 29328 28976
rect 29092 21344 29144 21350
rect 29092 21286 29144 21292
rect 29000 20528 29052 20534
rect 29000 20470 29052 20476
rect 29012 19922 29040 20470
rect 29104 20262 29132 21286
rect 29092 20256 29144 20262
rect 29092 20198 29144 20204
rect 29000 19916 29052 19922
rect 29000 19858 29052 19864
rect 29000 19440 29052 19446
rect 29000 19382 29052 19388
rect 29012 19242 29040 19382
rect 29000 19236 29052 19242
rect 29000 19178 29052 19184
rect 29000 18964 29052 18970
rect 29000 18906 29052 18912
rect 29012 18290 29040 18906
rect 29184 18760 29236 18766
rect 29184 18702 29236 18708
rect 29196 18426 29224 18702
rect 29184 18420 29236 18426
rect 29104 18380 29184 18408
rect 29000 18284 29052 18290
rect 29000 18226 29052 18232
rect 29104 16114 29132 18380
rect 29184 18362 29236 18368
rect 29184 16992 29236 16998
rect 29184 16934 29236 16940
rect 29196 16182 29224 16934
rect 29184 16176 29236 16182
rect 29184 16118 29236 16124
rect 29092 16108 29144 16114
rect 29092 16050 29144 16056
rect 29104 15706 29132 16050
rect 29092 15700 29144 15706
rect 29092 15642 29144 15648
rect 29104 15042 29132 15642
rect 29012 15014 29132 15042
rect 29012 14958 29040 15014
rect 29000 14952 29052 14958
rect 29000 14894 29052 14900
rect 29012 14006 29040 14894
rect 29000 14000 29052 14006
rect 29000 13942 29052 13948
rect 29184 12844 29236 12850
rect 29184 12786 29236 12792
rect 29196 11762 29224 12786
rect 29184 11756 29236 11762
rect 29184 11698 29236 11704
rect 29196 11218 29224 11698
rect 29184 11212 29236 11218
rect 29184 11154 29236 11160
rect 29092 9716 29144 9722
rect 29092 9658 29144 9664
rect 29000 9580 29052 9586
rect 29000 9522 29052 9528
rect 28906 9344 28962 9353
rect 28906 9279 28962 9288
rect 29012 9178 29040 9522
rect 29104 9178 29132 9658
rect 29000 9172 29052 9178
rect 29000 9114 29052 9120
rect 29092 9172 29144 9178
rect 29092 9114 29144 9120
rect 28632 8910 28684 8916
rect 28724 8946 28776 8952
rect 28540 8900 28592 8906
rect 28540 8842 28592 8848
rect 28368 8792 28488 8820
rect 28264 8628 28316 8634
rect 28264 8570 28316 8576
rect 28172 8560 28224 8566
rect 28172 8502 28224 8508
rect 27988 7744 28040 7750
rect 27988 7686 28040 7692
rect 28000 7410 28028 7686
rect 28184 7546 28212 8502
rect 28276 8090 28304 8570
rect 28264 8084 28316 8090
rect 28264 8026 28316 8032
rect 28276 7886 28304 8026
rect 28264 7880 28316 7886
rect 28264 7822 28316 7828
rect 28172 7540 28224 7546
rect 28172 7482 28224 7488
rect 28184 7410 28212 7482
rect 28276 7478 28304 7822
rect 28264 7472 28316 7478
rect 28264 7414 28316 7420
rect 27988 7404 28040 7410
rect 27988 7346 28040 7352
rect 28172 7404 28224 7410
rect 28172 7346 28224 7352
rect 27988 6724 28040 6730
rect 27988 6666 28040 6672
rect 28000 5914 28028 6666
rect 27988 5908 28040 5914
rect 27988 5850 28040 5856
rect 28356 3392 28408 3398
rect 28356 3334 28408 3340
rect 28368 3058 28396 3334
rect 28356 3052 28408 3058
rect 28356 2994 28408 3000
rect 27908 2746 28120 2774
rect 28092 2650 28120 2746
rect 28080 2644 28132 2650
rect 28080 2586 28132 2592
rect 28460 2446 28488 8792
rect 28552 8498 28580 8842
rect 28644 8786 28672 8910
rect 28724 8888 28776 8894
rect 28908 8900 28960 8906
rect 28908 8842 28960 8848
rect 28920 8786 28948 8842
rect 28644 8758 28948 8786
rect 29000 8560 29052 8566
rect 29104 8548 29132 9114
rect 29052 8520 29132 8548
rect 29000 8502 29052 8508
rect 28540 8492 28592 8498
rect 28540 8434 28592 8440
rect 28816 8492 28868 8498
rect 28816 8434 28868 8440
rect 28552 7818 28580 8434
rect 28828 7954 28856 8434
rect 28816 7948 28868 7954
rect 28816 7890 28868 7896
rect 28540 7812 28592 7818
rect 28540 7754 28592 7760
rect 29012 7410 29040 8502
rect 29000 7404 29052 7410
rect 29000 7346 29052 7352
rect 28908 7200 28960 7206
rect 28908 7142 28960 7148
rect 28920 3602 28948 7142
rect 29288 4010 29316 28970
rect 30380 28416 30432 28422
rect 30380 28358 30432 28364
rect 30392 28014 30420 28358
rect 30380 28008 30432 28014
rect 30380 27950 30432 27956
rect 30392 27878 30420 27950
rect 29644 27872 29696 27878
rect 29644 27814 29696 27820
rect 30380 27872 30432 27878
rect 30380 27814 30432 27820
rect 29656 27470 29684 27814
rect 29644 27464 29696 27470
rect 29644 27406 29696 27412
rect 29552 26784 29604 26790
rect 29552 26726 29604 26732
rect 29564 26518 29592 26726
rect 29552 26512 29604 26518
rect 29552 26454 29604 26460
rect 30392 25537 30420 27814
rect 30484 26926 30512 30738
rect 30932 30116 30984 30122
rect 30932 30058 30984 30064
rect 30840 29776 30892 29782
rect 30840 29718 30892 29724
rect 30656 29640 30708 29646
rect 30656 29582 30708 29588
rect 30564 27124 30616 27130
rect 30564 27066 30616 27072
rect 30472 26920 30524 26926
rect 30472 26862 30524 26868
rect 30576 26382 30604 27066
rect 30564 26376 30616 26382
rect 30564 26318 30616 26324
rect 30378 25528 30434 25537
rect 30378 25463 30434 25472
rect 30668 25430 30696 29582
rect 30748 28076 30800 28082
rect 30748 28018 30800 28024
rect 30760 27470 30788 28018
rect 30748 27464 30800 27470
rect 30748 27406 30800 27412
rect 30760 26382 30788 27406
rect 30748 26376 30800 26382
rect 30748 26318 30800 26324
rect 30760 25906 30788 26318
rect 30748 25900 30800 25906
rect 30748 25842 30800 25848
rect 30656 25424 30708 25430
rect 30656 25366 30708 25372
rect 29460 24064 29512 24070
rect 29460 24006 29512 24012
rect 29644 24064 29696 24070
rect 29644 24006 29696 24012
rect 29472 19174 29500 24006
rect 29656 23526 29684 24006
rect 29644 23520 29696 23526
rect 29642 23488 29644 23497
rect 29696 23488 29698 23497
rect 29642 23423 29698 23432
rect 30380 23112 30432 23118
rect 30380 23054 30432 23060
rect 30288 23044 30340 23050
rect 30288 22986 30340 22992
rect 29828 22976 29880 22982
rect 29828 22918 29880 22924
rect 29840 22642 29868 22918
rect 30300 22778 30328 22986
rect 30288 22772 30340 22778
rect 30288 22714 30340 22720
rect 30392 22642 30420 23054
rect 29828 22636 29880 22642
rect 29828 22578 29880 22584
rect 30380 22636 30432 22642
rect 30380 22578 30432 22584
rect 30852 22098 30880 29718
rect 30944 29714 30972 30058
rect 30932 29708 30984 29714
rect 30932 29650 30984 29656
rect 30932 29164 30984 29170
rect 30932 29106 30984 29112
rect 30944 27606 30972 29106
rect 30932 27600 30984 27606
rect 30932 27542 30984 27548
rect 31128 24750 31156 33390
rect 31220 32502 31248 33458
rect 31404 32978 31432 33594
rect 32416 33386 32444 33934
rect 35360 33930 35388 34478
rect 35440 33992 35492 33998
rect 35440 33934 35492 33940
rect 35348 33924 35400 33930
rect 35348 33866 35400 33872
rect 35452 33522 35480 33934
rect 35440 33516 35492 33522
rect 35440 33458 35492 33464
rect 32404 33380 32456 33386
rect 32404 33322 32456 33328
rect 34934 33212 35242 33232
rect 34934 33210 34940 33212
rect 34996 33210 35020 33212
rect 35076 33210 35100 33212
rect 35156 33210 35180 33212
rect 35236 33210 35242 33212
rect 34996 33158 34998 33210
rect 35178 33158 35180 33210
rect 34934 33156 34940 33158
rect 34996 33156 35020 33158
rect 35076 33156 35100 33158
rect 35156 33156 35180 33158
rect 35236 33156 35242 33158
rect 34934 33136 35242 33156
rect 31392 32972 31444 32978
rect 31392 32914 31444 32920
rect 34520 32904 34572 32910
rect 34520 32846 34572 32852
rect 33600 32768 33652 32774
rect 33600 32710 33652 32716
rect 33612 32570 33640 32710
rect 33600 32564 33652 32570
rect 33600 32506 33652 32512
rect 31208 32496 31260 32502
rect 31208 32438 31260 32444
rect 34532 32434 34560 32846
rect 35544 32774 35572 36042
rect 35992 35284 36044 35290
rect 35992 35226 36044 35232
rect 37372 35284 37424 35290
rect 37372 35226 37424 35232
rect 35900 35148 35952 35154
rect 35900 35090 35952 35096
rect 35912 34474 35940 35090
rect 36004 34950 36032 35226
rect 37188 35148 37240 35154
rect 37188 35090 37240 35096
rect 35992 34944 36044 34950
rect 35992 34886 36044 34892
rect 36004 34610 36032 34886
rect 35992 34604 36044 34610
rect 35992 34546 36044 34552
rect 35900 34468 35952 34474
rect 35900 34410 35952 34416
rect 35900 34060 35952 34066
rect 35900 34002 35952 34008
rect 35716 33652 35768 33658
rect 35716 33594 35768 33600
rect 35728 33318 35756 33594
rect 35912 33318 35940 34002
rect 37200 33998 37228 35090
rect 37384 33998 37412 35226
rect 37464 35080 37516 35086
rect 37464 35022 37516 35028
rect 37476 34542 37504 35022
rect 37464 34536 37516 34542
rect 37464 34478 37516 34484
rect 37188 33992 37240 33998
rect 37188 33934 37240 33940
rect 37372 33992 37424 33998
rect 37372 33934 37424 33940
rect 35716 33312 35768 33318
rect 35716 33254 35768 33260
rect 35900 33312 35952 33318
rect 35900 33254 35952 33260
rect 35912 32978 35940 33254
rect 35900 32972 35952 32978
rect 35900 32914 35952 32920
rect 35716 32904 35768 32910
rect 35716 32846 35768 32852
rect 37280 32904 37332 32910
rect 37280 32846 37332 32852
rect 35532 32768 35584 32774
rect 35532 32710 35584 32716
rect 35728 32502 35756 32846
rect 35716 32496 35768 32502
rect 35716 32438 35768 32444
rect 33784 32428 33836 32434
rect 33784 32370 33836 32376
rect 33968 32428 34020 32434
rect 33968 32370 34020 32376
rect 34520 32428 34572 32434
rect 34520 32370 34572 32376
rect 32128 31952 32180 31958
rect 32128 31894 32180 31900
rect 32140 31414 32168 31894
rect 32220 31748 32272 31754
rect 32220 31690 32272 31696
rect 32128 31408 32180 31414
rect 32128 31350 32180 31356
rect 32140 30870 32168 31350
rect 32232 31210 32260 31690
rect 33796 31482 33824 32370
rect 33980 32026 34008 32370
rect 34152 32360 34204 32366
rect 34152 32302 34204 32308
rect 34164 32026 34192 32302
rect 34934 32124 35242 32144
rect 34934 32122 34940 32124
rect 34996 32122 35020 32124
rect 35076 32122 35100 32124
rect 35156 32122 35180 32124
rect 35236 32122 35242 32124
rect 34996 32070 34998 32122
rect 35178 32070 35180 32122
rect 34934 32068 34940 32070
rect 34996 32068 35020 32070
rect 35076 32068 35100 32070
rect 35156 32068 35180 32070
rect 35236 32068 35242 32070
rect 34934 32048 35242 32068
rect 33968 32020 34020 32026
rect 33968 31962 34020 31968
rect 34152 32020 34204 32026
rect 34152 31962 34204 31968
rect 35728 31890 35756 32438
rect 37292 32434 37320 32846
rect 37464 32564 37516 32570
rect 37464 32506 37516 32512
rect 37280 32428 37332 32434
rect 37280 32370 37332 32376
rect 35716 31884 35768 31890
rect 35716 31826 35768 31832
rect 33968 31816 34020 31822
rect 33968 31758 34020 31764
rect 34152 31816 34204 31822
rect 34152 31758 34204 31764
rect 33784 31476 33836 31482
rect 33784 31418 33836 31424
rect 33980 31346 34008 31758
rect 33968 31340 34020 31346
rect 33968 31282 34020 31288
rect 32220 31204 32272 31210
rect 32220 31146 32272 31152
rect 32128 30864 32180 30870
rect 32128 30806 32180 30812
rect 32232 29306 32260 31146
rect 34164 30326 34192 31758
rect 34934 31036 35242 31056
rect 34934 31034 34940 31036
rect 34996 31034 35020 31036
rect 35076 31034 35100 31036
rect 35156 31034 35180 31036
rect 35236 31034 35242 31036
rect 34996 30982 34998 31034
rect 35178 30982 35180 31034
rect 34934 30980 34940 30982
rect 34996 30980 35020 30982
rect 35076 30980 35100 30982
rect 35156 30980 35180 30982
rect 35236 30980 35242 30982
rect 34934 30960 35242 30980
rect 34520 30728 34572 30734
rect 34520 30670 34572 30676
rect 37188 30728 37240 30734
rect 37188 30670 37240 30676
rect 34152 30320 34204 30326
rect 34152 30262 34204 30268
rect 32680 30252 32732 30258
rect 32680 30194 32732 30200
rect 34428 30252 34480 30258
rect 34428 30194 34480 30200
rect 32692 29714 32720 30194
rect 32772 30184 32824 30190
rect 32772 30126 32824 30132
rect 32956 30184 33008 30190
rect 32956 30126 33008 30132
rect 32784 29714 32812 30126
rect 32968 29850 32996 30126
rect 34440 30054 34468 30194
rect 34428 30048 34480 30054
rect 34428 29990 34480 29996
rect 32956 29844 33008 29850
rect 32956 29786 33008 29792
rect 32680 29708 32732 29714
rect 32680 29650 32732 29656
rect 32772 29708 32824 29714
rect 32772 29650 32824 29656
rect 32312 29504 32364 29510
rect 32312 29446 32364 29452
rect 32220 29300 32272 29306
rect 32220 29242 32272 29248
rect 32220 29164 32272 29170
rect 32220 29106 32272 29112
rect 31392 28484 31444 28490
rect 31392 28426 31444 28432
rect 31404 28082 31432 28426
rect 32232 28218 32260 29106
rect 32324 28694 32352 29446
rect 32692 29306 32720 29650
rect 32680 29300 32732 29306
rect 32680 29242 32732 29248
rect 33140 29096 33192 29102
rect 33140 29038 33192 29044
rect 32312 28688 32364 28694
rect 32312 28630 32364 28636
rect 32220 28212 32272 28218
rect 32220 28154 32272 28160
rect 31392 28076 31444 28082
rect 31392 28018 31444 28024
rect 32864 27600 32916 27606
rect 32864 27542 32916 27548
rect 32876 26994 32904 27542
rect 32864 26988 32916 26994
rect 32864 26930 32916 26936
rect 33152 26382 33180 29038
rect 33600 26784 33652 26790
rect 33600 26726 33652 26732
rect 33612 26382 33640 26726
rect 34440 26586 34468 29990
rect 34532 29170 34560 30670
rect 37200 30326 37228 30670
rect 37188 30320 37240 30326
rect 37188 30262 37240 30268
rect 34934 29948 35242 29968
rect 34934 29946 34940 29948
rect 34996 29946 35020 29948
rect 35076 29946 35100 29948
rect 35156 29946 35180 29948
rect 35236 29946 35242 29948
rect 34996 29894 34998 29946
rect 35178 29894 35180 29946
rect 34934 29892 34940 29894
rect 34996 29892 35020 29894
rect 35076 29892 35100 29894
rect 35156 29892 35180 29894
rect 35236 29892 35242 29894
rect 34934 29872 35242 29892
rect 37200 29850 37228 30262
rect 37188 29844 37240 29850
rect 37188 29786 37240 29792
rect 36452 29640 36504 29646
rect 36452 29582 36504 29588
rect 36636 29640 36688 29646
rect 36636 29582 36688 29588
rect 36464 29306 36492 29582
rect 36452 29300 36504 29306
rect 36452 29242 36504 29248
rect 34520 29164 34572 29170
rect 34520 29106 34572 29112
rect 34532 27538 34560 29106
rect 34934 28860 35242 28880
rect 34934 28858 34940 28860
rect 34996 28858 35020 28860
rect 35076 28858 35100 28860
rect 35156 28858 35180 28860
rect 35236 28858 35242 28860
rect 34996 28806 34998 28858
rect 35178 28806 35180 28858
rect 34934 28804 34940 28806
rect 34996 28804 35020 28806
rect 35076 28804 35100 28806
rect 35156 28804 35180 28806
rect 35236 28804 35242 28806
rect 34934 28784 35242 28804
rect 36648 28694 36676 29582
rect 36636 28688 36688 28694
rect 36636 28630 36688 28636
rect 34612 28620 34664 28626
rect 34612 28562 34664 28568
rect 34520 27532 34572 27538
rect 34520 27474 34572 27480
rect 34520 26920 34572 26926
rect 34520 26862 34572 26868
rect 34428 26580 34480 26586
rect 34428 26522 34480 26528
rect 33692 26444 33744 26450
rect 33692 26386 33744 26392
rect 33140 26376 33192 26382
rect 33140 26318 33192 26324
rect 33600 26376 33652 26382
rect 33600 26318 33652 26324
rect 31300 25356 31352 25362
rect 31300 25298 31352 25304
rect 31312 25265 31340 25298
rect 31392 25288 31444 25294
rect 31298 25256 31354 25265
rect 31392 25230 31444 25236
rect 31298 25191 31354 25200
rect 31404 24954 31432 25230
rect 31392 24948 31444 24954
rect 31392 24890 31444 24896
rect 31116 24744 31168 24750
rect 31116 24686 31168 24692
rect 33232 24608 33284 24614
rect 33232 24550 33284 24556
rect 31116 24404 31168 24410
rect 31116 24346 31168 24352
rect 31128 23662 31156 24346
rect 33244 24313 33272 24550
rect 33230 24304 33286 24313
rect 33230 24239 33286 24248
rect 31300 24064 31352 24070
rect 31300 24006 31352 24012
rect 31312 23866 31340 24006
rect 31300 23860 31352 23866
rect 31300 23802 31352 23808
rect 31116 23656 31168 23662
rect 31116 23598 31168 23604
rect 31128 23322 31156 23598
rect 31116 23316 31168 23322
rect 31116 23258 31168 23264
rect 31576 23112 31628 23118
rect 31576 23054 31628 23060
rect 30564 22094 30616 22098
rect 30840 22094 30892 22098
rect 30564 22092 30892 22094
rect 30616 22066 30840 22092
rect 30564 22034 30616 22040
rect 30840 22034 30892 22040
rect 29828 21888 29880 21894
rect 29828 21830 29880 21836
rect 29840 20942 29868 21830
rect 30564 21548 30616 21554
rect 30564 21490 30616 21496
rect 30380 21344 30432 21350
rect 30380 21286 30432 21292
rect 30392 20942 30420 21286
rect 30576 21185 30604 21490
rect 30562 21176 30618 21185
rect 30562 21111 30618 21120
rect 30748 21140 30800 21146
rect 30748 21082 30800 21088
rect 29552 20936 29604 20942
rect 29552 20878 29604 20884
rect 29644 20936 29696 20942
rect 29644 20878 29696 20884
rect 29828 20936 29880 20942
rect 29828 20878 29880 20884
rect 30380 20936 30432 20942
rect 30380 20878 30432 20884
rect 29564 20330 29592 20878
rect 29656 20602 29684 20878
rect 29644 20596 29696 20602
rect 29644 20538 29696 20544
rect 29644 20460 29696 20466
rect 29644 20402 29696 20408
rect 30104 20460 30156 20466
rect 30104 20402 30156 20408
rect 29552 20324 29604 20330
rect 29552 20266 29604 20272
rect 29656 20244 29684 20402
rect 29736 20256 29788 20262
rect 29656 20216 29736 20244
rect 29656 19786 29684 20216
rect 29736 20198 29788 20204
rect 29644 19780 29696 19786
rect 29644 19722 29696 19728
rect 29920 19712 29972 19718
rect 29920 19654 29972 19660
rect 29736 19508 29788 19514
rect 29736 19450 29788 19456
rect 29460 19168 29512 19174
rect 29460 19110 29512 19116
rect 29748 18766 29776 19450
rect 29932 18766 29960 19654
rect 30116 18766 30144 20402
rect 30392 20398 30420 20878
rect 30760 20466 30788 21082
rect 30852 20942 30880 22034
rect 31588 21690 31616 23054
rect 33508 22976 33560 22982
rect 33508 22918 33560 22924
rect 33520 22710 33548 22918
rect 33508 22704 33560 22710
rect 33506 22672 33508 22681
rect 33560 22672 33562 22681
rect 32956 22636 33008 22642
rect 33506 22607 33562 22616
rect 32956 22578 33008 22584
rect 33520 22581 33548 22607
rect 32680 21956 32732 21962
rect 32680 21898 32732 21904
rect 32692 21690 32720 21898
rect 32968 21690 32996 22578
rect 33324 22568 33376 22574
rect 33324 22510 33376 22516
rect 33336 21894 33364 22510
rect 33508 22500 33560 22506
rect 33508 22442 33560 22448
rect 33520 22166 33548 22442
rect 33612 22234 33640 26318
rect 33704 25430 33732 26386
rect 34532 25770 34560 26862
rect 34520 25764 34572 25770
rect 34520 25706 34572 25712
rect 34624 25430 34652 28562
rect 35348 28552 35400 28558
rect 35348 28494 35400 28500
rect 34934 27772 35242 27792
rect 34934 27770 34940 27772
rect 34996 27770 35020 27772
rect 35076 27770 35100 27772
rect 35156 27770 35180 27772
rect 35236 27770 35242 27772
rect 34996 27718 34998 27770
rect 35178 27718 35180 27770
rect 34934 27716 34940 27718
rect 34996 27716 35020 27718
rect 35076 27716 35100 27718
rect 35156 27716 35180 27718
rect 35236 27716 35242 27718
rect 34934 27696 35242 27716
rect 34704 27532 34756 27538
rect 34704 27474 34756 27480
rect 33692 25424 33744 25430
rect 33692 25366 33744 25372
rect 34612 25424 34664 25430
rect 34612 25366 34664 25372
rect 34716 25294 34744 27474
rect 35360 26994 35388 28494
rect 36360 28076 36412 28082
rect 36360 28018 36412 28024
rect 36452 28076 36504 28082
rect 36452 28018 36504 28024
rect 36372 27606 36400 28018
rect 36360 27600 36412 27606
rect 36360 27542 36412 27548
rect 36464 27470 36492 28018
rect 37292 27985 37320 32370
rect 37476 32366 37504 32506
rect 37464 32360 37516 32366
rect 37464 32302 37516 32308
rect 37372 31272 37424 31278
rect 37372 31214 37424 31220
rect 37384 30938 37412 31214
rect 37372 30932 37424 30938
rect 37372 30874 37424 30880
rect 37476 30818 37504 32302
rect 37556 31340 37608 31346
rect 37556 31282 37608 31288
rect 37384 30790 37504 30818
rect 37278 27976 37334 27985
rect 37278 27911 37334 27920
rect 36452 27464 36504 27470
rect 36452 27406 36504 27412
rect 36464 27130 36492 27406
rect 36452 27124 36504 27130
rect 36452 27066 36504 27072
rect 35348 26988 35400 26994
rect 35348 26930 35400 26936
rect 34796 26784 34848 26790
rect 34796 26726 34848 26732
rect 34808 26586 34836 26726
rect 34934 26684 35242 26704
rect 34934 26682 34940 26684
rect 34996 26682 35020 26684
rect 35076 26682 35100 26684
rect 35156 26682 35180 26684
rect 35236 26682 35242 26684
rect 34996 26630 34998 26682
rect 35178 26630 35180 26682
rect 34934 26628 34940 26630
rect 34996 26628 35020 26630
rect 35076 26628 35100 26630
rect 35156 26628 35180 26630
rect 35236 26628 35242 26630
rect 34934 26608 35242 26628
rect 34796 26580 34848 26586
rect 34796 26522 34848 26528
rect 34934 25596 35242 25616
rect 34934 25594 34940 25596
rect 34996 25594 35020 25596
rect 35076 25594 35100 25596
rect 35156 25594 35180 25596
rect 35236 25594 35242 25596
rect 34996 25542 34998 25594
rect 35178 25542 35180 25594
rect 34934 25540 34940 25542
rect 34996 25540 35020 25542
rect 35076 25540 35100 25542
rect 35156 25540 35180 25542
rect 35236 25540 35242 25542
rect 34934 25520 35242 25540
rect 34704 25288 34756 25294
rect 34704 25230 34756 25236
rect 34060 25152 34112 25158
rect 34060 25094 34112 25100
rect 34072 24886 34100 25094
rect 34716 24954 34744 25230
rect 34520 24948 34572 24954
rect 34520 24890 34572 24896
rect 34704 24948 34756 24954
rect 34704 24890 34756 24896
rect 34060 24880 34112 24886
rect 34060 24822 34112 24828
rect 33784 24812 33836 24818
rect 33784 24754 33836 24760
rect 33968 24812 34020 24818
rect 33968 24754 34020 24760
rect 33796 24070 33824 24754
rect 33876 24608 33928 24614
rect 33876 24550 33928 24556
rect 33888 24206 33916 24550
rect 33980 24410 34008 24754
rect 33968 24404 34020 24410
rect 33968 24346 34020 24352
rect 33876 24200 33928 24206
rect 33876 24142 33928 24148
rect 33784 24064 33836 24070
rect 33784 24006 33836 24012
rect 34336 24064 34388 24070
rect 34336 24006 34388 24012
rect 33600 22228 33652 22234
rect 33600 22170 33652 22176
rect 33508 22160 33560 22166
rect 33508 22102 33560 22108
rect 33048 21888 33100 21894
rect 33048 21830 33100 21836
rect 33324 21888 33376 21894
rect 33324 21830 33376 21836
rect 31576 21684 31628 21690
rect 31576 21626 31628 21632
rect 31668 21684 31720 21690
rect 31668 21626 31720 21632
rect 32680 21684 32732 21690
rect 32680 21626 32732 21632
rect 32956 21684 33008 21690
rect 32956 21626 33008 21632
rect 31680 21146 31708 21626
rect 31668 21140 31720 21146
rect 31668 21082 31720 21088
rect 31760 21140 31812 21146
rect 31760 21082 31812 21088
rect 31772 20942 31800 21082
rect 30840 20936 30892 20942
rect 30840 20878 30892 20884
rect 31760 20936 31812 20942
rect 31760 20878 31812 20884
rect 30748 20460 30800 20466
rect 30748 20402 30800 20408
rect 30852 20398 30880 20878
rect 31772 20602 31800 20878
rect 32680 20868 32732 20874
rect 32680 20810 32732 20816
rect 31760 20596 31812 20602
rect 31760 20538 31812 20544
rect 30380 20392 30432 20398
rect 30378 20360 30380 20369
rect 30840 20392 30892 20398
rect 30432 20360 30434 20369
rect 30840 20334 30892 20340
rect 30378 20295 30434 20304
rect 30392 20262 30420 20295
rect 30380 20256 30432 20262
rect 30380 20198 30432 20204
rect 30852 19922 30880 20334
rect 31760 20324 31812 20330
rect 31760 20266 31812 20272
rect 30840 19916 30892 19922
rect 30840 19858 30892 19864
rect 31772 19378 31800 20266
rect 31852 19780 31904 19786
rect 31852 19722 31904 19728
rect 31760 19372 31812 19378
rect 31760 19314 31812 19320
rect 31024 19304 31076 19310
rect 31024 19246 31076 19252
rect 31036 18970 31064 19246
rect 31392 19236 31444 19242
rect 31392 19178 31444 19184
rect 30656 18964 30708 18970
rect 30656 18906 30708 18912
rect 31024 18964 31076 18970
rect 31024 18906 31076 18912
rect 29736 18760 29788 18766
rect 29736 18702 29788 18708
rect 29920 18760 29972 18766
rect 29920 18702 29972 18708
rect 30104 18760 30156 18766
rect 30104 18702 30156 18708
rect 30196 18760 30248 18766
rect 30196 18702 30248 18708
rect 29644 18692 29696 18698
rect 29644 18634 29696 18640
rect 29368 18624 29420 18630
rect 29368 18566 29420 18572
rect 29380 18358 29408 18566
rect 29368 18352 29420 18358
rect 29368 18294 29420 18300
rect 29656 16114 29684 18634
rect 29932 17338 29960 18702
rect 30012 18080 30064 18086
rect 30012 18022 30064 18028
rect 29920 17332 29972 17338
rect 29920 17274 29972 17280
rect 30024 16998 30052 18022
rect 30116 17678 30144 18702
rect 30208 17882 30236 18702
rect 30668 18426 30696 18906
rect 31208 18896 31260 18902
rect 31208 18838 31260 18844
rect 30656 18420 30708 18426
rect 30656 18362 30708 18368
rect 30196 17876 30248 17882
rect 30196 17818 30248 17824
rect 30668 17678 30696 18362
rect 31024 18284 31076 18290
rect 31024 18226 31076 18232
rect 30104 17672 30156 17678
rect 30104 17614 30156 17620
rect 30656 17672 30708 17678
rect 30656 17614 30708 17620
rect 30840 17536 30892 17542
rect 30840 17478 30892 17484
rect 30852 17066 30880 17478
rect 31036 17202 31064 18226
rect 31024 17196 31076 17202
rect 31024 17138 31076 17144
rect 30840 17060 30892 17066
rect 30840 17002 30892 17008
rect 29828 16992 29880 16998
rect 29828 16934 29880 16940
rect 30012 16992 30064 16998
rect 30012 16934 30064 16940
rect 29840 16454 29868 16934
rect 30852 16658 30880 17002
rect 30840 16652 30892 16658
rect 30840 16594 30892 16600
rect 29828 16448 29880 16454
rect 29828 16390 29880 16396
rect 29644 16108 29696 16114
rect 29644 16050 29696 16056
rect 29656 15706 29684 16050
rect 29840 15910 29868 16390
rect 29828 15904 29880 15910
rect 29828 15846 29880 15852
rect 31022 15872 31078 15881
rect 29644 15700 29696 15706
rect 29644 15642 29696 15648
rect 29656 14362 29684 15642
rect 29656 14334 29776 14362
rect 29644 14272 29696 14278
rect 29644 14214 29696 14220
rect 29656 13326 29684 14214
rect 29748 14006 29776 14334
rect 29736 14000 29788 14006
rect 29736 13942 29788 13948
rect 29644 13320 29696 13326
rect 29644 13262 29696 13268
rect 29368 13184 29420 13190
rect 29368 13126 29420 13132
rect 29380 12850 29408 13126
rect 29368 12844 29420 12850
rect 29368 12786 29420 12792
rect 29460 12708 29512 12714
rect 29460 12650 29512 12656
rect 29368 11552 29420 11558
rect 29368 11494 29420 11500
rect 29380 10674 29408 11494
rect 29472 10810 29500 12650
rect 29644 12232 29696 12238
rect 29644 12174 29696 12180
rect 29656 11898 29684 12174
rect 29644 11892 29696 11898
rect 29644 11834 29696 11840
rect 29656 11762 29684 11834
rect 29644 11756 29696 11762
rect 29644 11698 29696 11704
rect 29840 11218 29868 15846
rect 31022 15807 31078 15816
rect 31036 15706 31064 15807
rect 31024 15700 31076 15706
rect 31024 15642 31076 15648
rect 30840 15632 30892 15638
rect 30840 15574 30892 15580
rect 30852 15026 30880 15574
rect 30932 15088 30984 15094
rect 30932 15030 30984 15036
rect 30012 15020 30064 15026
rect 30012 14962 30064 14968
rect 30840 15020 30892 15026
rect 30840 14962 30892 14968
rect 30024 14906 30052 14962
rect 29932 14878 30052 14906
rect 30104 14952 30156 14958
rect 30104 14894 30156 14900
rect 29932 14074 29960 14878
rect 30116 14618 30144 14894
rect 30840 14816 30892 14822
rect 30840 14758 30892 14764
rect 30104 14612 30156 14618
rect 30156 14572 30236 14600
rect 30104 14554 30156 14560
rect 29920 14068 29972 14074
rect 29920 14010 29972 14016
rect 30104 13932 30156 13938
rect 30104 13874 30156 13880
rect 30012 13320 30064 13326
rect 30012 13262 30064 13268
rect 30024 12306 30052 13262
rect 30012 12300 30064 12306
rect 30012 12242 30064 12248
rect 30116 12238 30144 13874
rect 30208 13326 30236 14572
rect 30564 14408 30616 14414
rect 30564 14350 30616 14356
rect 30196 13320 30248 13326
rect 30196 13262 30248 13268
rect 30286 13152 30342 13161
rect 30286 13087 30342 13096
rect 30300 12442 30328 13087
rect 30576 12850 30604 14350
rect 30564 12844 30616 12850
rect 30564 12786 30616 12792
rect 30196 12436 30248 12442
rect 30196 12378 30248 12384
rect 30288 12436 30340 12442
rect 30288 12378 30340 12384
rect 30104 12232 30156 12238
rect 30104 12174 30156 12180
rect 29920 12164 29972 12170
rect 29920 12106 29972 12112
rect 29932 11762 29960 12106
rect 30116 11898 30144 12174
rect 30104 11892 30156 11898
rect 30104 11834 30156 11840
rect 30208 11762 30236 12378
rect 29920 11756 29972 11762
rect 29920 11698 29972 11704
rect 30196 11756 30248 11762
rect 30196 11698 30248 11704
rect 29828 11212 29880 11218
rect 29828 11154 29880 11160
rect 29460 10804 29512 10810
rect 29460 10746 29512 10752
rect 29368 10668 29420 10674
rect 29368 10610 29420 10616
rect 29368 10124 29420 10130
rect 29368 10066 29420 10072
rect 29380 9654 29408 10066
rect 29472 9654 29500 10746
rect 29736 10668 29788 10674
rect 29736 10610 29788 10616
rect 29920 10668 29972 10674
rect 30208 10656 30236 11698
rect 30576 11694 30604 12786
rect 30656 12640 30708 12646
rect 30656 12582 30708 12588
rect 30668 12434 30696 12582
rect 30668 12406 30788 12434
rect 30656 12368 30708 12374
rect 30656 12310 30708 12316
rect 30668 11830 30696 12310
rect 30760 12102 30788 12406
rect 30852 12238 30880 14758
rect 30944 14346 30972 15030
rect 31036 14618 31064 15642
rect 31116 15020 31168 15026
rect 31116 14962 31168 14968
rect 31024 14612 31076 14618
rect 31024 14554 31076 14560
rect 31128 14550 31156 14962
rect 31116 14544 31168 14550
rect 31116 14486 31168 14492
rect 30932 14340 30984 14346
rect 30932 14282 30984 14288
rect 31116 14000 31168 14006
rect 31116 13942 31168 13948
rect 31128 13530 31156 13942
rect 31220 13530 31248 18838
rect 31404 18698 31432 19178
rect 31484 19168 31536 19174
rect 31484 19110 31536 19116
rect 31760 19168 31812 19174
rect 31760 19110 31812 19116
rect 31496 18902 31524 19110
rect 31484 18896 31536 18902
rect 31484 18838 31536 18844
rect 31392 18692 31444 18698
rect 31392 18634 31444 18640
rect 31300 18624 31352 18630
rect 31300 18566 31352 18572
rect 31312 17134 31340 18566
rect 31404 18290 31432 18634
rect 31772 18630 31800 19110
rect 31864 18766 31892 19722
rect 32692 19514 32720 20810
rect 32864 19780 32916 19786
rect 32864 19722 32916 19728
rect 32680 19508 32732 19514
rect 32680 19450 32732 19456
rect 32312 19304 32364 19310
rect 32312 19246 32364 19252
rect 31852 18760 31904 18766
rect 31852 18702 31904 18708
rect 32324 18698 32352 19246
rect 32876 18970 32904 19722
rect 32864 18964 32916 18970
rect 32864 18906 32916 18912
rect 32312 18692 32364 18698
rect 32312 18634 32364 18640
rect 31760 18624 31812 18630
rect 31760 18566 31812 18572
rect 32404 18624 32456 18630
rect 32404 18566 32456 18572
rect 31772 18358 31800 18566
rect 31760 18352 31812 18358
rect 31760 18294 31812 18300
rect 31392 18284 31444 18290
rect 31392 18226 31444 18232
rect 31484 18080 31536 18086
rect 31484 18022 31536 18028
rect 31300 17128 31352 17134
rect 31300 17070 31352 17076
rect 31392 16992 31444 16998
rect 31392 16934 31444 16940
rect 31404 16658 31432 16934
rect 31392 16652 31444 16658
rect 31392 16594 31444 16600
rect 31392 15360 31444 15366
rect 31392 15302 31444 15308
rect 31404 14385 31432 15302
rect 31496 14414 31524 18022
rect 32416 17678 32444 18566
rect 32876 18426 32904 18906
rect 33060 18578 33088 21830
rect 33336 21457 33364 21830
rect 33322 21448 33378 21457
rect 33322 21383 33378 21392
rect 33416 20528 33468 20534
rect 33416 20470 33468 20476
rect 33428 19786 33456 20470
rect 33508 20460 33560 20466
rect 33508 20402 33560 20408
rect 33520 19922 33548 20402
rect 33508 19916 33560 19922
rect 33508 19858 33560 19864
rect 33416 19780 33468 19786
rect 33416 19722 33468 19728
rect 33140 18624 33192 18630
rect 33060 18572 33140 18578
rect 33060 18566 33192 18572
rect 33060 18550 33180 18566
rect 32864 18420 32916 18426
rect 32864 18362 32916 18368
rect 33324 18284 33376 18290
rect 33324 18226 33376 18232
rect 33232 17876 33284 17882
rect 33232 17818 33284 17824
rect 32404 17672 32456 17678
rect 32404 17614 32456 17620
rect 32416 17202 32444 17614
rect 32588 17604 32640 17610
rect 32588 17546 32640 17552
rect 32404 17196 32456 17202
rect 32404 17138 32456 17144
rect 32496 16652 32548 16658
rect 32496 16594 32548 16600
rect 32508 16454 32536 16594
rect 32496 16448 32548 16454
rect 32496 16390 32548 16396
rect 32508 16250 32536 16390
rect 32496 16244 32548 16250
rect 32496 16186 32548 16192
rect 32036 15700 32088 15706
rect 32036 15642 32088 15648
rect 32404 15700 32456 15706
rect 32404 15642 32456 15648
rect 32048 15026 32076 15642
rect 32312 15496 32364 15502
rect 32312 15438 32364 15444
rect 32128 15360 32180 15366
rect 32128 15302 32180 15308
rect 32220 15360 32272 15366
rect 32220 15302 32272 15308
rect 32036 15020 32088 15026
rect 32036 14962 32088 14968
rect 32036 14816 32088 14822
rect 32036 14758 32088 14764
rect 32048 14414 32076 14758
rect 32140 14414 32168 15302
rect 32232 15094 32260 15302
rect 32220 15088 32272 15094
rect 32220 15030 32272 15036
rect 32232 14618 32260 15030
rect 32324 14890 32352 15438
rect 32416 15366 32444 15642
rect 32404 15360 32456 15366
rect 32404 15302 32456 15308
rect 32312 14884 32364 14890
rect 32312 14826 32364 14832
rect 32220 14612 32272 14618
rect 32220 14554 32272 14560
rect 31484 14408 31536 14414
rect 31390 14376 31446 14385
rect 31484 14350 31536 14356
rect 32036 14408 32088 14414
rect 32036 14350 32088 14356
rect 32128 14408 32180 14414
rect 32128 14350 32180 14356
rect 32312 14408 32364 14414
rect 32312 14350 32364 14356
rect 31390 14311 31446 14320
rect 31404 14278 31432 14311
rect 31392 14272 31444 14278
rect 31392 14214 31444 14220
rect 30932 13524 30984 13530
rect 30932 13466 30984 13472
rect 31116 13524 31168 13530
rect 31116 13466 31168 13472
rect 31208 13524 31260 13530
rect 31208 13466 31260 13472
rect 30840 12232 30892 12238
rect 30840 12174 30892 12180
rect 30748 12096 30800 12102
rect 30748 12038 30800 12044
rect 30656 11824 30708 11830
rect 30656 11766 30708 11772
rect 30564 11688 30616 11694
rect 30564 11630 30616 11636
rect 30380 11348 30432 11354
rect 30380 11290 30432 11296
rect 30288 11144 30340 11150
rect 30288 11086 30340 11092
rect 29972 10628 30236 10656
rect 29920 10610 29972 10616
rect 29748 10198 29776 10610
rect 30300 10470 30328 11086
rect 29828 10464 29880 10470
rect 29828 10406 29880 10412
rect 30288 10464 30340 10470
rect 30288 10406 30340 10412
rect 29736 10192 29788 10198
rect 29736 10134 29788 10140
rect 29748 9722 29776 10134
rect 29736 9716 29788 9722
rect 29736 9658 29788 9664
rect 29368 9648 29420 9654
rect 29368 9590 29420 9596
rect 29460 9648 29512 9654
rect 29460 9590 29512 9596
rect 29380 8634 29408 9590
rect 29460 9512 29512 9518
rect 29460 9454 29512 9460
rect 29472 8906 29500 9454
rect 29644 9104 29696 9110
rect 29644 9046 29696 9052
rect 29460 8900 29512 8906
rect 29460 8842 29512 8848
rect 29368 8628 29420 8634
rect 29368 8570 29420 8576
rect 29656 5778 29684 9046
rect 29748 8566 29776 9658
rect 29840 9625 29868 10406
rect 29920 9648 29972 9654
rect 29826 9616 29882 9625
rect 29920 9590 29972 9596
rect 29826 9551 29828 9560
rect 29880 9551 29882 9560
rect 29828 9522 29880 9528
rect 29840 9491 29868 9522
rect 29736 8560 29788 8566
rect 29736 8502 29788 8508
rect 29932 7886 29960 9590
rect 30300 8498 30328 10406
rect 30392 8634 30420 11290
rect 30760 10062 30788 12038
rect 30748 10056 30800 10062
rect 30748 9998 30800 10004
rect 30840 9920 30892 9926
rect 30840 9862 30892 9868
rect 30746 9616 30802 9625
rect 30746 9551 30802 9560
rect 30564 9376 30616 9382
rect 30564 9318 30616 9324
rect 30380 8628 30432 8634
rect 30380 8570 30432 8576
rect 30288 8492 30340 8498
rect 30288 8434 30340 8440
rect 30392 7954 30420 8570
rect 30380 7948 30432 7954
rect 30380 7890 30432 7896
rect 29920 7880 29972 7886
rect 29920 7822 29972 7828
rect 30576 7342 30604 9318
rect 30760 8906 30788 9551
rect 30852 8974 30880 9862
rect 30944 9042 30972 13466
rect 32048 13326 32076 14350
rect 32036 13320 32088 13326
rect 32036 13262 32088 13268
rect 31760 13184 31812 13190
rect 31760 13126 31812 13132
rect 31574 12472 31630 12481
rect 31574 12407 31630 12416
rect 31484 11552 31536 11558
rect 31484 11494 31536 11500
rect 31496 11150 31524 11494
rect 31484 11144 31536 11150
rect 31484 11086 31536 11092
rect 31484 10736 31536 10742
rect 31484 10678 31536 10684
rect 31024 10464 31076 10470
rect 31024 10406 31076 10412
rect 31036 9217 31064 10406
rect 31022 9208 31078 9217
rect 31022 9143 31078 9152
rect 30932 9036 30984 9042
rect 30932 8978 30984 8984
rect 30840 8968 30892 8974
rect 30840 8910 30892 8916
rect 30748 8900 30800 8906
rect 30748 8842 30800 8848
rect 31496 7546 31524 10678
rect 31588 10266 31616 12407
rect 31772 12238 31800 13126
rect 32048 12850 32076 13262
rect 32140 13258 32168 14350
rect 32324 14074 32352 14350
rect 32600 14226 32628 17546
rect 32956 17196 33008 17202
rect 32956 17138 33008 17144
rect 32680 16992 32732 16998
rect 32680 16934 32732 16940
rect 32692 16454 32720 16934
rect 32968 16590 32996 17138
rect 33048 16788 33100 16794
rect 33048 16730 33100 16736
rect 32956 16584 33008 16590
rect 32956 16526 33008 16532
rect 32680 16448 32732 16454
rect 32680 16390 32732 16396
rect 32692 15570 32720 16390
rect 33060 15609 33088 16730
rect 33046 15600 33102 15609
rect 32680 15564 32732 15570
rect 33046 15535 33102 15544
rect 32680 15506 32732 15512
rect 33140 15496 33192 15502
rect 33140 15438 33192 15444
rect 33152 15094 33180 15438
rect 33140 15088 33192 15094
rect 33140 15030 33192 15036
rect 32954 14376 33010 14385
rect 32954 14311 33010 14320
rect 32968 14278 32996 14311
rect 32508 14198 32628 14226
rect 32956 14272 33008 14278
rect 32956 14214 33008 14220
rect 32312 14068 32364 14074
rect 32312 14010 32364 14016
rect 32508 13938 32536 14198
rect 33244 14006 33272 17818
rect 33336 17660 33364 18226
rect 33428 17882 33456 19722
rect 34348 19378 34376 24006
rect 34532 22506 34560 24890
rect 34934 24508 35242 24528
rect 34934 24506 34940 24508
rect 34996 24506 35020 24508
rect 35076 24506 35100 24508
rect 35156 24506 35180 24508
rect 35236 24506 35242 24508
rect 34996 24454 34998 24506
rect 35178 24454 35180 24506
rect 34934 24452 34940 24454
rect 34996 24452 35020 24454
rect 35076 24452 35100 24454
rect 35156 24452 35180 24454
rect 35236 24452 35242 24454
rect 34934 24432 35242 24452
rect 34704 23724 34756 23730
rect 34704 23666 34756 23672
rect 34888 23724 34940 23730
rect 34888 23666 34940 23672
rect 34716 23050 34744 23666
rect 34900 23508 34928 23666
rect 34808 23480 34928 23508
rect 34704 23044 34756 23050
rect 34704 22986 34756 22992
rect 34808 23032 34836 23480
rect 34934 23420 35242 23440
rect 34934 23418 34940 23420
rect 34996 23418 35020 23420
rect 35076 23418 35100 23420
rect 35156 23418 35180 23420
rect 35236 23418 35242 23420
rect 34996 23366 34998 23418
rect 35178 23366 35180 23418
rect 34934 23364 34940 23366
rect 34996 23364 35020 23366
rect 35076 23364 35100 23366
rect 35156 23364 35180 23366
rect 35236 23364 35242 23366
rect 34934 23344 35242 23364
rect 34888 23044 34940 23050
rect 34808 23004 34888 23032
rect 34612 22976 34664 22982
rect 34612 22918 34664 22924
rect 34624 22642 34652 22918
rect 34716 22778 34744 22986
rect 34808 22778 34836 23004
rect 34888 22986 34940 22992
rect 34704 22772 34756 22778
rect 34704 22714 34756 22720
rect 34796 22772 34848 22778
rect 34796 22714 34848 22720
rect 34612 22636 34664 22642
rect 34612 22578 34664 22584
rect 34624 22506 34652 22578
rect 34520 22500 34572 22506
rect 34520 22442 34572 22448
rect 34612 22500 34664 22506
rect 34612 22442 34664 22448
rect 34532 22030 34560 22442
rect 34624 22094 34652 22442
rect 34934 22332 35242 22352
rect 34934 22330 34940 22332
rect 34996 22330 35020 22332
rect 35076 22330 35100 22332
rect 35156 22330 35180 22332
rect 35236 22330 35242 22332
rect 34996 22278 34998 22330
rect 35178 22278 35180 22330
rect 34934 22276 34940 22278
rect 34996 22276 35020 22278
rect 35076 22276 35100 22278
rect 35156 22276 35180 22278
rect 35236 22276 35242 22278
rect 34934 22256 35242 22276
rect 35360 22166 35388 26930
rect 37280 26308 37332 26314
rect 37280 26250 37332 26256
rect 37292 25838 37320 26250
rect 37280 25832 37332 25838
rect 37280 25774 37332 25780
rect 37188 25764 37240 25770
rect 37188 25706 37240 25712
rect 37200 25226 37228 25706
rect 37188 25220 37240 25226
rect 37188 25162 37240 25168
rect 36544 24812 36596 24818
rect 36544 24754 36596 24760
rect 35440 23792 35492 23798
rect 35440 23734 35492 23740
rect 35452 23322 35480 23734
rect 36556 23526 36584 24754
rect 36544 23520 36596 23526
rect 36544 23462 36596 23468
rect 36728 23520 36780 23526
rect 36728 23462 36780 23468
rect 35440 23316 35492 23322
rect 35440 23258 35492 23264
rect 35452 22778 35480 23258
rect 35624 22976 35676 22982
rect 35624 22918 35676 22924
rect 35440 22772 35492 22778
rect 35440 22714 35492 22720
rect 35636 22710 35664 22918
rect 35624 22704 35676 22710
rect 35624 22646 35676 22652
rect 35440 22636 35492 22642
rect 35440 22578 35492 22584
rect 35808 22636 35860 22642
rect 35808 22578 35860 22584
rect 35452 22234 35480 22578
rect 35820 22234 35848 22578
rect 36634 22536 36690 22545
rect 36634 22471 36636 22480
rect 36688 22471 36690 22480
rect 36636 22442 36688 22448
rect 36740 22438 36768 23462
rect 36728 22432 36780 22438
rect 36728 22374 36780 22380
rect 37200 22234 37228 25162
rect 37384 24614 37412 30790
rect 37464 30728 37516 30734
rect 37464 30670 37516 30676
rect 37476 30258 37504 30670
rect 37464 30252 37516 30258
rect 37464 30194 37516 30200
rect 37476 29850 37504 30194
rect 37568 30122 37596 31282
rect 37556 30116 37608 30122
rect 37556 30058 37608 30064
rect 37464 29844 37516 29850
rect 37464 29786 37516 29792
rect 37556 28620 37608 28626
rect 37556 28562 37608 28568
rect 37568 27334 37596 28562
rect 37660 27946 37688 37402
rect 38028 37194 38056 39200
rect 39120 37664 39172 37670
rect 39120 37606 39172 37612
rect 39132 37262 39160 37606
rect 39028 37256 39080 37262
rect 39028 37198 39080 37204
rect 39120 37256 39172 37262
rect 39120 37198 39172 37204
rect 39960 37210 39988 39200
rect 41892 37262 41920 39200
rect 46400 39114 46428 39200
rect 46492 39114 46520 39222
rect 46400 39086 46520 39114
rect 46756 37392 46808 37398
rect 46756 37334 46808 37340
rect 40132 37256 40184 37262
rect 38016 37188 38068 37194
rect 38016 37130 38068 37136
rect 38292 37120 38344 37126
rect 38292 37062 38344 37068
rect 38304 36786 38332 37062
rect 39040 36922 39068 37198
rect 39028 36916 39080 36922
rect 39028 36858 39080 36864
rect 38292 36780 38344 36786
rect 38292 36722 38344 36728
rect 38108 36236 38160 36242
rect 38108 36178 38160 36184
rect 37832 34604 37884 34610
rect 37832 34546 37884 34552
rect 37844 34066 37872 34546
rect 38120 34406 38148 36178
rect 38304 36174 38332 36722
rect 39040 36378 39068 36858
rect 39028 36372 39080 36378
rect 39028 36314 39080 36320
rect 38200 36168 38252 36174
rect 38200 36110 38252 36116
rect 38292 36168 38344 36174
rect 38292 36110 38344 36116
rect 38212 35834 38240 36110
rect 39132 36038 39160 37198
rect 39960 37182 40080 37210
rect 40132 37198 40184 37204
rect 41052 37256 41104 37262
rect 41052 37198 41104 37204
rect 41880 37256 41932 37262
rect 41880 37198 41932 37204
rect 42524 37256 42576 37262
rect 42524 37198 42576 37204
rect 40052 37126 40080 37182
rect 39212 37120 39264 37126
rect 39212 37062 39264 37068
rect 40040 37120 40092 37126
rect 40040 37062 40092 37068
rect 39224 36718 39252 37062
rect 40144 36922 40172 37198
rect 40132 36916 40184 36922
rect 40132 36858 40184 36864
rect 39212 36712 39264 36718
rect 40132 36712 40184 36718
rect 39264 36672 39436 36700
rect 39212 36654 39264 36660
rect 39408 36582 39436 36672
rect 40132 36654 40184 36660
rect 39304 36576 39356 36582
rect 39304 36518 39356 36524
rect 39396 36576 39448 36582
rect 39396 36518 39448 36524
rect 39316 36310 39344 36518
rect 39304 36304 39356 36310
rect 39304 36246 39356 36252
rect 40144 36038 40172 36654
rect 40316 36576 40368 36582
rect 40316 36518 40368 36524
rect 40328 36174 40356 36518
rect 40316 36168 40368 36174
rect 40316 36110 40368 36116
rect 39120 36032 39172 36038
rect 39120 35974 39172 35980
rect 40132 36032 40184 36038
rect 40132 35974 40184 35980
rect 40144 35834 40172 35974
rect 38200 35828 38252 35834
rect 38200 35770 38252 35776
rect 40132 35828 40184 35834
rect 40132 35770 40184 35776
rect 38212 34610 38240 35770
rect 41064 35494 41092 37198
rect 42536 36825 42564 37198
rect 43720 37188 43772 37194
rect 43720 37130 43772 37136
rect 46112 37188 46164 37194
rect 46112 37130 46164 37136
rect 42616 37120 42668 37126
rect 42616 37062 42668 37068
rect 42522 36816 42578 36825
rect 41880 36780 41932 36786
rect 42522 36751 42578 36760
rect 41880 36722 41932 36728
rect 41420 36576 41472 36582
rect 41420 36518 41472 36524
rect 41432 36378 41460 36518
rect 41420 36372 41472 36378
rect 41420 36314 41472 36320
rect 41420 36236 41472 36242
rect 41420 36178 41472 36184
rect 41052 35488 41104 35494
rect 41052 35430 41104 35436
rect 40316 35012 40368 35018
rect 40316 34954 40368 34960
rect 38936 34944 38988 34950
rect 38936 34886 38988 34892
rect 38948 34610 38976 34886
rect 40328 34678 40356 34954
rect 40316 34672 40368 34678
rect 40316 34614 40368 34620
rect 38200 34604 38252 34610
rect 38200 34546 38252 34552
rect 38936 34604 38988 34610
rect 38936 34546 38988 34552
rect 40040 34604 40092 34610
rect 40040 34546 40092 34552
rect 38292 34536 38344 34542
rect 38292 34478 38344 34484
rect 38108 34400 38160 34406
rect 38108 34342 38160 34348
rect 38304 34134 38332 34478
rect 38384 34468 38436 34474
rect 38384 34410 38436 34416
rect 38396 34202 38424 34410
rect 38384 34196 38436 34202
rect 38384 34138 38436 34144
rect 38292 34128 38344 34134
rect 38292 34070 38344 34076
rect 40052 34082 40080 34546
rect 40132 34536 40184 34542
rect 40132 34478 40184 34484
rect 40144 34202 40172 34478
rect 40316 34468 40368 34474
rect 40316 34410 40368 34416
rect 40132 34196 40184 34202
rect 40132 34138 40184 34144
rect 40224 34128 40276 34134
rect 40052 34076 40224 34082
rect 40052 34070 40276 34076
rect 37832 34060 37884 34066
rect 37832 34002 37884 34008
rect 40052 34054 40264 34070
rect 39948 33992 40000 33998
rect 39948 33934 40000 33940
rect 39960 33454 39988 33934
rect 39948 33448 40000 33454
rect 39948 33390 40000 33396
rect 38660 33040 38712 33046
rect 38660 32982 38712 32988
rect 38292 32836 38344 32842
rect 38292 32778 38344 32784
rect 38304 32570 38332 32778
rect 38292 32564 38344 32570
rect 38292 32506 38344 32512
rect 38200 32428 38252 32434
rect 38200 32370 38252 32376
rect 38016 32292 38068 32298
rect 38016 32234 38068 32240
rect 38028 31822 38056 32234
rect 38212 31822 38240 32370
rect 38672 31890 38700 32982
rect 39028 32768 39080 32774
rect 39028 32710 39080 32716
rect 39040 32434 39068 32710
rect 40052 32570 40080 34054
rect 40328 33998 40356 34410
rect 40316 33992 40368 33998
rect 40316 33934 40368 33940
rect 40040 32564 40092 32570
rect 40040 32506 40092 32512
rect 39028 32428 39080 32434
rect 39028 32370 39080 32376
rect 39212 32428 39264 32434
rect 39212 32370 39264 32376
rect 39040 31958 39068 32370
rect 39028 31952 39080 31958
rect 39028 31894 39080 31900
rect 38660 31884 38712 31890
rect 38660 31826 38712 31832
rect 39224 31822 39252 32370
rect 41064 31958 41092 35430
rect 41328 32428 41380 32434
rect 41328 32370 41380 32376
rect 41236 32360 41288 32366
rect 41236 32302 41288 32308
rect 41052 31952 41104 31958
rect 41052 31894 41104 31900
rect 41248 31890 41276 32302
rect 41340 31890 41368 32370
rect 41236 31884 41288 31890
rect 41236 31826 41288 31832
rect 41328 31884 41380 31890
rect 41328 31826 41380 31832
rect 38016 31816 38068 31822
rect 38016 31758 38068 31764
rect 38200 31816 38252 31822
rect 38200 31758 38252 31764
rect 39212 31816 39264 31822
rect 39212 31758 39264 31764
rect 38212 31482 38240 31758
rect 38200 31476 38252 31482
rect 38200 31418 38252 31424
rect 40500 31340 40552 31346
rect 40500 31282 40552 31288
rect 40408 30388 40460 30394
rect 40408 30330 40460 30336
rect 39672 30184 39724 30190
rect 39856 30184 39908 30190
rect 39724 30132 39856 30138
rect 39672 30126 39908 30132
rect 39684 30110 39896 30126
rect 39684 28694 39712 30110
rect 40420 29646 40448 30330
rect 40512 30326 40540 31282
rect 41340 31278 41368 31826
rect 40684 31272 40736 31278
rect 40684 31214 40736 31220
rect 41328 31272 41380 31278
rect 41328 31214 41380 31220
rect 40696 30394 40724 31214
rect 40684 30388 40736 30394
rect 40684 30330 40736 30336
rect 40500 30320 40552 30326
rect 40500 30262 40552 30268
rect 40408 29640 40460 29646
rect 40408 29582 40460 29588
rect 40512 29510 40540 30262
rect 40592 30048 40644 30054
rect 40592 29990 40644 29996
rect 40604 29646 40632 29990
rect 40592 29640 40644 29646
rect 40592 29582 40644 29588
rect 40500 29504 40552 29510
rect 40500 29446 40552 29452
rect 39672 28688 39724 28694
rect 39672 28630 39724 28636
rect 39120 28620 39172 28626
rect 39120 28562 39172 28568
rect 37740 28552 37792 28558
rect 37740 28494 37792 28500
rect 37752 28218 37780 28494
rect 37740 28212 37792 28218
rect 37740 28154 37792 28160
rect 39132 28082 39160 28562
rect 39304 28552 39356 28558
rect 39304 28494 39356 28500
rect 39316 28082 39344 28494
rect 39120 28076 39172 28082
rect 39120 28018 39172 28024
rect 39304 28076 39356 28082
rect 39304 28018 39356 28024
rect 41052 28076 41104 28082
rect 41052 28018 41104 28024
rect 41144 28076 41196 28082
rect 41144 28018 41196 28024
rect 41328 28076 41380 28082
rect 41328 28018 41380 28024
rect 37648 27940 37700 27946
rect 37648 27882 37700 27888
rect 39316 27606 39344 28018
rect 41064 27674 41092 28018
rect 41052 27668 41104 27674
rect 41052 27610 41104 27616
rect 39304 27600 39356 27606
rect 39304 27542 39356 27548
rect 38108 27532 38160 27538
rect 38108 27474 38160 27480
rect 37556 27328 37608 27334
rect 37556 27270 37608 27276
rect 38120 26994 38148 27474
rect 38200 27464 38252 27470
rect 38200 27406 38252 27412
rect 40868 27464 40920 27470
rect 40868 27406 40920 27412
rect 38212 27062 38240 27406
rect 40880 27130 40908 27406
rect 40868 27124 40920 27130
rect 40868 27066 40920 27072
rect 38200 27056 38252 27062
rect 38200 26998 38252 27004
rect 39948 27056 40000 27062
rect 39948 26998 40000 27004
rect 37648 26988 37700 26994
rect 37648 26930 37700 26936
rect 38108 26988 38160 26994
rect 38108 26930 38160 26936
rect 37464 26376 37516 26382
rect 37464 26318 37516 26324
rect 37476 25906 37504 26318
rect 37464 25900 37516 25906
rect 37464 25842 37516 25848
rect 37476 25430 37504 25842
rect 37464 25424 37516 25430
rect 37464 25366 37516 25372
rect 37372 24608 37424 24614
rect 37372 24550 37424 24556
rect 37384 24070 37412 24550
rect 37660 24342 37688 26930
rect 38212 26586 38240 26998
rect 38200 26580 38252 26586
rect 38200 26522 38252 26528
rect 38108 26376 38160 26382
rect 38108 26318 38160 26324
rect 38752 26376 38804 26382
rect 38752 26318 38804 26324
rect 38016 25832 38068 25838
rect 38016 25774 38068 25780
rect 38028 25430 38056 25774
rect 38120 25430 38148 26318
rect 38764 26042 38792 26318
rect 39960 26246 39988 26998
rect 40224 26988 40276 26994
rect 40224 26930 40276 26936
rect 40500 26988 40552 26994
rect 40500 26930 40552 26936
rect 40236 26382 40264 26930
rect 40512 26450 40540 26930
rect 41064 26858 41092 27610
rect 41156 27402 41184 28018
rect 41236 28008 41288 28014
rect 41236 27950 41288 27956
rect 41248 27538 41276 27950
rect 41236 27532 41288 27538
rect 41236 27474 41288 27480
rect 41340 27470 41368 28018
rect 41328 27464 41380 27470
rect 41328 27406 41380 27412
rect 41144 27396 41196 27402
rect 41144 27338 41196 27344
rect 41156 27282 41184 27338
rect 41156 27254 41368 27282
rect 41340 27130 41368 27254
rect 41328 27124 41380 27130
rect 41328 27066 41380 27072
rect 41052 26852 41104 26858
rect 41052 26794 41104 26800
rect 41144 26784 41196 26790
rect 41144 26726 41196 26732
rect 40500 26444 40552 26450
rect 40500 26386 40552 26392
rect 41156 26382 41184 26726
rect 40224 26376 40276 26382
rect 40224 26318 40276 26324
rect 41144 26376 41196 26382
rect 41144 26318 41196 26324
rect 39948 26240 40000 26246
rect 39948 26182 40000 26188
rect 38752 26036 38804 26042
rect 38752 25978 38804 25984
rect 38016 25424 38068 25430
rect 38016 25366 38068 25372
rect 38108 25424 38160 25430
rect 38108 25366 38160 25372
rect 39120 24812 39172 24818
rect 39120 24754 39172 24760
rect 38568 24744 38620 24750
rect 38568 24686 38620 24692
rect 37740 24608 37792 24614
rect 37740 24550 37792 24556
rect 37648 24336 37700 24342
rect 37648 24278 37700 24284
rect 37752 24138 37780 24550
rect 38580 24410 38608 24686
rect 39132 24410 39160 24754
rect 39960 24614 39988 26182
rect 40132 25696 40184 25702
rect 40132 25638 40184 25644
rect 40144 25294 40172 25638
rect 40132 25288 40184 25294
rect 40132 25230 40184 25236
rect 40144 24818 40172 25230
rect 40132 24812 40184 24818
rect 40132 24754 40184 24760
rect 39948 24608 40000 24614
rect 39948 24550 40000 24556
rect 40236 24410 40264 26318
rect 40960 25288 41012 25294
rect 40960 25230 41012 25236
rect 40316 25220 40368 25226
rect 40316 25162 40368 25168
rect 40328 24818 40356 25162
rect 40972 24954 41000 25230
rect 40960 24948 41012 24954
rect 40960 24890 41012 24896
rect 40316 24812 40368 24818
rect 40316 24754 40368 24760
rect 40972 24614 41000 24890
rect 40960 24608 41012 24614
rect 40960 24550 41012 24556
rect 38568 24404 38620 24410
rect 38568 24346 38620 24352
rect 39120 24404 39172 24410
rect 39120 24346 39172 24352
rect 40224 24404 40276 24410
rect 40224 24346 40276 24352
rect 40592 24268 40644 24274
rect 40592 24210 40644 24216
rect 38108 24200 38160 24206
rect 38108 24142 38160 24148
rect 37740 24132 37792 24138
rect 37740 24074 37792 24080
rect 37372 24064 37424 24070
rect 37372 24006 37424 24012
rect 37752 23730 37780 24074
rect 37280 23724 37332 23730
rect 37280 23666 37332 23672
rect 37464 23724 37516 23730
rect 37464 23666 37516 23672
rect 37740 23724 37792 23730
rect 37740 23666 37792 23672
rect 35440 22228 35492 22234
rect 35440 22170 35492 22176
rect 35808 22228 35860 22234
rect 35808 22170 35860 22176
rect 37188 22228 37240 22234
rect 37188 22170 37240 22176
rect 34796 22160 34848 22166
rect 34796 22102 34848 22108
rect 35348 22160 35400 22166
rect 35348 22102 35400 22108
rect 34624 22066 34744 22094
rect 34520 22024 34572 22030
rect 34520 21966 34572 21972
rect 34532 21690 34560 21966
rect 34716 21894 34744 22066
rect 34704 21888 34756 21894
rect 34704 21830 34756 21836
rect 34520 21684 34572 21690
rect 34520 21626 34572 21632
rect 34612 21684 34664 21690
rect 34612 21626 34664 21632
rect 34624 21146 34652 21626
rect 34612 21140 34664 21146
rect 34612 21082 34664 21088
rect 34716 21026 34744 21830
rect 34808 21554 34836 22102
rect 36820 22092 36872 22098
rect 36820 22034 36872 22040
rect 35348 21616 35400 21622
rect 35348 21558 35400 21564
rect 34796 21548 34848 21554
rect 34796 21490 34848 21496
rect 34934 21244 35242 21264
rect 34934 21242 34940 21244
rect 34996 21242 35020 21244
rect 35076 21242 35100 21244
rect 35156 21242 35180 21244
rect 35236 21242 35242 21244
rect 34996 21190 34998 21242
rect 35178 21190 35180 21242
rect 34934 21188 34940 21190
rect 34996 21188 35020 21190
rect 35076 21188 35100 21190
rect 35156 21188 35180 21190
rect 35236 21188 35242 21190
rect 34934 21168 35242 21188
rect 35360 21146 35388 21558
rect 36832 21418 36860 22034
rect 37292 22030 37320 23666
rect 37476 23526 37504 23666
rect 37464 23520 37516 23526
rect 37464 23462 37516 23468
rect 37752 23254 37780 23666
rect 37740 23248 37792 23254
rect 37740 23190 37792 23196
rect 38120 22778 38148 24142
rect 38384 24064 38436 24070
rect 38384 24006 38436 24012
rect 38108 22772 38160 22778
rect 38108 22714 38160 22720
rect 38200 22092 38252 22098
rect 38200 22034 38252 22040
rect 37280 22024 37332 22030
rect 37280 21966 37332 21972
rect 37292 21486 37320 21966
rect 38212 21894 38240 22034
rect 38200 21888 38252 21894
rect 38200 21830 38252 21836
rect 37280 21480 37332 21486
rect 37280 21422 37332 21428
rect 36820 21412 36872 21418
rect 36820 21354 36872 21360
rect 37004 21344 37056 21350
rect 37004 21286 37056 21292
rect 35348 21140 35400 21146
rect 35348 21082 35400 21088
rect 34624 20998 34744 21026
rect 34520 20868 34572 20874
rect 34520 20810 34572 20816
rect 34532 20466 34560 20810
rect 34624 20505 34652 20998
rect 37016 20942 37044 21286
rect 34796 20936 34848 20942
rect 34716 20884 34796 20890
rect 34716 20878 34848 20884
rect 37004 20936 37056 20942
rect 38212 20913 38240 21830
rect 37004 20878 37056 20884
rect 38198 20904 38254 20913
rect 34716 20862 34836 20878
rect 34888 20868 34940 20874
rect 34610 20496 34666 20505
rect 34520 20460 34572 20466
rect 34716 20466 34744 20862
rect 34888 20810 34940 20816
rect 34900 20602 34928 20810
rect 34888 20596 34940 20602
rect 34888 20538 34940 20544
rect 34610 20431 34666 20440
rect 34704 20460 34756 20466
rect 34520 20402 34572 20408
rect 34704 20402 34756 20408
rect 34532 20058 34560 20402
rect 34520 20052 34572 20058
rect 34520 19994 34572 20000
rect 34336 19372 34388 19378
rect 34336 19314 34388 19320
rect 34716 18970 34744 20402
rect 34796 20392 34848 20398
rect 34796 20334 34848 20340
rect 34808 19854 34836 20334
rect 34934 20156 35242 20176
rect 34934 20154 34940 20156
rect 34996 20154 35020 20156
rect 35076 20154 35100 20156
rect 35156 20154 35180 20156
rect 35236 20154 35242 20156
rect 34996 20102 34998 20154
rect 35178 20102 35180 20154
rect 34934 20100 34940 20102
rect 34996 20100 35020 20102
rect 35076 20100 35100 20102
rect 35156 20100 35180 20102
rect 35236 20100 35242 20102
rect 34934 20080 35242 20100
rect 34796 19848 34848 19854
rect 34796 19790 34848 19796
rect 35992 19848 36044 19854
rect 35992 19790 36044 19796
rect 36176 19848 36228 19854
rect 36176 19790 36228 19796
rect 34808 19514 34836 19790
rect 34796 19508 34848 19514
rect 34796 19450 34848 19456
rect 36004 19446 36032 19790
rect 35992 19440 36044 19446
rect 35992 19382 36044 19388
rect 36188 19378 36216 19790
rect 37016 19378 37044 20878
rect 38198 20839 38254 20848
rect 37372 20800 37424 20806
rect 37372 20742 37424 20748
rect 37384 20466 37412 20742
rect 37372 20460 37424 20466
rect 37372 20402 37424 20408
rect 38292 20460 38344 20466
rect 38292 20402 38344 20408
rect 38304 19922 38332 20402
rect 38292 19916 38344 19922
rect 38292 19858 38344 19864
rect 36176 19372 36228 19378
rect 36176 19314 36228 19320
rect 37004 19372 37056 19378
rect 37004 19314 37056 19320
rect 37188 19372 37240 19378
rect 37188 19314 37240 19320
rect 34934 19068 35242 19088
rect 34934 19066 34940 19068
rect 34996 19066 35020 19068
rect 35076 19066 35100 19068
rect 35156 19066 35180 19068
rect 35236 19066 35242 19068
rect 34996 19014 34998 19066
rect 35178 19014 35180 19066
rect 34934 19012 34940 19014
rect 34996 19012 35020 19014
rect 35076 19012 35100 19014
rect 35156 19012 35180 19014
rect 35236 19012 35242 19014
rect 34934 18992 35242 19012
rect 34704 18964 34756 18970
rect 34704 18906 34756 18912
rect 34520 18896 34572 18902
rect 34520 18838 34572 18844
rect 35992 18896 36044 18902
rect 35992 18838 36044 18844
rect 33600 18760 33652 18766
rect 33600 18702 33652 18708
rect 33968 18760 34020 18766
rect 33968 18702 34020 18708
rect 33612 18154 33640 18702
rect 33600 18148 33652 18154
rect 33600 18090 33652 18096
rect 33980 18086 34008 18702
rect 34336 18692 34388 18698
rect 34336 18634 34388 18640
rect 34348 18426 34376 18634
rect 34532 18630 34560 18838
rect 35716 18760 35768 18766
rect 35716 18702 35768 18708
rect 34520 18624 34572 18630
rect 34520 18566 34572 18572
rect 34532 18426 34560 18566
rect 35728 18426 35756 18702
rect 35900 18624 35952 18630
rect 35900 18566 35952 18572
rect 34336 18420 34388 18426
rect 34336 18362 34388 18368
rect 34520 18420 34572 18426
rect 34520 18362 34572 18368
rect 35716 18420 35768 18426
rect 35716 18362 35768 18368
rect 34348 18290 34376 18362
rect 34336 18284 34388 18290
rect 34336 18226 34388 18232
rect 34428 18284 34480 18290
rect 34428 18226 34480 18232
rect 33968 18080 34020 18086
rect 33968 18022 34020 18028
rect 33416 17876 33468 17882
rect 33416 17818 33468 17824
rect 33416 17672 33468 17678
rect 33336 17632 33416 17660
rect 33416 17614 33468 17620
rect 33324 15360 33376 15366
rect 33324 15302 33376 15308
rect 33336 14958 33364 15302
rect 33324 14952 33376 14958
rect 33324 14894 33376 14900
rect 33336 14278 33364 14894
rect 33428 14482 33456 17614
rect 33784 17536 33836 17542
rect 33836 17484 33916 17490
rect 33784 17478 33916 17484
rect 33796 17462 33916 17478
rect 33520 17202 33732 17218
rect 33508 17196 33744 17202
rect 33560 17190 33692 17196
rect 33508 17138 33560 17144
rect 33692 17138 33744 17144
rect 33784 16992 33836 16998
rect 33784 16934 33836 16940
rect 33796 16658 33824 16934
rect 33784 16652 33836 16658
rect 33784 16594 33836 16600
rect 33508 15360 33560 15366
rect 33508 15302 33560 15308
rect 33520 15026 33548 15302
rect 33508 15020 33560 15026
rect 33508 14962 33560 14968
rect 33888 14958 33916 17462
rect 33980 16590 34008 18022
rect 34440 17542 34468 18226
rect 35728 18222 35756 18362
rect 35716 18216 35768 18222
rect 35716 18158 35768 18164
rect 35808 18148 35860 18154
rect 35808 18090 35860 18096
rect 34934 17980 35242 18000
rect 34934 17978 34940 17980
rect 34996 17978 35020 17980
rect 35076 17978 35100 17980
rect 35156 17978 35180 17980
rect 35236 17978 35242 17980
rect 34996 17926 34998 17978
rect 35178 17926 35180 17978
rect 34934 17924 34940 17926
rect 34996 17924 35020 17926
rect 35076 17924 35100 17926
rect 35156 17924 35180 17926
rect 35236 17924 35242 17926
rect 34934 17904 35242 17924
rect 34428 17536 34480 17542
rect 34428 17478 34480 17484
rect 34428 17196 34480 17202
rect 34428 17138 34480 17144
rect 33968 16584 34020 16590
rect 33968 16526 34020 16532
rect 34440 16250 34468 17138
rect 35348 17060 35400 17066
rect 35348 17002 35400 17008
rect 34934 16892 35242 16912
rect 34934 16890 34940 16892
rect 34996 16890 35020 16892
rect 35076 16890 35100 16892
rect 35156 16890 35180 16892
rect 35236 16890 35242 16892
rect 34996 16838 34998 16890
rect 35178 16838 35180 16890
rect 34934 16836 34940 16838
rect 34996 16836 35020 16838
rect 35076 16836 35100 16838
rect 35156 16836 35180 16838
rect 35236 16836 35242 16838
rect 34934 16816 35242 16836
rect 35256 16652 35308 16658
rect 35360 16640 35388 17002
rect 35308 16612 35388 16640
rect 35256 16594 35308 16600
rect 34520 16448 34572 16454
rect 34520 16390 34572 16396
rect 34428 16244 34480 16250
rect 34428 16186 34480 16192
rect 34532 16114 34560 16390
rect 35268 16182 35296 16594
rect 35256 16176 35308 16182
rect 35256 16118 35308 16124
rect 35820 16114 35848 18090
rect 35912 17610 35940 18566
rect 36004 18290 36032 18838
rect 35992 18284 36044 18290
rect 35992 18226 36044 18232
rect 36084 18284 36136 18290
rect 36084 18226 36136 18232
rect 36096 17814 36124 18226
rect 36084 17808 36136 17814
rect 36084 17750 36136 17756
rect 35900 17604 35952 17610
rect 35900 17546 35952 17552
rect 36188 16980 36216 19314
rect 36360 18760 36412 18766
rect 36360 18702 36412 18708
rect 36268 18692 36320 18698
rect 36268 18634 36320 18640
rect 36280 17882 36308 18634
rect 36268 17876 36320 17882
rect 36268 17818 36320 17824
rect 36096 16952 36216 16980
rect 36096 16590 36124 16952
rect 36084 16584 36136 16590
rect 36084 16526 36136 16532
rect 34520 16108 34572 16114
rect 34520 16050 34572 16056
rect 35808 16108 35860 16114
rect 35808 16050 35860 16056
rect 34060 16040 34112 16046
rect 34060 15982 34112 15988
rect 34336 16040 34388 16046
rect 34336 15982 34388 15988
rect 33876 14952 33928 14958
rect 33876 14894 33928 14900
rect 33784 14884 33836 14890
rect 33784 14826 33836 14832
rect 33416 14476 33468 14482
rect 33416 14418 33468 14424
rect 33796 14278 33824 14826
rect 33888 14550 33916 14894
rect 33876 14544 33928 14550
rect 33876 14486 33928 14492
rect 33324 14272 33376 14278
rect 33324 14214 33376 14220
rect 33784 14272 33836 14278
rect 33784 14214 33836 14220
rect 33232 14000 33284 14006
rect 33232 13942 33284 13948
rect 32496 13932 32548 13938
rect 32496 13874 32548 13880
rect 32588 13932 32640 13938
rect 32588 13874 32640 13880
rect 32128 13252 32180 13258
rect 32128 13194 32180 13200
rect 32312 13252 32364 13258
rect 32312 13194 32364 13200
rect 32324 12850 32352 13194
rect 32508 13190 32536 13874
rect 32600 13326 32628 13874
rect 33244 13734 33272 13942
rect 33796 13938 33824 14214
rect 33784 13932 33836 13938
rect 33784 13874 33836 13880
rect 34072 13734 34100 15982
rect 34348 15026 34376 15982
rect 34934 15804 35242 15824
rect 34934 15802 34940 15804
rect 34996 15802 35020 15804
rect 35076 15802 35100 15804
rect 35156 15802 35180 15804
rect 35236 15802 35242 15804
rect 34996 15750 34998 15802
rect 35178 15750 35180 15802
rect 34934 15748 34940 15750
rect 34996 15748 35020 15750
rect 35076 15748 35100 15750
rect 35156 15748 35180 15750
rect 35236 15748 35242 15750
rect 34934 15728 35242 15748
rect 34336 15020 34388 15026
rect 34336 14962 34388 14968
rect 34520 14816 34572 14822
rect 34520 14758 34572 14764
rect 34612 14816 34664 14822
rect 34612 14758 34664 14764
rect 34532 14346 34560 14758
rect 34624 14482 34652 14758
rect 34934 14716 35242 14736
rect 34934 14714 34940 14716
rect 34996 14714 35020 14716
rect 35076 14714 35100 14716
rect 35156 14714 35180 14716
rect 35236 14714 35242 14716
rect 34996 14662 34998 14714
rect 35178 14662 35180 14714
rect 34934 14660 34940 14662
rect 34996 14660 35020 14662
rect 35076 14660 35100 14662
rect 35156 14660 35180 14662
rect 35236 14660 35242 14662
rect 34934 14640 35242 14660
rect 34612 14476 34664 14482
rect 34612 14418 34664 14424
rect 34980 14408 35032 14414
rect 34980 14350 35032 14356
rect 34520 14340 34572 14346
rect 34520 14282 34572 14288
rect 34532 13870 34560 14282
rect 34992 13938 35020 14350
rect 35820 13938 35848 16050
rect 34980 13932 35032 13938
rect 34980 13874 35032 13880
rect 35808 13932 35860 13938
rect 35808 13874 35860 13880
rect 34520 13864 34572 13870
rect 34520 13806 34572 13812
rect 32680 13728 32732 13734
rect 32680 13670 32732 13676
rect 33232 13728 33284 13734
rect 33232 13670 33284 13676
rect 34060 13728 34112 13734
rect 34060 13670 34112 13676
rect 32588 13320 32640 13326
rect 32588 13262 32640 13268
rect 32496 13184 32548 13190
rect 32496 13126 32548 13132
rect 32036 12844 32088 12850
rect 32036 12786 32088 12792
rect 32312 12844 32364 12850
rect 32312 12786 32364 12792
rect 32692 12782 32720 13670
rect 34934 13628 35242 13648
rect 34934 13626 34940 13628
rect 34996 13626 35020 13628
rect 35076 13626 35100 13628
rect 35156 13626 35180 13628
rect 35236 13626 35242 13628
rect 34996 13574 34998 13626
rect 35178 13574 35180 13626
rect 34934 13572 34940 13574
rect 34996 13572 35020 13574
rect 35076 13572 35100 13574
rect 35156 13572 35180 13574
rect 35236 13572 35242 13574
rect 34934 13552 35242 13572
rect 34796 13184 34848 13190
rect 34796 13126 34848 13132
rect 32496 12776 32548 12782
rect 32496 12718 32548 12724
rect 32680 12776 32732 12782
rect 32680 12718 32732 12724
rect 33140 12776 33192 12782
rect 33140 12718 33192 12724
rect 32508 12442 32536 12718
rect 32496 12436 32548 12442
rect 32496 12378 32548 12384
rect 31760 12232 31812 12238
rect 31760 12174 31812 12180
rect 31944 12096 31996 12102
rect 31944 12038 31996 12044
rect 31956 11218 31984 12038
rect 32508 11898 32536 12378
rect 32496 11892 32548 11898
rect 32496 11834 32548 11840
rect 31944 11212 31996 11218
rect 31944 11154 31996 11160
rect 32680 11076 32732 11082
rect 32680 11018 32732 11024
rect 31576 10260 31628 10266
rect 31576 10202 31628 10208
rect 32692 10062 32720 11018
rect 32680 10056 32732 10062
rect 32680 9998 32732 10004
rect 33152 9110 33180 12718
rect 34808 12442 34836 13126
rect 34934 12540 35242 12560
rect 34934 12538 34940 12540
rect 34996 12538 35020 12540
rect 35076 12538 35100 12540
rect 35156 12538 35180 12540
rect 35236 12538 35242 12540
rect 34996 12486 34998 12538
rect 35178 12486 35180 12538
rect 34934 12484 34940 12486
rect 34996 12484 35020 12486
rect 35076 12484 35100 12486
rect 35156 12484 35180 12486
rect 35236 12484 35242 12486
rect 34934 12464 35242 12484
rect 34796 12436 34848 12442
rect 34796 12378 34848 12384
rect 34520 12300 34572 12306
rect 34520 12242 34572 12248
rect 33784 12096 33836 12102
rect 33784 12038 33836 12044
rect 33692 11892 33744 11898
rect 33692 11834 33744 11840
rect 33600 11824 33652 11830
rect 33600 11766 33652 11772
rect 33612 11082 33640 11766
rect 33704 11150 33732 11834
rect 33796 11558 33824 12038
rect 34532 11762 34560 12242
rect 34704 12164 34756 12170
rect 34704 12106 34756 12112
rect 34716 11762 34744 12106
rect 34808 11898 34836 12378
rect 35348 12096 35400 12102
rect 35348 12038 35400 12044
rect 34796 11892 34848 11898
rect 34796 11834 34848 11840
rect 34520 11756 34572 11762
rect 34520 11698 34572 11704
rect 34704 11756 34756 11762
rect 34704 11698 34756 11704
rect 33784 11552 33836 11558
rect 33784 11494 33836 11500
rect 34704 11552 34756 11558
rect 34704 11494 34756 11500
rect 33796 11150 33824 11494
rect 33692 11144 33744 11150
rect 33692 11086 33744 11092
rect 33784 11144 33836 11150
rect 33784 11086 33836 11092
rect 34716 11082 34744 11494
rect 34934 11452 35242 11472
rect 34934 11450 34940 11452
rect 34996 11450 35020 11452
rect 35076 11450 35100 11452
rect 35156 11450 35180 11452
rect 35236 11450 35242 11452
rect 34996 11398 34998 11450
rect 35178 11398 35180 11450
rect 34934 11396 34940 11398
rect 34996 11396 35020 11398
rect 35076 11396 35100 11398
rect 35156 11396 35180 11398
rect 35236 11396 35242 11398
rect 34934 11376 35242 11396
rect 35360 11218 35388 12038
rect 36096 11762 36124 16526
rect 36176 13728 36228 13734
rect 36176 13670 36228 13676
rect 36188 13326 36216 13670
rect 36176 13320 36228 13326
rect 36176 13262 36228 13268
rect 36084 11756 36136 11762
rect 36084 11698 36136 11704
rect 35440 11552 35492 11558
rect 35440 11494 35492 11500
rect 35348 11212 35400 11218
rect 35348 11154 35400 11160
rect 34796 11144 34848 11150
rect 34796 11086 34848 11092
rect 33600 11076 33652 11082
rect 33600 11018 33652 11024
rect 34704 11076 34756 11082
rect 34704 11018 34756 11024
rect 33612 10674 33640 11018
rect 34716 10742 34744 11018
rect 34704 10736 34756 10742
rect 34704 10678 34756 10684
rect 33600 10668 33652 10674
rect 33600 10610 33652 10616
rect 34808 10606 34836 11086
rect 35360 10724 35388 11154
rect 35452 11150 35480 11494
rect 35808 11280 35860 11286
rect 35808 11222 35860 11228
rect 35440 11144 35492 11150
rect 35440 11086 35492 11092
rect 35268 10696 35388 10724
rect 34796 10600 34848 10606
rect 34796 10542 34848 10548
rect 35268 10538 35296 10696
rect 35452 10674 35480 11086
rect 35532 11008 35584 11014
rect 35532 10950 35584 10956
rect 35440 10668 35492 10674
rect 35440 10610 35492 10616
rect 35256 10532 35308 10538
rect 35256 10474 35308 10480
rect 35544 10470 35572 10950
rect 35532 10464 35584 10470
rect 35532 10406 35584 10412
rect 34934 10364 35242 10384
rect 34934 10362 34940 10364
rect 34996 10362 35020 10364
rect 35076 10362 35100 10364
rect 35156 10362 35180 10364
rect 35236 10362 35242 10364
rect 34996 10310 34998 10362
rect 35178 10310 35180 10362
rect 34934 10308 34940 10310
rect 34996 10308 35020 10310
rect 35076 10308 35100 10310
rect 35156 10308 35180 10310
rect 35236 10308 35242 10310
rect 34934 10288 35242 10308
rect 33416 10056 33468 10062
rect 33416 9998 33468 10004
rect 33232 9172 33284 9178
rect 33232 9114 33284 9120
rect 33140 9104 33192 9110
rect 33140 9046 33192 9052
rect 33152 8974 33180 9046
rect 32128 8968 32180 8974
rect 32128 8910 32180 8916
rect 33140 8968 33192 8974
rect 33140 8910 33192 8916
rect 31576 8356 31628 8362
rect 31576 8298 31628 8304
rect 31588 7954 31616 8298
rect 31668 8288 31720 8294
rect 31668 8230 31720 8236
rect 31576 7948 31628 7954
rect 31576 7890 31628 7896
rect 31680 7546 31708 8230
rect 32140 7954 32168 8910
rect 33152 7954 33180 8910
rect 32128 7948 32180 7954
rect 32128 7890 32180 7896
rect 33140 7948 33192 7954
rect 33140 7890 33192 7896
rect 31944 7744 31996 7750
rect 31944 7686 31996 7692
rect 31484 7540 31536 7546
rect 31484 7482 31536 7488
rect 31668 7540 31720 7546
rect 31668 7482 31720 7488
rect 31496 7410 31524 7482
rect 31956 7478 31984 7686
rect 31944 7472 31996 7478
rect 31944 7414 31996 7420
rect 31484 7404 31536 7410
rect 31484 7346 31536 7352
rect 32312 7404 32364 7410
rect 32312 7346 32364 7352
rect 30564 7336 30616 7342
rect 30564 7278 30616 7284
rect 31024 7268 31076 7274
rect 31024 7210 31076 7216
rect 31036 6798 31064 7210
rect 32324 7206 32352 7346
rect 32312 7200 32364 7206
rect 32312 7142 32364 7148
rect 32324 6866 32352 7142
rect 33152 7002 33180 7890
rect 33244 7342 33272 9114
rect 33428 7886 33456 9998
rect 35360 9926 35388 9957
rect 33692 9920 33744 9926
rect 35348 9920 35400 9926
rect 33692 9862 33744 9868
rect 35346 9888 35348 9897
rect 35400 9888 35402 9897
rect 33704 8974 33732 9862
rect 35346 9823 35402 9832
rect 35360 9722 35388 9823
rect 35348 9716 35400 9722
rect 35348 9658 35400 9664
rect 34934 9276 35242 9296
rect 34934 9274 34940 9276
rect 34996 9274 35020 9276
rect 35076 9274 35100 9276
rect 35156 9274 35180 9276
rect 35236 9274 35242 9276
rect 34996 9222 34998 9274
rect 35178 9222 35180 9274
rect 34934 9220 34940 9222
rect 34996 9220 35020 9222
rect 35076 9220 35100 9222
rect 35156 9220 35180 9222
rect 35236 9220 35242 9222
rect 34934 9200 35242 9220
rect 34612 9036 34664 9042
rect 34612 8978 34664 8984
rect 33692 8968 33744 8974
rect 33692 8910 33744 8916
rect 34428 8968 34480 8974
rect 34428 8910 34480 8916
rect 34440 8498 34468 8910
rect 34624 8498 34652 8978
rect 34428 8492 34480 8498
rect 34428 8434 34480 8440
rect 34612 8492 34664 8498
rect 34612 8434 34664 8440
rect 34934 8188 35242 8208
rect 34934 8186 34940 8188
rect 34996 8186 35020 8188
rect 35076 8186 35100 8188
rect 35156 8186 35180 8188
rect 35236 8186 35242 8188
rect 34996 8134 34998 8186
rect 35178 8134 35180 8186
rect 34934 8132 34940 8134
rect 34996 8132 35020 8134
rect 35076 8132 35100 8134
rect 35156 8132 35180 8134
rect 35236 8132 35242 8134
rect 34934 8112 35242 8132
rect 35624 8084 35676 8090
rect 35624 8026 35676 8032
rect 33416 7880 33468 7886
rect 33416 7822 33468 7828
rect 33968 7744 34020 7750
rect 33968 7686 34020 7692
rect 34888 7744 34940 7750
rect 34888 7686 34940 7692
rect 33980 7410 34008 7686
rect 34900 7410 34928 7686
rect 35532 7540 35584 7546
rect 35532 7482 35584 7488
rect 33968 7404 34020 7410
rect 33968 7346 34020 7352
rect 34888 7404 34940 7410
rect 34888 7346 34940 7352
rect 33232 7336 33284 7342
rect 33232 7278 33284 7284
rect 34704 7268 34756 7274
rect 34704 7210 34756 7216
rect 33140 6996 33192 7002
rect 33140 6938 33192 6944
rect 32312 6860 32364 6866
rect 32312 6802 32364 6808
rect 34716 6798 34744 7210
rect 34934 7100 35242 7120
rect 34934 7098 34940 7100
rect 34996 7098 35020 7100
rect 35076 7098 35100 7100
rect 35156 7098 35180 7100
rect 35236 7098 35242 7100
rect 34996 7046 34998 7098
rect 35178 7046 35180 7098
rect 34934 7044 34940 7046
rect 34996 7044 35020 7046
rect 35076 7044 35100 7046
rect 35156 7044 35180 7046
rect 35236 7044 35242 7046
rect 34934 7024 35242 7044
rect 35544 6798 35572 7482
rect 35636 7342 35664 8026
rect 35716 7880 35768 7886
rect 35716 7822 35768 7828
rect 35728 7410 35756 7822
rect 35820 7750 35848 11222
rect 36096 11150 36124 11698
rect 36188 11286 36216 13262
rect 36280 11830 36308 17818
rect 36372 16998 36400 18702
rect 36544 17604 36596 17610
rect 36544 17546 36596 17552
rect 36556 17270 36584 17546
rect 36452 17264 36504 17270
rect 36452 17206 36504 17212
rect 36544 17264 36596 17270
rect 36544 17206 36596 17212
rect 36360 16992 36412 16998
rect 36360 16934 36412 16940
rect 36372 16114 36400 16934
rect 36360 16108 36412 16114
rect 36464 16096 36492 17206
rect 37200 16590 37228 19314
rect 38016 19304 38068 19310
rect 38014 19272 38016 19281
rect 38068 19272 38070 19281
rect 38014 19207 38070 19216
rect 37372 18420 37424 18426
rect 37372 18362 37424 18368
rect 37384 17202 37412 18362
rect 37464 18080 37516 18086
rect 37464 18022 37516 18028
rect 37476 17338 37504 18022
rect 37464 17332 37516 17338
rect 37464 17274 37516 17280
rect 37372 17196 37424 17202
rect 37372 17138 37424 17144
rect 37188 16584 37240 16590
rect 37188 16526 37240 16532
rect 36544 16108 36596 16114
rect 36464 16068 36544 16096
rect 36360 16050 36412 16056
rect 36544 16050 36596 16056
rect 36372 15638 36400 16050
rect 36360 15632 36412 15638
rect 36360 15574 36412 15580
rect 36360 14816 36412 14822
rect 36360 14758 36412 14764
rect 36372 14414 36400 14758
rect 36360 14408 36412 14414
rect 36360 14350 36412 14356
rect 37200 13938 37228 16526
rect 37372 15632 37424 15638
rect 37372 15574 37424 15580
rect 37384 13938 37412 15574
rect 38396 15162 38424 24006
rect 40132 23724 40184 23730
rect 40132 23666 40184 23672
rect 40144 22930 40172 23666
rect 40052 22902 40172 22930
rect 38936 22636 38988 22642
rect 38936 22578 38988 22584
rect 38948 22030 38976 22578
rect 40052 22094 40080 22902
rect 40224 22636 40276 22642
rect 40224 22578 40276 22584
rect 40132 22568 40184 22574
rect 40132 22510 40184 22516
rect 40144 22234 40172 22510
rect 40236 22386 40264 22578
rect 40604 22574 40632 24210
rect 41052 24200 41104 24206
rect 41052 24142 41104 24148
rect 41064 23798 41092 24142
rect 41052 23792 41104 23798
rect 41052 23734 41104 23740
rect 40592 22568 40644 22574
rect 40592 22510 40644 22516
rect 40236 22358 40356 22386
rect 40132 22228 40184 22234
rect 40132 22170 40184 22176
rect 40052 22066 40264 22094
rect 38936 22024 38988 22030
rect 38936 21966 38988 21972
rect 39028 22024 39080 22030
rect 39028 21966 39080 21972
rect 38476 20392 38528 20398
rect 38476 20334 38528 20340
rect 38488 19854 38516 20334
rect 38476 19848 38528 19854
rect 38476 19790 38528 19796
rect 38844 19712 38896 19718
rect 38844 19654 38896 19660
rect 38856 18290 38884 19654
rect 38844 18284 38896 18290
rect 38844 18226 38896 18232
rect 38750 17096 38806 17105
rect 38750 17031 38806 17040
rect 38764 16658 38792 17031
rect 38752 16652 38804 16658
rect 38752 16594 38804 16600
rect 38660 16584 38712 16590
rect 38660 16526 38712 16532
rect 38568 16176 38620 16182
rect 38568 16118 38620 16124
rect 38384 15156 38436 15162
rect 38384 15098 38436 15104
rect 37464 15020 37516 15026
rect 37464 14962 37516 14968
rect 37476 14414 37504 14962
rect 38016 14952 38068 14958
rect 38016 14894 38068 14900
rect 38028 14414 38056 14894
rect 37464 14408 37516 14414
rect 37464 14350 37516 14356
rect 38016 14408 38068 14414
rect 38016 14350 38068 14356
rect 38028 14074 38056 14350
rect 38396 14278 38424 15098
rect 38384 14272 38436 14278
rect 38384 14214 38436 14220
rect 38016 14068 38068 14074
rect 38016 14010 38068 14016
rect 37188 13932 37240 13938
rect 37188 13874 37240 13880
rect 37372 13932 37424 13938
rect 37372 13874 37424 13880
rect 37740 13252 37792 13258
rect 37740 13194 37792 13200
rect 37556 13184 37608 13190
rect 37556 13126 37608 13132
rect 37568 12986 37596 13126
rect 37188 12980 37240 12986
rect 37188 12922 37240 12928
rect 37556 12980 37608 12986
rect 37556 12922 37608 12928
rect 37200 12170 37228 12922
rect 37568 12753 37596 12922
rect 37752 12850 37780 13194
rect 38476 13184 38528 13190
rect 38476 13126 38528 13132
rect 37740 12844 37792 12850
rect 37740 12786 37792 12792
rect 37554 12744 37610 12753
rect 38488 12714 38516 13126
rect 37554 12679 37610 12688
rect 38476 12708 38528 12714
rect 37568 12442 37596 12679
rect 38476 12650 38528 12656
rect 38292 12640 38344 12646
rect 38292 12582 38344 12588
rect 37556 12436 37608 12442
rect 37556 12378 37608 12384
rect 38304 12238 38332 12582
rect 38292 12232 38344 12238
rect 38292 12174 38344 12180
rect 37188 12164 37240 12170
rect 37188 12106 37240 12112
rect 38304 11830 38332 12174
rect 38384 12164 38436 12170
rect 38384 12106 38436 12112
rect 36268 11824 36320 11830
rect 36268 11766 36320 11772
rect 38292 11824 38344 11830
rect 38292 11766 38344 11772
rect 38396 11762 38424 12106
rect 38384 11756 38436 11762
rect 38384 11698 38436 11704
rect 38476 11620 38528 11626
rect 38476 11562 38528 11568
rect 36176 11280 36228 11286
rect 36176 11222 36228 11228
rect 37370 11248 37426 11257
rect 37370 11183 37426 11192
rect 36084 11144 36136 11150
rect 36084 11086 36136 11092
rect 37384 10674 37412 11183
rect 38488 11082 38516 11562
rect 38580 11150 38608 16118
rect 38672 16114 38700 16526
rect 38660 16108 38712 16114
rect 38660 16050 38712 16056
rect 38752 14340 38804 14346
rect 38752 14282 38804 14288
rect 38764 13938 38792 14282
rect 38752 13932 38804 13938
rect 38752 13874 38804 13880
rect 38764 12918 38792 13874
rect 38752 12912 38804 12918
rect 38752 12854 38804 12860
rect 38752 12640 38804 12646
rect 38752 12582 38804 12588
rect 38764 12306 38792 12582
rect 38752 12300 38804 12306
rect 38752 12242 38804 12248
rect 38764 11830 38792 12242
rect 38752 11824 38804 11830
rect 38752 11766 38804 11772
rect 38568 11144 38620 11150
rect 38856 11132 38884 18226
rect 38948 16114 38976 21966
rect 39040 21690 39068 21966
rect 39028 21684 39080 21690
rect 39028 21626 39080 21632
rect 40236 20942 40264 22066
rect 40328 21962 40356 22358
rect 40316 21956 40368 21962
rect 40316 21898 40368 21904
rect 40224 20936 40276 20942
rect 40224 20878 40276 20884
rect 40500 20868 40552 20874
rect 40500 20810 40552 20816
rect 40512 20466 40540 20810
rect 40500 20460 40552 20466
rect 40500 20402 40552 20408
rect 39764 20392 39816 20398
rect 39764 20334 39816 20340
rect 39776 20262 39804 20334
rect 39764 20256 39816 20262
rect 39764 20198 39816 20204
rect 39776 19990 39804 20198
rect 39764 19984 39816 19990
rect 39764 19926 39816 19932
rect 40316 19168 40368 19174
rect 40316 19110 40368 19116
rect 40328 18834 40356 19110
rect 40316 18828 40368 18834
rect 40316 18770 40368 18776
rect 40328 18290 40356 18770
rect 40316 18284 40368 18290
rect 40316 18226 40368 18232
rect 40224 17740 40276 17746
rect 40224 17682 40276 17688
rect 40236 17542 40264 17682
rect 40512 17678 40540 20402
rect 40684 18760 40736 18766
rect 40684 18702 40736 18708
rect 40696 18290 40724 18702
rect 40684 18284 40736 18290
rect 40684 18226 40736 18232
rect 40500 17672 40552 17678
rect 40500 17614 40552 17620
rect 40224 17536 40276 17542
rect 40222 17504 40224 17513
rect 40276 17504 40278 17513
rect 40222 17439 40278 17448
rect 40512 17202 40540 17614
rect 40500 17196 40552 17202
rect 40500 17138 40552 17144
rect 40512 17082 40540 17138
rect 40512 17054 40632 17082
rect 40040 16992 40092 16998
rect 40040 16934 40092 16940
rect 40052 16697 40080 16934
rect 40038 16688 40094 16697
rect 40038 16623 40094 16632
rect 39212 16448 39264 16454
rect 39212 16390 39264 16396
rect 38936 16108 38988 16114
rect 38936 16050 38988 16056
rect 39224 15910 39252 16390
rect 39854 16008 39910 16017
rect 39854 15943 39910 15952
rect 39212 15904 39264 15910
rect 39212 15846 39264 15852
rect 39868 15706 39896 15943
rect 39856 15700 39908 15706
rect 39856 15642 39908 15648
rect 40604 15502 40632 17054
rect 41432 16574 41460 36178
rect 41892 36106 41920 36722
rect 42628 36718 42656 37062
rect 42706 36816 42762 36825
rect 43732 36786 43760 37130
rect 46124 36786 46152 37130
rect 46572 37120 46624 37126
rect 46572 37062 46624 37068
rect 46768 37074 46796 37334
rect 46860 37210 46888 39222
rect 48318 39200 48374 40000
rect 50250 39200 50306 40000
rect 52182 39200 52238 40000
rect 54114 39200 54170 40000
rect 56046 39200 56102 40000
rect 57978 39200 58034 40000
rect 59910 39200 59966 40000
rect 48332 37346 48360 39200
rect 48596 37460 48648 37466
rect 48596 37402 48648 37408
rect 47032 37324 47084 37330
rect 48332 37318 48452 37346
rect 47032 37266 47084 37272
rect 46860 37194 46980 37210
rect 46860 37188 46992 37194
rect 46860 37182 46940 37188
rect 46940 37130 46992 37136
rect 46388 36848 46440 36854
rect 46388 36790 46440 36796
rect 42706 36751 42708 36760
rect 42760 36751 42762 36760
rect 43720 36780 43772 36786
rect 42708 36722 42760 36728
rect 43720 36722 43772 36728
rect 46112 36780 46164 36786
rect 46112 36722 46164 36728
rect 42616 36712 42668 36718
rect 42616 36654 42668 36660
rect 42628 36582 42656 36654
rect 42616 36576 42668 36582
rect 42616 36518 42668 36524
rect 42984 36576 43036 36582
rect 42984 36518 43036 36524
rect 42996 36174 43024 36518
rect 46124 36310 46152 36722
rect 46112 36304 46164 36310
rect 46112 36246 46164 36252
rect 42984 36168 43036 36174
rect 42984 36110 43036 36116
rect 41880 36100 41932 36106
rect 41880 36042 41932 36048
rect 44640 36100 44692 36106
rect 44640 36042 44692 36048
rect 43628 35624 43680 35630
rect 43628 35566 43680 35572
rect 43640 35290 43668 35566
rect 43628 35284 43680 35290
rect 43628 35226 43680 35232
rect 43260 35148 43312 35154
rect 43260 35090 43312 35096
rect 42892 34604 42944 34610
rect 42892 34546 42944 34552
rect 43168 34604 43220 34610
rect 43168 34546 43220 34552
rect 42904 34134 42932 34546
rect 43180 34202 43208 34546
rect 43272 34474 43300 35090
rect 43352 35080 43404 35086
rect 43352 35022 43404 35028
rect 43260 34468 43312 34474
rect 43260 34410 43312 34416
rect 43168 34196 43220 34202
rect 43168 34138 43220 34144
rect 42892 34128 42944 34134
rect 42892 34070 42944 34076
rect 41788 34060 41840 34066
rect 41788 34002 41840 34008
rect 41800 33522 41828 34002
rect 42904 33998 42932 34070
rect 42892 33992 42944 33998
rect 42892 33934 42944 33940
rect 42616 33924 42668 33930
rect 42616 33866 42668 33872
rect 42628 33522 42656 33866
rect 43180 33862 43208 34138
rect 43364 33998 43392 35022
rect 43352 33992 43404 33998
rect 43352 33934 43404 33940
rect 43168 33856 43220 33862
rect 43168 33798 43220 33804
rect 43352 33856 43404 33862
rect 43352 33798 43404 33804
rect 43364 33522 43392 33798
rect 41788 33516 41840 33522
rect 41788 33458 41840 33464
rect 42616 33516 42668 33522
rect 42616 33458 42668 33464
rect 43352 33516 43404 33522
rect 43352 33458 43404 33464
rect 41800 32366 41828 33458
rect 43352 32428 43404 32434
rect 43352 32370 43404 32376
rect 41788 32360 41840 32366
rect 41788 32302 41840 32308
rect 43364 32026 43392 32370
rect 43352 32020 43404 32026
rect 43352 31962 43404 31968
rect 44364 30728 44416 30734
rect 44364 30670 44416 30676
rect 44376 30394 44404 30670
rect 44364 30388 44416 30394
rect 44364 30330 44416 30336
rect 43076 30320 43128 30326
rect 43076 30262 43128 30268
rect 42432 30252 42484 30258
rect 42432 30194 42484 30200
rect 42444 29510 42472 30194
rect 42524 30184 42576 30190
rect 42524 30126 42576 30132
rect 42536 29850 42564 30126
rect 42524 29844 42576 29850
rect 42524 29786 42576 29792
rect 42432 29504 42484 29510
rect 42432 29446 42484 29452
rect 42536 28762 42564 29786
rect 43088 29578 43116 30262
rect 44272 30252 44324 30258
rect 44272 30194 44324 30200
rect 44284 29714 44312 30194
rect 44272 29708 44324 29714
rect 44272 29650 44324 29656
rect 43076 29572 43128 29578
rect 43076 29514 43128 29520
rect 43088 29170 43116 29514
rect 43076 29164 43128 29170
rect 43076 29106 43128 29112
rect 42892 29096 42944 29102
rect 42892 29038 42944 29044
rect 42524 28756 42576 28762
rect 42524 28698 42576 28704
rect 42904 28626 42932 29038
rect 42892 28620 42944 28626
rect 42892 28562 42944 28568
rect 42340 28552 42392 28558
rect 42340 28494 42392 28500
rect 41880 28416 41932 28422
rect 41880 28358 41932 28364
rect 41892 28082 41920 28358
rect 41880 28076 41932 28082
rect 41880 28018 41932 28024
rect 42352 28014 42380 28494
rect 42904 28082 42932 28562
rect 43088 28218 43116 29106
rect 43076 28212 43128 28218
rect 43076 28154 43128 28160
rect 42892 28076 42944 28082
rect 42892 28018 42944 28024
rect 42340 28008 42392 28014
rect 42340 27950 42392 27956
rect 42352 27334 42380 27950
rect 42340 27328 42392 27334
rect 42340 27270 42392 27276
rect 44272 26988 44324 26994
rect 44272 26930 44324 26936
rect 44180 26920 44232 26926
rect 44180 26862 44232 26868
rect 43168 26512 43220 26518
rect 43168 26454 43220 26460
rect 41880 25288 41932 25294
rect 41880 25230 41932 25236
rect 42800 25288 42852 25294
rect 42800 25230 42852 25236
rect 41604 25220 41656 25226
rect 41604 25162 41656 25168
rect 41616 24818 41644 25162
rect 41892 24818 41920 25230
rect 41604 24812 41656 24818
rect 41604 24754 41656 24760
rect 41880 24812 41932 24818
rect 41880 24754 41932 24760
rect 41616 23526 41644 24754
rect 42812 24750 42840 25230
rect 42800 24744 42852 24750
rect 42800 24686 42852 24692
rect 41604 23520 41656 23526
rect 41604 23462 41656 23468
rect 42800 23112 42852 23118
rect 42800 23054 42852 23060
rect 42524 22636 42576 22642
rect 42524 22578 42576 22584
rect 42536 22234 42564 22578
rect 42812 22234 42840 23054
rect 42984 22636 43036 22642
rect 42984 22578 43036 22584
rect 42892 22432 42944 22438
rect 42892 22374 42944 22380
rect 42524 22228 42576 22234
rect 42524 22170 42576 22176
rect 42800 22228 42852 22234
rect 42800 22170 42852 22176
rect 42904 22030 42932 22374
rect 42996 22030 43024 22578
rect 42892 22024 42944 22030
rect 42892 21966 42944 21972
rect 42984 22024 43036 22030
rect 42984 21966 43036 21972
rect 42996 21146 43024 21966
rect 42984 21140 43036 21146
rect 42984 21082 43036 21088
rect 41972 20936 42024 20942
rect 41972 20878 42024 20884
rect 42156 20936 42208 20942
rect 42156 20878 42208 20884
rect 41984 20602 42012 20878
rect 41972 20596 42024 20602
rect 41972 20538 42024 20544
rect 41984 20330 42012 20538
rect 42168 20534 42196 20878
rect 42156 20528 42208 20534
rect 42156 20470 42208 20476
rect 41972 20324 42024 20330
rect 41972 20266 42024 20272
rect 42800 20052 42852 20058
rect 42800 19994 42852 20000
rect 42708 19780 42760 19786
rect 42708 19722 42760 19728
rect 41788 19712 41840 19718
rect 41788 19654 41840 19660
rect 41800 19174 41828 19654
rect 42720 19378 42748 19722
rect 42708 19372 42760 19378
rect 42708 19314 42760 19320
rect 41788 19168 41840 19174
rect 41788 19110 41840 19116
rect 41696 18760 41748 18766
rect 41800 18737 41828 19110
rect 41696 18702 41748 18708
rect 41786 18728 41842 18737
rect 41708 17814 41736 18702
rect 41786 18663 41842 18672
rect 42720 18426 42748 19314
rect 42812 19310 42840 19994
rect 42800 19304 42852 19310
rect 42800 19246 42852 19252
rect 42812 18902 42840 19246
rect 42800 18896 42852 18902
rect 42800 18838 42852 18844
rect 42708 18420 42760 18426
rect 42708 18362 42760 18368
rect 41696 17808 41748 17814
rect 41696 17750 41748 17756
rect 41432 16546 41644 16574
rect 40592 15496 40644 15502
rect 40592 15438 40644 15444
rect 40038 15192 40094 15201
rect 40038 15127 40094 15136
rect 40052 14618 40080 15127
rect 40604 15026 40632 15438
rect 40592 15020 40644 15026
rect 40592 14962 40644 14968
rect 40776 14816 40828 14822
rect 40776 14758 40828 14764
rect 40040 14612 40092 14618
rect 40040 14554 40092 14560
rect 40052 14482 40080 14554
rect 40040 14476 40092 14482
rect 40040 14418 40092 14424
rect 40788 14414 40816 14758
rect 40776 14408 40828 14414
rect 40696 14368 40776 14396
rect 39120 14000 39172 14006
rect 39120 13942 39172 13948
rect 39132 11762 39160 13942
rect 40696 12238 40724 14368
rect 40776 14350 40828 14356
rect 40776 13728 40828 13734
rect 40776 13670 40828 13676
rect 40788 13326 40816 13670
rect 41144 13388 41196 13394
rect 41144 13330 41196 13336
rect 40776 13320 40828 13326
rect 40776 13262 40828 13268
rect 40788 12850 40816 13262
rect 40776 12844 40828 12850
rect 40776 12786 40828 12792
rect 41156 12782 41184 13330
rect 41144 12776 41196 12782
rect 41144 12718 41196 12724
rect 40684 12232 40736 12238
rect 40314 12200 40370 12209
rect 40684 12174 40736 12180
rect 41144 12232 41196 12238
rect 41144 12174 41196 12180
rect 40314 12135 40370 12144
rect 39120 11756 39172 11762
rect 39040 11716 39120 11744
rect 39040 11218 39068 11716
rect 39120 11698 39172 11704
rect 39304 11552 39356 11558
rect 39304 11494 39356 11500
rect 39856 11552 39908 11558
rect 39856 11494 39908 11500
rect 39028 11212 39080 11218
rect 39028 11154 39080 11160
rect 38936 11144 38988 11150
rect 38856 11104 38936 11132
rect 38568 11086 38620 11092
rect 38936 11086 38988 11092
rect 38476 11076 38528 11082
rect 38476 11018 38528 11024
rect 37372 10668 37424 10674
rect 37372 10610 37424 10616
rect 38292 10600 38344 10606
rect 38292 10542 38344 10548
rect 36360 10260 36412 10266
rect 36360 10202 36412 10208
rect 35900 9648 35952 9654
rect 35900 9590 35952 9596
rect 35912 9489 35940 9590
rect 36372 9586 36400 10202
rect 36544 10056 36596 10062
rect 36544 9998 36596 10004
rect 36360 9580 36412 9586
rect 36360 9522 36412 9528
rect 35898 9480 35954 9489
rect 35898 9415 35954 9424
rect 35912 9042 35940 9415
rect 36372 9178 36400 9522
rect 36556 9518 36584 9998
rect 36728 9920 36780 9926
rect 36728 9862 36780 9868
rect 36544 9512 36596 9518
rect 36544 9454 36596 9460
rect 36360 9172 36412 9178
rect 36360 9114 36412 9120
rect 35900 9036 35952 9042
rect 35900 8978 35952 8984
rect 36268 9036 36320 9042
rect 36268 8978 36320 8984
rect 36280 8566 36308 8978
rect 36556 8634 36584 9454
rect 36740 9110 36768 9862
rect 36728 9104 36780 9110
rect 36728 9046 36780 9052
rect 38304 9042 38332 10542
rect 38488 9994 38516 11018
rect 38580 10010 38608 11086
rect 38948 10674 38976 11086
rect 38936 10668 38988 10674
rect 38936 10610 38988 10616
rect 38936 10532 38988 10538
rect 38936 10474 38988 10480
rect 38580 9994 38700 10010
rect 38476 9988 38528 9994
rect 38580 9988 38712 9994
rect 38580 9982 38660 9988
rect 38476 9930 38528 9936
rect 38660 9930 38712 9936
rect 37924 9036 37976 9042
rect 37924 8978 37976 8984
rect 38292 9036 38344 9042
rect 38292 8978 38344 8984
rect 37556 8968 37608 8974
rect 37556 8910 37608 8916
rect 36544 8628 36596 8634
rect 36544 8570 36596 8576
rect 36268 8560 36320 8566
rect 36268 8502 36320 8508
rect 37568 8498 37596 8910
rect 37936 8498 37964 8978
rect 37556 8492 37608 8498
rect 37556 8434 37608 8440
rect 37924 8492 37976 8498
rect 37924 8434 37976 8440
rect 38108 8492 38160 8498
rect 38108 8434 38160 8440
rect 35900 7880 35952 7886
rect 35900 7822 35952 7828
rect 35808 7744 35860 7750
rect 35808 7686 35860 7692
rect 35716 7404 35768 7410
rect 35716 7346 35768 7352
rect 35624 7336 35676 7342
rect 35624 7278 35676 7284
rect 35624 7200 35676 7206
rect 35624 7142 35676 7148
rect 31024 6792 31076 6798
rect 31024 6734 31076 6740
rect 31484 6792 31536 6798
rect 31484 6734 31536 6740
rect 34704 6792 34756 6798
rect 34704 6734 34756 6740
rect 35532 6792 35584 6798
rect 35532 6734 35584 6740
rect 31036 6322 31064 6734
rect 31208 6656 31260 6662
rect 31208 6598 31260 6604
rect 31024 6316 31076 6322
rect 31024 6258 31076 6264
rect 29644 5772 29696 5778
rect 29644 5714 29696 5720
rect 31220 5710 31248 6598
rect 31496 6322 31524 6734
rect 33600 6452 33652 6458
rect 33600 6394 33652 6400
rect 31484 6316 31536 6322
rect 31484 6258 31536 6264
rect 31392 6112 31444 6118
rect 31392 6054 31444 6060
rect 32036 6112 32088 6118
rect 32036 6054 32088 6060
rect 31404 5914 31432 6054
rect 32048 5914 32076 6054
rect 31392 5908 31444 5914
rect 31392 5850 31444 5856
rect 32036 5908 32088 5914
rect 32036 5850 32088 5856
rect 31404 5710 31432 5850
rect 31944 5840 31996 5846
rect 31944 5782 31996 5788
rect 31956 5710 31984 5782
rect 33612 5710 33640 6394
rect 34716 6322 34744 6734
rect 34704 6316 34756 6322
rect 34704 6258 34756 6264
rect 35440 6112 35492 6118
rect 35440 6054 35492 6060
rect 34934 6012 35242 6032
rect 34934 6010 34940 6012
rect 34996 6010 35020 6012
rect 35076 6010 35100 6012
rect 35156 6010 35180 6012
rect 35236 6010 35242 6012
rect 34996 5958 34998 6010
rect 35178 5958 35180 6010
rect 34934 5956 34940 5958
rect 34996 5956 35020 5958
rect 35076 5956 35100 5958
rect 35156 5956 35180 5958
rect 35236 5956 35242 5958
rect 34934 5936 35242 5956
rect 35452 5778 35480 6054
rect 35440 5772 35492 5778
rect 35440 5714 35492 5720
rect 35544 5710 35572 6734
rect 31208 5704 31260 5710
rect 31208 5646 31260 5652
rect 31392 5704 31444 5710
rect 31392 5646 31444 5652
rect 31944 5704 31996 5710
rect 31944 5646 31996 5652
rect 33140 5704 33192 5710
rect 33140 5646 33192 5652
rect 33600 5704 33652 5710
rect 33600 5646 33652 5652
rect 35532 5704 35584 5710
rect 35532 5646 35584 5652
rect 30472 5568 30524 5574
rect 30472 5510 30524 5516
rect 31576 5568 31628 5574
rect 31576 5510 31628 5516
rect 32404 5568 32456 5574
rect 32404 5510 32456 5516
rect 30484 5234 30512 5510
rect 31588 5302 31616 5510
rect 31576 5296 31628 5302
rect 31576 5238 31628 5244
rect 32416 5234 32444 5510
rect 33152 5302 33180 5646
rect 33232 5568 33284 5574
rect 33232 5510 33284 5516
rect 33140 5296 33192 5302
rect 33140 5238 33192 5244
rect 30472 5228 30524 5234
rect 30472 5170 30524 5176
rect 32404 5228 32456 5234
rect 32404 5170 32456 5176
rect 32220 5160 32272 5166
rect 32220 5102 32272 5108
rect 32864 5160 32916 5166
rect 32864 5102 32916 5108
rect 31576 5024 31628 5030
rect 31576 4966 31628 4972
rect 31588 4622 31616 4966
rect 31576 4616 31628 4622
rect 31576 4558 31628 4564
rect 29276 4004 29328 4010
rect 29276 3946 29328 3952
rect 28540 3596 28592 3602
rect 28540 3538 28592 3544
rect 28908 3596 28960 3602
rect 28908 3538 28960 3544
rect 28552 3398 28580 3538
rect 32232 3534 32260 5102
rect 32876 4554 32904 5102
rect 33152 4826 33180 5238
rect 33244 5234 33272 5510
rect 33232 5228 33284 5234
rect 33232 5170 33284 5176
rect 34934 4924 35242 4944
rect 34934 4922 34940 4924
rect 34996 4922 35020 4924
rect 35076 4922 35100 4924
rect 35156 4922 35180 4924
rect 35236 4922 35242 4924
rect 34996 4870 34998 4922
rect 35178 4870 35180 4922
rect 34934 4868 34940 4870
rect 34996 4868 35020 4870
rect 35076 4868 35100 4870
rect 35156 4868 35180 4870
rect 35236 4868 35242 4870
rect 34934 4848 35242 4868
rect 33140 4820 33192 4826
rect 33140 4762 33192 4768
rect 32864 4548 32916 4554
rect 32864 4490 32916 4496
rect 33140 4480 33192 4486
rect 33140 4422 33192 4428
rect 33152 4146 33180 4422
rect 33140 4140 33192 4146
rect 33140 4082 33192 4088
rect 33600 4140 33652 4146
rect 33600 4082 33652 4088
rect 33692 4140 33744 4146
rect 35636 4128 35664 7142
rect 35820 6798 35848 7686
rect 35912 7478 35940 7822
rect 37740 7812 37792 7818
rect 37740 7754 37792 7760
rect 36452 7744 36504 7750
rect 36452 7686 36504 7692
rect 35900 7472 35952 7478
rect 35900 7414 35952 7420
rect 35912 7002 35940 7414
rect 35900 6996 35952 7002
rect 35900 6938 35952 6944
rect 35808 6792 35860 6798
rect 35808 6734 35860 6740
rect 35820 6390 35848 6734
rect 35808 6384 35860 6390
rect 35808 6326 35860 6332
rect 35716 6316 35768 6322
rect 35716 6258 35768 6264
rect 35728 5778 35756 6258
rect 35716 5772 35768 5778
rect 35716 5714 35768 5720
rect 35900 5568 35952 5574
rect 35900 5510 35952 5516
rect 35912 5234 35940 5510
rect 35900 5228 35952 5234
rect 35900 5170 35952 5176
rect 36464 4146 36492 7686
rect 37004 6656 37056 6662
rect 37004 6598 37056 6604
rect 37016 6322 37044 6598
rect 37004 6316 37056 6322
rect 37004 6258 37056 6264
rect 37464 6316 37516 6322
rect 37464 6258 37516 6264
rect 37016 5710 37044 6258
rect 37476 6186 37504 6258
rect 37752 6254 37780 7754
rect 38120 6662 38148 8434
rect 38660 7948 38712 7954
rect 38660 7890 38712 7896
rect 38476 7200 38528 7206
rect 38476 7142 38528 7148
rect 38488 6730 38516 7142
rect 38476 6724 38528 6730
rect 38476 6666 38528 6672
rect 38108 6656 38160 6662
rect 38108 6598 38160 6604
rect 37740 6248 37792 6254
rect 37740 6190 37792 6196
rect 37464 6180 37516 6186
rect 37464 6122 37516 6128
rect 37476 5710 37504 6122
rect 37832 6112 37884 6118
rect 37832 6054 37884 6060
rect 37844 5710 37872 6054
rect 37004 5704 37056 5710
rect 37004 5646 37056 5652
rect 37464 5704 37516 5710
rect 37464 5646 37516 5652
rect 37832 5704 37884 5710
rect 37832 5646 37884 5652
rect 37096 5568 37148 5574
rect 37096 5510 37148 5516
rect 37832 5568 37884 5574
rect 37832 5510 37884 5516
rect 37108 4554 37136 5510
rect 37648 4820 37700 4826
rect 37648 4762 37700 4768
rect 37280 4684 37332 4690
rect 37280 4626 37332 4632
rect 37096 4548 37148 4554
rect 37096 4490 37148 4496
rect 35808 4140 35860 4146
rect 35636 4100 35808 4128
rect 33692 4082 33744 4088
rect 35808 4082 35860 4088
rect 36452 4140 36504 4146
rect 36452 4082 36504 4088
rect 33232 3936 33284 3942
rect 33232 3878 33284 3884
rect 33048 3596 33100 3602
rect 33048 3538 33100 3544
rect 32220 3528 32272 3534
rect 32220 3470 32272 3476
rect 28540 3392 28592 3398
rect 28540 3334 28592 3340
rect 33060 3058 33088 3538
rect 33244 3058 33272 3878
rect 33612 3534 33640 4082
rect 33704 3670 33732 4082
rect 34934 3836 35242 3856
rect 34934 3834 34940 3836
rect 34996 3834 35020 3836
rect 35076 3834 35100 3836
rect 35156 3834 35180 3836
rect 35236 3834 35242 3836
rect 34996 3782 34998 3834
rect 35178 3782 35180 3834
rect 34934 3780 34940 3782
rect 34996 3780 35020 3782
rect 35076 3780 35100 3782
rect 35156 3780 35180 3782
rect 35236 3780 35242 3782
rect 34934 3760 35242 3780
rect 33692 3664 33744 3670
rect 33692 3606 33744 3612
rect 33600 3528 33652 3534
rect 33600 3470 33652 3476
rect 33876 3528 33928 3534
rect 33876 3470 33928 3476
rect 33888 3126 33916 3470
rect 34244 3460 34296 3466
rect 34244 3402 34296 3408
rect 34256 3126 34284 3402
rect 33876 3120 33928 3126
rect 33876 3062 33928 3068
rect 34244 3120 34296 3126
rect 34244 3062 34296 3068
rect 35820 3058 35848 4082
rect 36544 3936 36596 3942
rect 36544 3878 36596 3884
rect 36556 3738 36584 3878
rect 36544 3732 36596 3738
rect 36544 3674 36596 3680
rect 36360 3596 36412 3602
rect 36360 3538 36412 3544
rect 36372 3194 36400 3538
rect 37108 3534 37136 4490
rect 37292 3534 37320 4626
rect 37660 4622 37688 4762
rect 37844 4622 37872 5510
rect 38120 4826 38148 6598
rect 38672 6458 38700 7890
rect 38948 7750 38976 10474
rect 39316 10266 39344 11494
rect 39868 11082 39896 11494
rect 40328 11218 40356 12135
rect 41052 11348 41104 11354
rect 41052 11290 41104 11296
rect 40316 11212 40368 11218
rect 40316 11154 40368 11160
rect 39856 11076 39908 11082
rect 39856 11018 39908 11024
rect 39868 10742 39896 11018
rect 39856 10736 39908 10742
rect 39856 10678 39908 10684
rect 40328 10674 40356 11154
rect 40316 10668 40368 10674
rect 40316 10610 40368 10616
rect 39856 10464 39908 10470
rect 39856 10406 39908 10412
rect 40960 10464 41012 10470
rect 40960 10406 41012 10412
rect 39304 10260 39356 10266
rect 39304 10202 39356 10208
rect 39118 8936 39174 8945
rect 39118 8871 39174 8880
rect 39132 8634 39160 8871
rect 39672 8832 39724 8838
rect 39672 8774 39724 8780
rect 39120 8628 39172 8634
rect 39120 8570 39172 8576
rect 39120 8424 39172 8430
rect 39120 8366 39172 8372
rect 39132 7886 39160 8366
rect 39684 8362 39712 8774
rect 39672 8356 39724 8362
rect 39672 8298 39724 8304
rect 39684 7886 39712 8298
rect 39868 7954 39896 10406
rect 40972 10062 41000 10406
rect 41064 10266 41092 11290
rect 41156 10742 41184 12174
rect 41420 11008 41472 11014
rect 41420 10950 41472 10956
rect 41144 10736 41196 10742
rect 41144 10678 41196 10684
rect 41052 10260 41104 10266
rect 41052 10202 41104 10208
rect 41064 10062 41092 10202
rect 41432 10062 41460 10950
rect 40960 10056 41012 10062
rect 40960 9998 41012 10004
rect 41052 10056 41104 10062
rect 41052 9998 41104 10004
rect 41420 10056 41472 10062
rect 41420 9998 41472 10004
rect 41512 9920 41564 9926
rect 41512 9862 41564 9868
rect 41524 9654 41552 9862
rect 41512 9648 41564 9654
rect 41512 9590 41564 9596
rect 40132 9104 40184 9110
rect 40132 9046 40184 9052
rect 40144 8498 40172 9046
rect 41052 8968 41104 8974
rect 41052 8910 41104 8916
rect 41064 8498 41092 8910
rect 40132 8492 40184 8498
rect 40132 8434 40184 8440
rect 41052 8492 41104 8498
rect 41052 8434 41104 8440
rect 41064 7954 41092 8434
rect 39856 7948 39908 7954
rect 39856 7890 39908 7896
rect 41052 7948 41104 7954
rect 41052 7890 41104 7896
rect 39120 7880 39172 7886
rect 39120 7822 39172 7828
rect 39672 7880 39724 7886
rect 39672 7822 39724 7828
rect 38936 7744 38988 7750
rect 38936 7686 38988 7692
rect 38948 7410 38976 7686
rect 38936 7404 38988 7410
rect 38936 7346 38988 7352
rect 39684 7342 39712 7822
rect 39672 7336 39724 7342
rect 39670 7304 39672 7313
rect 39724 7304 39726 7313
rect 39670 7239 39726 7248
rect 38844 6928 38896 6934
rect 38844 6870 38896 6876
rect 40132 6928 40184 6934
rect 40132 6870 40184 6876
rect 38856 6458 38884 6870
rect 39948 6792 40000 6798
rect 39948 6734 40000 6740
rect 38660 6452 38712 6458
rect 38660 6394 38712 6400
rect 38844 6452 38896 6458
rect 38844 6394 38896 6400
rect 38672 5098 38700 6394
rect 38856 6322 38884 6394
rect 39960 6322 39988 6734
rect 40040 6724 40092 6730
rect 40040 6666 40092 6672
rect 38844 6316 38896 6322
rect 38844 6258 38896 6264
rect 39948 6316 40000 6322
rect 39948 6258 40000 6264
rect 40052 5710 40080 6666
rect 40144 6186 40172 6870
rect 40224 6248 40276 6254
rect 40224 6190 40276 6196
rect 40408 6248 40460 6254
rect 40408 6190 40460 6196
rect 40132 6180 40184 6186
rect 40132 6122 40184 6128
rect 40236 5710 40264 6190
rect 40040 5704 40092 5710
rect 40040 5646 40092 5652
rect 40224 5704 40276 5710
rect 40224 5646 40276 5652
rect 38660 5092 38712 5098
rect 38660 5034 38712 5040
rect 38108 4820 38160 4826
rect 38108 4762 38160 4768
rect 40420 4622 40448 6190
rect 40500 5568 40552 5574
rect 40500 5510 40552 5516
rect 40868 5568 40920 5574
rect 40868 5510 40920 5516
rect 40512 5234 40540 5510
rect 40880 5234 40908 5510
rect 40500 5228 40552 5234
rect 40500 5170 40552 5176
rect 40868 5228 40920 5234
rect 40868 5170 40920 5176
rect 41236 5160 41288 5166
rect 41236 5102 41288 5108
rect 40500 5092 40552 5098
rect 40500 5034 40552 5040
rect 37556 4616 37608 4622
rect 37556 4558 37608 4564
rect 37648 4616 37700 4622
rect 37648 4558 37700 4564
rect 37832 4616 37884 4622
rect 37832 4558 37884 4564
rect 40408 4616 40460 4622
rect 40408 4558 40460 4564
rect 37568 4078 37596 4558
rect 37844 4078 37872 4558
rect 40512 4146 40540 5034
rect 40684 4616 40736 4622
rect 40684 4558 40736 4564
rect 40500 4140 40552 4146
rect 40500 4082 40552 4088
rect 40696 4078 40724 4558
rect 40868 4480 40920 4486
rect 40868 4422 40920 4428
rect 40880 4214 40908 4422
rect 40868 4208 40920 4214
rect 40868 4150 40920 4156
rect 37372 4072 37424 4078
rect 37372 4014 37424 4020
rect 37556 4072 37608 4078
rect 37556 4014 37608 4020
rect 37832 4072 37884 4078
rect 37832 4014 37884 4020
rect 40684 4072 40736 4078
rect 40684 4014 40736 4020
rect 37096 3528 37148 3534
rect 37096 3470 37148 3476
rect 37280 3528 37332 3534
rect 37280 3470 37332 3476
rect 37384 3466 37412 4014
rect 37464 3936 37516 3942
rect 37464 3878 37516 3884
rect 37476 3534 37504 3878
rect 37740 3664 37792 3670
rect 37740 3606 37792 3612
rect 37464 3528 37516 3534
rect 37464 3470 37516 3476
rect 37372 3460 37424 3466
rect 37372 3402 37424 3408
rect 36360 3188 36412 3194
rect 36360 3130 36412 3136
rect 37384 3058 37412 3402
rect 33048 3052 33100 3058
rect 33048 2994 33100 3000
rect 33232 3052 33284 3058
rect 33232 2994 33284 3000
rect 33416 3052 33468 3058
rect 33416 2994 33468 3000
rect 35808 3052 35860 3058
rect 35808 2994 35860 3000
rect 37372 3052 37424 3058
rect 37372 2994 37424 3000
rect 32588 2916 32640 2922
rect 32588 2858 32640 2864
rect 31576 2848 31628 2854
rect 31576 2790 31628 2796
rect 31588 2446 31616 2790
rect 32600 2446 32628 2858
rect 33060 2650 33088 2994
rect 33048 2644 33100 2650
rect 33048 2586 33100 2592
rect 32680 2576 32732 2582
rect 32680 2518 32732 2524
rect 27712 2440 27764 2446
rect 27712 2382 27764 2388
rect 28448 2440 28500 2446
rect 28448 2382 28500 2388
rect 31576 2440 31628 2446
rect 31576 2382 31628 2388
rect 32588 2440 32640 2446
rect 32588 2382 32640 2388
rect 26240 1760 26292 1766
rect 26160 1708 26240 1714
rect 26160 1702 26292 1708
rect 26976 1760 27028 1766
rect 26976 1702 27028 1708
rect 27528 1760 27580 1766
rect 27528 1702 27580 1708
rect 26160 1686 26280 1702
rect 25792 870 25912 898
rect 25792 800 25820 870
rect 18 0 74 800
rect 1950 0 2006 800
rect 3882 0 3938 800
rect 5814 0 5870 800
rect 7746 0 7802 800
rect 9678 0 9734 800
rect 11610 0 11666 800
rect 13542 0 13598 800
rect 15474 0 15530 800
rect 18050 0 18106 800
rect 19982 0 20038 800
rect 21914 0 21970 800
rect 23846 0 23902 800
rect 25778 0 25834 800
rect 25884 762 25912 870
rect 26160 762 26188 1686
rect 27724 800 27752 2382
rect 29644 2372 29696 2378
rect 29644 2314 29696 2320
rect 29656 800 29684 2314
rect 30104 2304 30156 2310
rect 30104 2246 30156 2252
rect 30116 1902 30144 2246
rect 30104 1896 30156 1902
rect 30104 1838 30156 1844
rect 31588 800 31616 2382
rect 32692 2310 32720 2518
rect 33244 2446 33272 2994
rect 33428 2854 33456 2994
rect 37476 2990 37504 3470
rect 37752 3398 37780 3606
rect 40880 3534 40908 4150
rect 41248 4026 41276 5102
rect 41512 5024 41564 5030
rect 41512 4966 41564 4972
rect 41524 4622 41552 4966
rect 41328 4616 41380 4622
rect 41328 4558 41380 4564
rect 41512 4616 41564 4622
rect 41512 4558 41564 4564
rect 41340 4146 41368 4558
rect 41524 4146 41552 4558
rect 41328 4140 41380 4146
rect 41328 4082 41380 4088
rect 41512 4140 41564 4146
rect 41512 4082 41564 4088
rect 41248 3998 41460 4026
rect 41432 3942 41460 3998
rect 41052 3936 41104 3942
rect 41052 3878 41104 3884
rect 41420 3936 41472 3942
rect 41420 3878 41472 3884
rect 41064 3534 41092 3878
rect 41616 3670 41644 16546
rect 42524 16516 42576 16522
rect 42524 16458 42576 16464
rect 41972 16448 42024 16454
rect 41972 16390 42024 16396
rect 41984 15502 42012 16390
rect 42536 15502 42564 16458
rect 42800 16108 42852 16114
rect 42800 16050 42852 16056
rect 42812 15502 42840 16050
rect 41972 15496 42024 15502
rect 41970 15464 41972 15473
rect 42524 15496 42576 15502
rect 42024 15464 42026 15473
rect 42524 15438 42576 15444
rect 42800 15496 42852 15502
rect 42800 15438 42852 15444
rect 41970 15399 42026 15408
rect 42340 14272 42392 14278
rect 42340 14214 42392 14220
rect 42352 13326 42380 14214
rect 42340 13320 42392 13326
rect 42340 13262 42392 13268
rect 42352 12714 42380 13262
rect 42892 13252 42944 13258
rect 42892 13194 42944 13200
rect 42904 12918 42932 13194
rect 42892 12912 42944 12918
rect 42892 12854 42944 12860
rect 42340 12708 42392 12714
rect 42340 12650 42392 12656
rect 43180 12434 43208 26454
rect 44192 26042 44220 26862
rect 44284 26586 44312 26930
rect 44272 26580 44324 26586
rect 44272 26522 44324 26528
rect 44180 26036 44232 26042
rect 44180 25978 44232 25984
rect 43812 25900 43864 25906
rect 43812 25842 43864 25848
rect 43720 25832 43772 25838
rect 43720 25774 43772 25780
rect 43732 25294 43760 25774
rect 43824 25498 43852 25842
rect 43812 25492 43864 25498
rect 43812 25434 43864 25440
rect 43720 25288 43772 25294
rect 43720 25230 43772 25236
rect 43824 24342 43852 25434
rect 44180 25152 44232 25158
rect 44180 25094 44232 25100
rect 44192 24818 44220 25094
rect 44180 24812 44232 24818
rect 44180 24754 44232 24760
rect 44548 24812 44600 24818
rect 44548 24754 44600 24760
rect 43812 24336 43864 24342
rect 43812 24278 43864 24284
rect 44192 24206 44220 24754
rect 44560 24410 44588 24754
rect 44548 24404 44600 24410
rect 44548 24346 44600 24352
rect 43812 24200 43864 24206
rect 44180 24200 44232 24206
rect 43864 24160 43944 24188
rect 43812 24142 43864 24148
rect 43536 24064 43588 24070
rect 43536 24006 43588 24012
rect 43548 23798 43576 24006
rect 43536 23792 43588 23798
rect 43536 23734 43588 23740
rect 43548 22982 43576 23734
rect 43916 23526 43944 24160
rect 44180 24142 44232 24148
rect 44560 24138 44588 24346
rect 43996 24132 44048 24138
rect 43996 24074 44048 24080
rect 44548 24132 44600 24138
rect 44548 24074 44600 24080
rect 44008 23798 44036 24074
rect 43996 23792 44048 23798
rect 43996 23734 44048 23740
rect 43904 23520 43956 23526
rect 43904 23462 43956 23468
rect 43916 23118 43944 23462
rect 44008 23186 44036 23734
rect 43996 23180 44048 23186
rect 43996 23122 44048 23128
rect 43904 23112 43956 23118
rect 43904 23054 43956 23060
rect 43536 22976 43588 22982
rect 43536 22918 43588 22924
rect 43548 22778 43576 22918
rect 43536 22772 43588 22778
rect 43536 22714 43588 22720
rect 43352 21344 43404 21350
rect 43352 21286 43404 21292
rect 43364 20466 43392 21286
rect 43444 20936 43496 20942
rect 43444 20878 43496 20884
rect 43628 20936 43680 20942
rect 43628 20878 43680 20884
rect 43352 20460 43404 20466
rect 43352 20402 43404 20408
rect 43364 19417 43392 20402
rect 43456 20398 43484 20878
rect 43444 20392 43496 20398
rect 43444 20334 43496 20340
rect 43456 19922 43484 20334
rect 43640 20262 43668 20878
rect 43996 20868 44048 20874
rect 43996 20810 44048 20816
rect 44008 20466 44036 20810
rect 43996 20460 44048 20466
rect 43996 20402 44048 20408
rect 43628 20256 43680 20262
rect 43628 20198 43680 20204
rect 43444 19916 43496 19922
rect 43444 19858 43496 19864
rect 44180 19848 44232 19854
rect 44180 19790 44232 19796
rect 44192 19514 44220 19790
rect 44180 19508 44232 19514
rect 44180 19450 44232 19456
rect 43350 19408 43406 19417
rect 43350 19343 43406 19352
rect 43996 19372 44048 19378
rect 43996 19314 44048 19320
rect 44008 18970 44036 19314
rect 43996 18964 44048 18970
rect 43996 18906 44048 18912
rect 43996 17740 44048 17746
rect 43996 17682 44048 17688
rect 43904 17264 43956 17270
rect 43904 17206 43956 17212
rect 43916 16590 43944 17206
rect 44008 17202 44036 17682
rect 44180 17672 44232 17678
rect 44180 17614 44232 17620
rect 44088 17604 44140 17610
rect 44088 17546 44140 17552
rect 44100 17270 44128 17546
rect 44088 17264 44140 17270
rect 44088 17206 44140 17212
rect 43996 17196 44048 17202
rect 43996 17138 44048 17144
rect 44008 16726 44036 17138
rect 44192 16998 44220 17614
rect 44272 17332 44324 17338
rect 44272 17274 44324 17280
rect 44180 16992 44232 16998
rect 44180 16934 44232 16940
rect 43996 16720 44048 16726
rect 43996 16662 44048 16668
rect 43260 16584 43312 16590
rect 43260 16526 43312 16532
rect 43904 16584 43956 16590
rect 43904 16526 43956 16532
rect 43272 16114 43300 16526
rect 43812 16448 43864 16454
rect 43812 16390 43864 16396
rect 43824 16182 43852 16390
rect 43812 16176 43864 16182
rect 43812 16118 43864 16124
rect 43260 16108 43312 16114
rect 43260 16050 43312 16056
rect 43272 15094 43300 16050
rect 43824 15706 43852 16118
rect 43916 16114 43944 16526
rect 43996 16244 44048 16250
rect 43996 16186 44048 16192
rect 43904 16108 43956 16114
rect 43904 16050 43956 16056
rect 43812 15700 43864 15706
rect 43812 15642 43864 15648
rect 43916 15434 43944 16050
rect 43904 15428 43956 15434
rect 43904 15370 43956 15376
rect 43260 15088 43312 15094
rect 43260 15030 43312 15036
rect 43904 14544 43956 14550
rect 43904 14486 43956 14492
rect 43916 13938 43944 14486
rect 44008 14414 44036 16186
rect 44088 16040 44140 16046
rect 44284 15994 44312 17274
rect 44456 16516 44508 16522
rect 44456 16458 44508 16464
rect 44468 16046 44496 16458
rect 44140 15988 44312 15994
rect 44088 15982 44312 15988
rect 44456 16040 44508 16046
rect 44456 15982 44508 15988
rect 44100 15966 44312 15982
rect 44180 15904 44232 15910
rect 44180 15846 44232 15852
rect 44088 15088 44140 15094
rect 44088 15030 44140 15036
rect 44100 14482 44128 15030
rect 44192 15026 44220 15846
rect 44180 15020 44232 15026
rect 44180 14962 44232 14968
rect 44284 14482 44312 15966
rect 44468 15434 44496 15982
rect 44456 15428 44508 15434
rect 44456 15370 44508 15376
rect 44364 15020 44416 15026
rect 44364 14962 44416 14968
rect 44376 14822 44404 14962
rect 44364 14816 44416 14822
rect 44364 14758 44416 14764
rect 44088 14476 44140 14482
rect 44088 14418 44140 14424
rect 44272 14476 44324 14482
rect 44272 14418 44324 14424
rect 43996 14408 44048 14414
rect 43996 14350 44048 14356
rect 44008 13938 44036 14350
rect 43904 13932 43956 13938
rect 43904 13874 43956 13880
rect 43996 13932 44048 13938
rect 43996 13874 44048 13880
rect 44100 13870 44128 14418
rect 44376 14385 44404 14758
rect 44362 14376 44418 14385
rect 44362 14311 44418 14320
rect 44088 13864 44140 13870
rect 44088 13806 44140 13812
rect 43352 13184 43404 13190
rect 43352 13126 43404 13132
rect 43364 12986 43392 13126
rect 43352 12980 43404 12986
rect 43352 12922 43404 12928
rect 43180 12406 43300 12434
rect 43168 12096 43220 12102
rect 43168 12038 43220 12044
rect 43076 11824 43128 11830
rect 43076 11766 43128 11772
rect 43088 11150 43116 11766
rect 43180 11762 43208 12038
rect 43168 11756 43220 11762
rect 43168 11698 43220 11704
rect 43180 11286 43208 11698
rect 43168 11280 43220 11286
rect 43168 11222 43220 11228
rect 42340 11144 42392 11150
rect 42340 11086 42392 11092
rect 43076 11144 43128 11150
rect 43076 11086 43128 11092
rect 41880 10192 41932 10198
rect 41880 10134 41932 10140
rect 41788 10056 41840 10062
rect 41788 9998 41840 10004
rect 41800 9926 41828 9998
rect 41696 9920 41748 9926
rect 41696 9862 41748 9868
rect 41788 9920 41840 9926
rect 41788 9862 41840 9868
rect 41708 9586 41736 9862
rect 41696 9580 41748 9586
rect 41696 9522 41748 9528
rect 41892 7886 41920 10134
rect 42352 8498 42380 11086
rect 43168 10804 43220 10810
rect 43168 10746 43220 10752
rect 43180 10130 43208 10746
rect 43168 10124 43220 10130
rect 43168 10066 43220 10072
rect 42892 9988 42944 9994
rect 42892 9930 42944 9936
rect 42708 9920 42760 9926
rect 42708 9862 42760 9868
rect 42720 9654 42748 9862
rect 42708 9648 42760 9654
rect 42708 9590 42760 9596
rect 42904 9382 42932 9930
rect 43180 9586 43208 10066
rect 43168 9580 43220 9586
rect 43168 9522 43220 9528
rect 42524 9376 42576 9382
rect 42524 9318 42576 9324
rect 42892 9376 42944 9382
rect 42892 9318 42944 9324
rect 42340 8492 42392 8498
rect 42340 8434 42392 8440
rect 42352 7886 42380 8434
rect 42536 7886 42564 9318
rect 43180 9178 43208 9522
rect 43168 9172 43220 9178
rect 43168 9114 43220 9120
rect 41880 7880 41932 7886
rect 41880 7822 41932 7828
rect 42340 7880 42392 7886
rect 42340 7822 42392 7828
rect 42524 7880 42576 7886
rect 42524 7822 42576 7828
rect 42536 7478 42564 7822
rect 42616 7744 42668 7750
rect 42616 7686 42668 7692
rect 42524 7472 42576 7478
rect 42524 7414 42576 7420
rect 42628 7410 42656 7686
rect 42616 7404 42668 7410
rect 42616 7346 42668 7352
rect 42248 4208 42300 4214
rect 42248 4150 42300 4156
rect 42064 4004 42116 4010
rect 42064 3946 42116 3952
rect 42076 3670 42104 3946
rect 41604 3664 41656 3670
rect 41604 3606 41656 3612
rect 42064 3664 42116 3670
rect 42064 3606 42116 3612
rect 40040 3528 40092 3534
rect 40040 3470 40092 3476
rect 40868 3528 40920 3534
rect 40868 3470 40920 3476
rect 41052 3528 41104 3534
rect 41052 3470 41104 3476
rect 37740 3392 37792 3398
rect 37740 3334 37792 3340
rect 40052 3058 40080 3470
rect 40224 3392 40276 3398
rect 40224 3334 40276 3340
rect 40868 3392 40920 3398
rect 40868 3334 40920 3340
rect 41328 3392 41380 3398
rect 41328 3334 41380 3340
rect 40236 3194 40264 3334
rect 40224 3188 40276 3194
rect 40224 3130 40276 3136
rect 40040 3052 40092 3058
rect 40040 2994 40092 3000
rect 37464 2984 37516 2990
rect 37464 2926 37516 2932
rect 39948 2916 40000 2922
rect 39948 2858 40000 2864
rect 33416 2848 33468 2854
rect 33416 2790 33468 2796
rect 33428 2446 33456 2790
rect 34934 2748 35242 2768
rect 34934 2746 34940 2748
rect 34996 2746 35020 2748
rect 35076 2746 35100 2748
rect 35156 2746 35180 2748
rect 35236 2746 35242 2748
rect 34996 2694 34998 2746
rect 35178 2694 35180 2746
rect 34934 2692 34940 2694
rect 34996 2692 35020 2694
rect 35076 2692 35100 2694
rect 35156 2692 35180 2694
rect 35236 2692 35242 2694
rect 34934 2672 35242 2692
rect 39960 2650 39988 2858
rect 40132 2848 40184 2854
rect 40132 2790 40184 2796
rect 39948 2644 40000 2650
rect 39948 2586 40000 2592
rect 40144 2446 40172 2790
rect 40236 2446 40264 3130
rect 40880 3058 40908 3334
rect 41340 3126 41368 3334
rect 41328 3120 41380 3126
rect 41328 3062 41380 3068
rect 40868 3052 40920 3058
rect 40868 2994 40920 3000
rect 41616 2446 41644 3606
rect 42260 3466 42288 4150
rect 43272 3534 43300 12406
rect 43812 12164 43864 12170
rect 43812 12106 43864 12112
rect 43720 12096 43772 12102
rect 43720 12038 43772 12044
rect 43732 11830 43760 12038
rect 43720 11824 43772 11830
rect 43720 11766 43772 11772
rect 43824 11762 43852 12106
rect 43812 11756 43864 11762
rect 43812 11698 43864 11704
rect 43824 11082 43852 11698
rect 43812 11076 43864 11082
rect 43812 11018 43864 11024
rect 44180 9920 44232 9926
rect 44180 9862 44232 9868
rect 44192 9654 44220 9862
rect 44180 9648 44232 9654
rect 44180 9590 44232 9596
rect 43536 7540 43588 7546
rect 43536 7482 43588 7488
rect 43548 6390 43576 7482
rect 44652 6390 44680 36042
rect 45100 35692 45152 35698
rect 45100 35634 45152 35640
rect 45112 34542 45140 35634
rect 45100 34536 45152 34542
rect 45100 34478 45152 34484
rect 45112 33998 45140 34478
rect 45008 33992 45060 33998
rect 45008 33934 45060 33940
rect 45100 33992 45152 33998
rect 45152 33952 45232 33980
rect 45100 33934 45152 33940
rect 44732 33516 44784 33522
rect 44732 33458 44784 33464
rect 44916 33516 44968 33522
rect 44916 33458 44968 33464
rect 44744 22094 44772 33458
rect 44928 32910 44956 33458
rect 45020 33454 45048 33934
rect 45204 33522 45232 33952
rect 45836 33856 45888 33862
rect 45836 33798 45888 33804
rect 45100 33516 45152 33522
rect 45100 33458 45152 33464
rect 45192 33516 45244 33522
rect 45192 33458 45244 33464
rect 45008 33448 45060 33454
rect 45008 33390 45060 33396
rect 44916 32904 44968 32910
rect 44916 32846 44968 32852
rect 44928 32434 44956 32846
rect 44916 32428 44968 32434
rect 44916 32370 44968 32376
rect 45112 32366 45140 33458
rect 45560 33380 45612 33386
rect 45560 33322 45612 33328
rect 45192 32904 45244 32910
rect 45192 32846 45244 32852
rect 45100 32360 45152 32366
rect 45100 32302 45152 32308
rect 45204 32230 45232 32846
rect 45192 32224 45244 32230
rect 45192 32166 45244 32172
rect 45008 32020 45060 32026
rect 45008 31962 45060 31968
rect 44824 31204 44876 31210
rect 44824 31146 44876 31152
rect 44836 30666 44864 31146
rect 45020 30802 45048 31962
rect 45100 31816 45152 31822
rect 45100 31758 45152 31764
rect 45112 31278 45140 31758
rect 45100 31272 45152 31278
rect 45100 31214 45152 31220
rect 45204 30938 45232 32166
rect 45572 31822 45600 33322
rect 45848 32910 45876 33798
rect 45836 32904 45888 32910
rect 45836 32846 45888 32852
rect 46204 32904 46256 32910
rect 46204 32846 46256 32852
rect 45652 32768 45704 32774
rect 45652 32710 45704 32716
rect 45664 32434 45692 32710
rect 46216 32570 46244 32846
rect 46204 32564 46256 32570
rect 46204 32506 46256 32512
rect 45652 32428 45704 32434
rect 45652 32370 45704 32376
rect 45664 31890 45692 32370
rect 45652 31884 45704 31890
rect 45652 31826 45704 31832
rect 45560 31816 45612 31822
rect 45560 31758 45612 31764
rect 45376 31748 45428 31754
rect 45376 31690 45428 31696
rect 45388 31346 45416 31690
rect 45376 31340 45428 31346
rect 45376 31282 45428 31288
rect 45284 31272 45336 31278
rect 45284 31214 45336 31220
rect 45572 31226 45600 31758
rect 45664 31346 45692 31826
rect 45652 31340 45704 31346
rect 45652 31282 45704 31288
rect 45296 30938 45324 31214
rect 45572 31210 45692 31226
rect 45572 31204 45704 31210
rect 45572 31198 45652 31204
rect 45652 31146 45704 31152
rect 45192 30932 45244 30938
rect 45192 30874 45244 30880
rect 45284 30932 45336 30938
rect 45284 30874 45336 30880
rect 45008 30796 45060 30802
rect 45008 30738 45060 30744
rect 44824 30660 44876 30666
rect 44824 30602 44876 30608
rect 44836 30394 44864 30602
rect 45020 30410 45048 30738
rect 44824 30388 44876 30394
rect 45020 30382 45140 30410
rect 44824 30330 44876 30336
rect 45112 30258 45140 30382
rect 45008 30252 45060 30258
rect 45008 30194 45060 30200
rect 45100 30252 45152 30258
rect 45100 30194 45152 30200
rect 45020 29646 45048 30194
rect 45204 30054 45232 30874
rect 45376 30728 45428 30734
rect 45376 30670 45428 30676
rect 45388 30054 45416 30670
rect 45468 30592 45520 30598
rect 45468 30534 45520 30540
rect 45192 30048 45244 30054
rect 45192 29990 45244 29996
rect 45376 30048 45428 30054
rect 45376 29990 45428 29996
rect 45480 29850 45508 30534
rect 45468 29844 45520 29850
rect 45468 29786 45520 29792
rect 45008 29640 45060 29646
rect 45008 29582 45060 29588
rect 45020 29238 45048 29582
rect 45008 29232 45060 29238
rect 45008 29174 45060 29180
rect 45468 29164 45520 29170
rect 45468 29106 45520 29112
rect 45192 29096 45244 29102
rect 45192 29038 45244 29044
rect 45204 28626 45232 29038
rect 45192 28620 45244 28626
rect 45192 28562 45244 28568
rect 45480 28558 45508 29106
rect 45468 28552 45520 28558
rect 45468 28494 45520 28500
rect 44916 28076 44968 28082
rect 44916 28018 44968 28024
rect 44928 27470 44956 28018
rect 45008 28008 45060 28014
rect 45008 27950 45060 27956
rect 44916 27464 44968 27470
rect 44916 27406 44968 27412
rect 44928 27130 44956 27406
rect 45020 27130 45048 27950
rect 45100 27940 45152 27946
rect 45100 27882 45152 27888
rect 45112 27538 45140 27882
rect 45480 27674 45508 28494
rect 45468 27668 45520 27674
rect 45468 27610 45520 27616
rect 45100 27532 45152 27538
rect 45100 27474 45152 27480
rect 44916 27124 44968 27130
rect 44916 27066 44968 27072
rect 45008 27124 45060 27130
rect 45008 27066 45060 27072
rect 45112 26314 45140 27474
rect 45100 26308 45152 26314
rect 45100 26250 45152 26256
rect 45744 25288 45796 25294
rect 45928 25288 45980 25294
rect 45744 25230 45796 25236
rect 45848 25248 45928 25276
rect 45756 24818 45784 25230
rect 45848 24818 45876 25248
rect 45928 25230 45980 25236
rect 46112 25288 46164 25294
rect 46112 25230 46164 25236
rect 46296 25288 46348 25294
rect 46296 25230 46348 25236
rect 45376 24812 45428 24818
rect 45376 24754 45428 24760
rect 45744 24812 45796 24818
rect 45744 24754 45796 24760
rect 45836 24812 45888 24818
rect 45836 24754 45888 24760
rect 45100 24744 45152 24750
rect 45100 24686 45152 24692
rect 45112 24274 45140 24686
rect 45100 24268 45152 24274
rect 45100 24210 45152 24216
rect 45388 24206 45416 24754
rect 45652 24744 45704 24750
rect 45652 24686 45704 24692
rect 45664 24410 45692 24686
rect 45848 24614 45876 24754
rect 46124 24750 46152 25230
rect 46308 24818 46336 25230
rect 46296 24812 46348 24818
rect 46296 24754 46348 24760
rect 46112 24744 46164 24750
rect 46112 24686 46164 24692
rect 45836 24608 45888 24614
rect 45836 24550 45888 24556
rect 45652 24404 45704 24410
rect 45652 24346 45704 24352
rect 45376 24200 45428 24206
rect 45376 24142 45428 24148
rect 45388 23594 45416 24142
rect 45376 23588 45428 23594
rect 45376 23530 45428 23536
rect 46020 23112 46072 23118
rect 46020 23054 46072 23060
rect 46296 23112 46348 23118
rect 46296 23054 46348 23060
rect 46032 22778 46060 23054
rect 46112 22976 46164 22982
rect 46112 22918 46164 22924
rect 46020 22772 46072 22778
rect 46020 22714 46072 22720
rect 46032 22234 46060 22714
rect 46124 22438 46152 22918
rect 46308 22710 46336 23054
rect 46296 22704 46348 22710
rect 46296 22646 46348 22652
rect 46112 22432 46164 22438
rect 46112 22374 46164 22380
rect 46020 22228 46072 22234
rect 46020 22170 46072 22176
rect 44744 22066 44956 22094
rect 44732 18284 44784 18290
rect 44732 18226 44784 18232
rect 44744 17678 44772 18226
rect 44732 17672 44784 17678
rect 44732 17614 44784 17620
rect 44928 12434 44956 22066
rect 45652 22024 45704 22030
rect 45652 21966 45704 21972
rect 45008 21616 45060 21622
rect 45008 21558 45060 21564
rect 45020 20942 45048 21558
rect 45664 21554 45692 21966
rect 45836 21888 45888 21894
rect 45836 21830 45888 21836
rect 45652 21548 45704 21554
rect 45652 21490 45704 21496
rect 45664 21146 45692 21490
rect 45848 21486 45876 21830
rect 45836 21480 45888 21486
rect 45836 21422 45888 21428
rect 45652 21140 45704 21146
rect 45652 21082 45704 21088
rect 45284 21072 45336 21078
rect 45284 21014 45336 21020
rect 45296 20942 45324 21014
rect 45008 20936 45060 20942
rect 45008 20878 45060 20884
rect 45284 20936 45336 20942
rect 45284 20878 45336 20884
rect 45020 20534 45048 20878
rect 45100 20800 45152 20806
rect 45100 20742 45152 20748
rect 45008 20528 45060 20534
rect 45008 20470 45060 20476
rect 45112 20466 45140 20742
rect 45296 20466 45324 20878
rect 45100 20460 45152 20466
rect 45100 20402 45152 20408
rect 45284 20460 45336 20466
rect 45284 20402 45336 20408
rect 45112 19310 45140 20402
rect 45848 20330 45876 21422
rect 45836 20324 45888 20330
rect 45836 20266 45888 20272
rect 46020 19372 46072 19378
rect 46020 19314 46072 19320
rect 45100 19304 45152 19310
rect 45100 19246 45152 19252
rect 45112 18766 45140 19246
rect 46032 18766 46060 19314
rect 45100 18760 45152 18766
rect 45100 18702 45152 18708
rect 46020 18760 46072 18766
rect 46020 18702 46072 18708
rect 46032 18358 46060 18702
rect 46020 18352 46072 18358
rect 46020 18294 46072 18300
rect 45100 18148 45152 18154
rect 45100 18090 45152 18096
rect 45112 17882 45140 18090
rect 45100 17876 45152 17882
rect 45100 17818 45152 17824
rect 45376 17740 45428 17746
rect 45376 17682 45428 17688
rect 45388 17202 45416 17682
rect 45376 17196 45428 17202
rect 45376 17138 45428 17144
rect 45284 16992 45336 16998
rect 45284 16934 45336 16940
rect 45296 15366 45324 16934
rect 45928 16788 45980 16794
rect 45928 16730 45980 16736
rect 45940 16590 45968 16730
rect 45928 16584 45980 16590
rect 46400 16574 46428 36790
rect 46584 36786 46612 37062
rect 46768 37046 46980 37074
rect 46572 36780 46624 36786
rect 46572 36722 46624 36728
rect 46584 36106 46612 36722
rect 46572 36100 46624 36106
rect 46572 36042 46624 36048
rect 46952 34134 46980 37046
rect 46940 34128 46992 34134
rect 46940 34070 46992 34076
rect 47044 32842 47072 37266
rect 48424 37262 48452 37318
rect 47584 37256 47636 37262
rect 47584 37198 47636 37204
rect 48412 37256 48464 37262
rect 48412 37198 48464 37204
rect 47596 36922 47624 37198
rect 48228 37188 48280 37194
rect 48228 37130 48280 37136
rect 48240 36922 48268 37130
rect 47400 36916 47452 36922
rect 47400 36858 47452 36864
rect 47584 36916 47636 36922
rect 47584 36858 47636 36864
rect 48228 36916 48280 36922
rect 48228 36858 48280 36864
rect 47124 36780 47176 36786
rect 47124 36722 47176 36728
rect 47136 36174 47164 36722
rect 47412 36378 47440 36858
rect 47676 36712 47728 36718
rect 47676 36654 47728 36660
rect 47400 36372 47452 36378
rect 47400 36314 47452 36320
rect 47688 36174 47716 36654
rect 47124 36168 47176 36174
rect 47124 36110 47176 36116
rect 47676 36168 47728 36174
rect 47676 36110 47728 36116
rect 47136 35834 47164 36110
rect 47124 35828 47176 35834
rect 47124 35770 47176 35776
rect 48504 35080 48556 35086
rect 48504 35022 48556 35028
rect 48412 34944 48464 34950
rect 48412 34886 48464 34892
rect 48424 34610 48452 34886
rect 48412 34604 48464 34610
rect 48412 34546 48464 34552
rect 48516 34474 48544 35022
rect 48608 34746 48636 37402
rect 50264 37262 50292 39200
rect 48964 37256 49016 37262
rect 50252 37256 50304 37262
rect 48964 37198 49016 37204
rect 50172 37204 50252 37210
rect 50172 37198 50304 37204
rect 48976 36922 49004 37198
rect 50172 37182 50292 37198
rect 50068 37120 50120 37126
rect 50068 37062 50120 37068
rect 48964 36916 49016 36922
rect 48964 36858 49016 36864
rect 49056 36236 49108 36242
rect 49056 36178 49108 36184
rect 48964 36168 49016 36174
rect 48964 36110 49016 36116
rect 48688 35012 48740 35018
rect 48688 34954 48740 34960
rect 48596 34740 48648 34746
rect 48596 34682 48648 34688
rect 48700 34678 48728 34954
rect 48976 34746 49004 36110
rect 49068 35834 49096 36178
rect 49056 35828 49108 35834
rect 49056 35770 49108 35776
rect 49424 35692 49476 35698
rect 49424 35634 49476 35640
rect 49056 35080 49108 35086
rect 49056 35022 49108 35028
rect 48964 34740 49016 34746
rect 48964 34682 49016 34688
rect 48688 34672 48740 34678
rect 48688 34614 48740 34620
rect 48504 34468 48556 34474
rect 48504 34410 48556 34416
rect 48516 33590 48544 34410
rect 48700 34202 48728 34614
rect 48872 34536 48924 34542
rect 48872 34478 48924 34484
rect 48688 34196 48740 34202
rect 48688 34138 48740 34144
rect 48700 33998 48728 34138
rect 48688 33992 48740 33998
rect 48688 33934 48740 33940
rect 48504 33584 48556 33590
rect 48504 33526 48556 33532
rect 48884 33114 48912 34478
rect 49068 33930 49096 35022
rect 49436 34406 49464 35634
rect 49976 35624 50028 35630
rect 49976 35566 50028 35572
rect 49516 35148 49568 35154
rect 49516 35090 49568 35096
rect 49528 34542 49556 35090
rect 49988 34950 50016 35566
rect 49976 34944 50028 34950
rect 49976 34886 50028 34892
rect 49988 34610 50016 34886
rect 49976 34604 50028 34610
rect 49976 34546 50028 34552
rect 49516 34536 49568 34542
rect 49516 34478 49568 34484
rect 49424 34400 49476 34406
rect 49424 34342 49476 34348
rect 49436 34202 49464 34342
rect 49424 34196 49476 34202
rect 49424 34138 49476 34144
rect 49056 33924 49108 33930
rect 49056 33866 49108 33872
rect 48964 33516 49016 33522
rect 48964 33458 49016 33464
rect 48872 33108 48924 33114
rect 48872 33050 48924 33056
rect 48976 32910 49004 33458
rect 48780 32904 48832 32910
rect 48964 32904 49016 32910
rect 48832 32864 48912 32892
rect 48780 32846 48832 32852
rect 47032 32836 47084 32842
rect 47032 32778 47084 32784
rect 47952 32428 48004 32434
rect 47952 32370 48004 32376
rect 47964 32026 47992 32370
rect 47952 32020 48004 32026
rect 47952 31962 48004 31968
rect 48228 31884 48280 31890
rect 48228 31826 48280 31832
rect 48412 31884 48464 31890
rect 48412 31826 48464 31832
rect 48240 31278 48268 31826
rect 48320 31340 48372 31346
rect 48320 31282 48372 31288
rect 48228 31272 48280 31278
rect 48228 31214 48280 31220
rect 48240 30666 48268 31214
rect 48332 31142 48360 31282
rect 48320 31136 48372 31142
rect 48320 31078 48372 31084
rect 48332 30734 48360 31078
rect 48424 30734 48452 31826
rect 48688 31816 48740 31822
rect 48688 31758 48740 31764
rect 48596 31748 48648 31754
rect 48596 31690 48648 31696
rect 48608 31482 48636 31690
rect 48700 31482 48728 31758
rect 48596 31476 48648 31482
rect 48596 31418 48648 31424
rect 48688 31476 48740 31482
rect 48688 31418 48740 31424
rect 48608 30734 48636 31418
rect 48780 31272 48832 31278
rect 48780 31214 48832 31220
rect 48792 30734 48820 31214
rect 48320 30728 48372 30734
rect 48320 30670 48372 30676
rect 48412 30728 48464 30734
rect 48412 30670 48464 30676
rect 48596 30728 48648 30734
rect 48596 30670 48648 30676
rect 48780 30728 48832 30734
rect 48780 30670 48832 30676
rect 48228 30660 48280 30666
rect 48228 30602 48280 30608
rect 48044 30252 48096 30258
rect 48044 30194 48096 30200
rect 48056 29646 48084 30194
rect 48332 29850 48360 30670
rect 48320 29844 48372 29850
rect 48320 29786 48372 29792
rect 47676 29640 47728 29646
rect 47676 29582 47728 29588
rect 48044 29640 48096 29646
rect 48044 29582 48096 29588
rect 47688 29238 47716 29582
rect 47676 29232 47728 29238
rect 47676 29174 47728 29180
rect 47688 28490 47716 29174
rect 48056 28966 48084 29582
rect 48424 29034 48452 30670
rect 48792 30394 48820 30670
rect 48780 30388 48832 30394
rect 48780 30330 48832 30336
rect 48504 30048 48556 30054
rect 48504 29990 48556 29996
rect 48516 29646 48544 29990
rect 48504 29640 48556 29646
rect 48504 29582 48556 29588
rect 48780 29640 48832 29646
rect 48780 29582 48832 29588
rect 48792 29306 48820 29582
rect 48780 29300 48832 29306
rect 48780 29242 48832 29248
rect 48504 29096 48556 29102
rect 48504 29038 48556 29044
rect 48412 29028 48464 29034
rect 48412 28970 48464 28976
rect 48044 28960 48096 28966
rect 48044 28902 48096 28908
rect 48056 28558 48084 28902
rect 48516 28762 48544 29038
rect 48504 28756 48556 28762
rect 48504 28698 48556 28704
rect 48044 28552 48096 28558
rect 48044 28494 48096 28500
rect 48320 28552 48372 28558
rect 48320 28494 48372 28500
rect 47676 28484 47728 28490
rect 47676 28426 47728 28432
rect 46848 27872 46900 27878
rect 46848 27814 46900 27820
rect 46860 27538 46888 27814
rect 48056 27606 48084 28494
rect 48332 27674 48360 28494
rect 48320 27668 48372 27674
rect 48320 27610 48372 27616
rect 48044 27600 48096 27606
rect 48044 27542 48096 27548
rect 46848 27532 46900 27538
rect 46848 27474 46900 27480
rect 47400 27464 47452 27470
rect 47400 27406 47452 27412
rect 47412 27334 47440 27406
rect 47952 27396 48004 27402
rect 47952 27338 48004 27344
rect 47400 27328 47452 27334
rect 47400 27270 47452 27276
rect 47964 26042 47992 27338
rect 47952 26036 48004 26042
rect 47952 25978 48004 25984
rect 46848 25900 46900 25906
rect 46848 25842 46900 25848
rect 47032 25900 47084 25906
rect 47032 25842 47084 25848
rect 47584 25900 47636 25906
rect 47584 25842 47636 25848
rect 46860 25294 46888 25842
rect 46848 25288 46900 25294
rect 46848 25230 46900 25236
rect 47044 24886 47072 25842
rect 47596 25498 47624 25842
rect 47584 25492 47636 25498
rect 47584 25434 47636 25440
rect 47032 24880 47084 24886
rect 47032 24822 47084 24828
rect 47860 24200 47912 24206
rect 47860 24142 47912 24148
rect 48044 24200 48096 24206
rect 48044 24142 48096 24148
rect 47872 23866 47900 24142
rect 48056 23866 48084 24142
rect 47308 23860 47360 23866
rect 47308 23802 47360 23808
rect 47860 23860 47912 23866
rect 47860 23802 47912 23808
rect 48044 23860 48096 23866
rect 48044 23802 48096 23808
rect 47320 23118 47348 23802
rect 47584 23656 47636 23662
rect 47584 23598 47636 23604
rect 47400 23588 47452 23594
rect 47400 23530 47452 23536
rect 47412 23118 47440 23530
rect 47596 23118 47624 23598
rect 47308 23112 47360 23118
rect 47308 23054 47360 23060
rect 47400 23112 47452 23118
rect 47400 23054 47452 23060
rect 47584 23112 47636 23118
rect 47584 23054 47636 23060
rect 47596 22778 47624 23054
rect 47584 22772 47636 22778
rect 47584 22714 47636 22720
rect 46572 22432 46624 22438
rect 46572 22374 46624 22380
rect 46584 22234 46612 22374
rect 46572 22228 46624 22234
rect 46572 22170 46624 22176
rect 46480 22024 46532 22030
rect 46480 21966 46532 21972
rect 46492 21486 46520 21966
rect 48412 21548 48464 21554
rect 48412 21490 48464 21496
rect 46480 21480 46532 21486
rect 46480 21422 46532 21428
rect 48320 21480 48372 21486
rect 48320 21422 48372 21428
rect 46492 21010 46520 21422
rect 46480 21004 46532 21010
rect 46480 20946 46532 20952
rect 48332 20942 48360 21422
rect 48424 21146 48452 21490
rect 48412 21140 48464 21146
rect 48412 21082 48464 21088
rect 48320 20936 48372 20942
rect 48320 20878 48372 20884
rect 47492 20868 47544 20874
rect 47492 20810 47544 20816
rect 47504 20602 47532 20810
rect 47492 20596 47544 20602
rect 47492 20538 47544 20544
rect 48332 19922 48360 20878
rect 46940 19916 46992 19922
rect 46940 19858 46992 19864
rect 48320 19916 48372 19922
rect 48320 19858 48372 19864
rect 46952 19378 46980 19858
rect 47768 19848 47820 19854
rect 47768 19790 47820 19796
rect 47780 19378 47808 19790
rect 48780 19712 48832 19718
rect 48780 19654 48832 19660
rect 48792 19378 48820 19654
rect 46940 19372 46992 19378
rect 46940 19314 46992 19320
rect 47768 19372 47820 19378
rect 47768 19314 47820 19320
rect 48780 19372 48832 19378
rect 48780 19314 48832 19320
rect 48780 18284 48832 18290
rect 48780 18226 48832 18232
rect 48320 17604 48372 17610
rect 48320 17546 48372 17552
rect 48504 17604 48556 17610
rect 48504 17546 48556 17552
rect 48332 17338 48360 17546
rect 48320 17332 48372 17338
rect 48320 17274 48372 17280
rect 48136 17196 48188 17202
rect 48136 17138 48188 17144
rect 48148 17066 48176 17138
rect 48516 17134 48544 17546
rect 48792 17542 48820 18226
rect 48780 17536 48832 17542
rect 48780 17478 48832 17484
rect 48504 17128 48556 17134
rect 48504 17070 48556 17076
rect 48136 17060 48188 17066
rect 48136 17002 48188 17008
rect 48148 16794 48176 17002
rect 48136 16788 48188 16794
rect 48136 16730 48188 16736
rect 46400 16546 46520 16574
rect 45928 16526 45980 16532
rect 45284 15360 45336 15366
rect 45284 15302 45336 15308
rect 45376 15020 45428 15026
rect 45376 14962 45428 14968
rect 45388 14822 45416 14962
rect 45928 14952 45980 14958
rect 45928 14894 45980 14900
rect 45376 14816 45428 14822
rect 45376 14758 45428 14764
rect 45836 14816 45888 14822
rect 45836 14758 45888 14764
rect 45284 14476 45336 14482
rect 45284 14418 45336 14424
rect 45008 14272 45060 14278
rect 45008 14214 45060 14220
rect 45020 13326 45048 14214
rect 45100 14000 45152 14006
rect 45100 13942 45152 13948
rect 45112 13326 45140 13942
rect 45296 13326 45324 14418
rect 45848 14414 45876 14758
rect 45940 14414 45968 14894
rect 45836 14408 45888 14414
rect 45836 14350 45888 14356
rect 45928 14408 45980 14414
rect 45928 14350 45980 14356
rect 45008 13320 45060 13326
rect 45008 13262 45060 13268
rect 45100 13320 45152 13326
rect 45100 13262 45152 13268
rect 45284 13320 45336 13326
rect 45284 13262 45336 13268
rect 45020 12850 45048 13262
rect 45112 12918 45140 13262
rect 45100 12912 45152 12918
rect 45100 12854 45152 12860
rect 45296 12850 45324 13262
rect 45468 13184 45520 13190
rect 45468 13126 45520 13132
rect 45008 12844 45060 12850
rect 45008 12786 45060 12792
rect 45284 12844 45336 12850
rect 45284 12786 45336 12792
rect 44928 12406 45140 12434
rect 44916 11688 44968 11694
rect 44916 11630 44968 11636
rect 44928 11354 44956 11630
rect 44916 11348 44968 11354
rect 44916 11290 44968 11296
rect 45008 8356 45060 8362
rect 45008 8298 45060 8304
rect 45020 7410 45048 8298
rect 45008 7404 45060 7410
rect 45008 7346 45060 7352
rect 45020 6730 45048 7346
rect 45008 6724 45060 6730
rect 45008 6666 45060 6672
rect 43536 6384 43588 6390
rect 43456 6332 43536 6338
rect 43456 6326 43588 6332
rect 44640 6384 44692 6390
rect 44640 6326 44692 6332
rect 43456 6310 43576 6326
rect 43456 5778 43484 6310
rect 43536 6112 43588 6118
rect 43536 6054 43588 6060
rect 44456 6112 44508 6118
rect 44456 6054 44508 6060
rect 43444 5772 43496 5778
rect 43444 5714 43496 5720
rect 43548 5710 43576 6054
rect 43536 5704 43588 5710
rect 43536 5646 43588 5652
rect 44180 5568 44232 5574
rect 44180 5510 44232 5516
rect 44192 5234 44220 5510
rect 44468 5234 44496 6054
rect 44180 5228 44232 5234
rect 44180 5170 44232 5176
rect 44272 5228 44324 5234
rect 44272 5170 44324 5176
rect 44456 5228 44508 5234
rect 44456 5170 44508 5176
rect 43812 5024 43864 5030
rect 43812 4966 43864 4972
rect 43076 3528 43128 3534
rect 43076 3470 43128 3476
rect 43260 3528 43312 3534
rect 43260 3470 43312 3476
rect 42248 3460 42300 3466
rect 42248 3402 42300 3408
rect 42432 3460 42484 3466
rect 42432 3402 42484 3408
rect 42616 3460 42668 3466
rect 42616 3402 42668 3408
rect 41696 3188 41748 3194
rect 41696 3130 41748 3136
rect 41708 2990 41736 3130
rect 41696 2984 41748 2990
rect 41696 2926 41748 2932
rect 42260 2854 42288 3402
rect 42444 3194 42472 3402
rect 42432 3188 42484 3194
rect 42432 3130 42484 3136
rect 42628 3126 42656 3402
rect 43088 3126 43116 3470
rect 43168 3392 43220 3398
rect 43168 3334 43220 3340
rect 43352 3392 43404 3398
rect 43352 3334 43404 3340
rect 43180 3194 43208 3334
rect 43168 3188 43220 3194
rect 43168 3130 43220 3136
rect 42616 3120 42668 3126
rect 42616 3062 42668 3068
rect 43076 3120 43128 3126
rect 43076 3062 43128 3068
rect 42248 2848 42300 2854
rect 42248 2790 42300 2796
rect 43364 2446 43392 3334
rect 43444 3052 43496 3058
rect 43444 2994 43496 3000
rect 33232 2440 33284 2446
rect 33232 2382 33284 2388
rect 33416 2440 33468 2446
rect 33416 2382 33468 2388
rect 36084 2440 36136 2446
rect 36084 2382 36136 2388
rect 40132 2440 40184 2446
rect 40132 2382 40184 2388
rect 40224 2440 40276 2446
rect 40224 2382 40276 2388
rect 41604 2440 41656 2446
rect 41604 2382 41656 2388
rect 43352 2440 43404 2446
rect 43352 2382 43404 2388
rect 32680 2304 32732 2310
rect 32680 2246 32732 2252
rect 34152 2304 34204 2310
rect 34152 2246 34204 2252
rect 34164 800 34192 2246
rect 36096 800 36124 2382
rect 42708 2372 42760 2378
rect 42708 2314 42760 2320
rect 37556 2304 37608 2310
rect 37556 2246 37608 2252
rect 38016 2304 38068 2310
rect 40040 2304 40092 2310
rect 38016 2246 38068 2252
rect 39960 2264 40040 2292
rect 37568 2106 37596 2246
rect 37556 2100 37608 2106
rect 37556 2042 37608 2048
rect 38028 800 38056 2246
rect 39960 800 39988 2264
rect 40040 2246 40092 2252
rect 41880 2304 41932 2310
rect 41880 2246 41932 2252
rect 41892 800 41920 2246
rect 42720 1970 42748 2314
rect 43352 2304 43404 2310
rect 43456 2292 43484 2994
rect 43824 2990 43852 4966
rect 44284 4690 44312 5170
rect 44364 5160 44416 5166
rect 44364 5102 44416 5108
rect 44376 4826 44404 5102
rect 44364 4820 44416 4826
rect 44364 4762 44416 4768
rect 44272 4684 44324 4690
rect 44272 4626 44324 4632
rect 44376 4554 44404 4762
rect 44364 4548 44416 4554
rect 44364 4490 44416 4496
rect 45112 3126 45140 12406
rect 45376 12164 45428 12170
rect 45376 12106 45428 12112
rect 45388 11898 45416 12106
rect 45376 11892 45428 11898
rect 45376 11834 45428 11840
rect 45388 11082 45416 11834
rect 45480 11762 45508 13126
rect 46112 12776 46164 12782
rect 46112 12718 46164 12724
rect 45744 12232 45796 12238
rect 45744 12174 45796 12180
rect 45468 11756 45520 11762
rect 45468 11698 45520 11704
rect 45756 11150 45784 12174
rect 45836 12096 45888 12102
rect 45836 12038 45888 12044
rect 45848 11354 45876 12038
rect 46124 11762 46152 12718
rect 46112 11756 46164 11762
rect 46112 11698 46164 11704
rect 45928 11688 45980 11694
rect 45928 11630 45980 11636
rect 45836 11348 45888 11354
rect 45836 11290 45888 11296
rect 45940 11286 45968 11630
rect 45928 11280 45980 11286
rect 45928 11222 45980 11228
rect 45744 11144 45796 11150
rect 45744 11086 45796 11092
rect 45376 11076 45428 11082
rect 45376 11018 45428 11024
rect 45560 10124 45612 10130
rect 45560 10066 45612 10072
rect 45572 9586 45600 10066
rect 45560 9580 45612 9586
rect 45560 9522 45612 9528
rect 45836 9580 45888 9586
rect 45836 9522 45888 9528
rect 46020 9580 46072 9586
rect 46020 9522 46072 9528
rect 45572 9110 45600 9522
rect 45560 9104 45612 9110
rect 45560 9046 45612 9052
rect 45848 9042 45876 9522
rect 45928 9376 45980 9382
rect 45928 9318 45980 9324
rect 45836 9036 45888 9042
rect 45836 8978 45888 8984
rect 45848 8022 45876 8978
rect 45940 8430 45968 9318
rect 46032 9110 46060 9522
rect 46020 9104 46072 9110
rect 46020 9046 46072 9052
rect 46020 8492 46072 8498
rect 46020 8434 46072 8440
rect 45928 8424 45980 8430
rect 45928 8366 45980 8372
rect 45836 8016 45888 8022
rect 45836 7958 45888 7964
rect 45940 7886 45968 8366
rect 46032 7886 46060 8434
rect 45560 7880 45612 7886
rect 45560 7822 45612 7828
rect 45928 7880 45980 7886
rect 45928 7822 45980 7828
rect 46020 7880 46072 7886
rect 46020 7822 46072 7828
rect 45192 7744 45244 7750
rect 45192 7686 45244 7692
rect 45204 7410 45232 7686
rect 45192 7404 45244 7410
rect 45192 7346 45244 7352
rect 45204 6866 45232 7346
rect 45468 7336 45520 7342
rect 45468 7278 45520 7284
rect 45480 6866 45508 7278
rect 45572 7002 45600 7822
rect 46032 7546 46060 7822
rect 46020 7540 46072 7546
rect 46020 7482 46072 7488
rect 45560 6996 45612 7002
rect 45560 6938 45612 6944
rect 45192 6860 45244 6866
rect 45192 6802 45244 6808
rect 45468 6860 45520 6866
rect 45468 6802 45520 6808
rect 45192 5228 45244 5234
rect 45192 5170 45244 5176
rect 45204 4826 45232 5170
rect 45560 5092 45612 5098
rect 45560 5034 45612 5040
rect 45192 4820 45244 4826
rect 45192 4762 45244 4768
rect 45572 4622 45600 5034
rect 46296 4684 46348 4690
rect 46296 4626 46348 4632
rect 46388 4684 46440 4690
rect 46388 4626 46440 4632
rect 45560 4616 45612 4622
rect 45560 4558 45612 4564
rect 46204 4548 46256 4554
rect 46204 4490 46256 4496
rect 46216 4146 46244 4490
rect 46308 4214 46336 4626
rect 46296 4208 46348 4214
rect 46296 4150 46348 4156
rect 46204 4140 46256 4146
rect 46204 4082 46256 4088
rect 46112 4004 46164 4010
rect 46112 3946 46164 3952
rect 45192 3936 45244 3942
rect 45192 3878 45244 3884
rect 45100 3120 45152 3126
rect 45100 3062 45152 3068
rect 45204 3058 45232 3878
rect 46124 3534 46152 3946
rect 46308 3602 46336 4150
rect 46400 4078 46428 4626
rect 46388 4072 46440 4078
rect 46388 4014 46440 4020
rect 46296 3596 46348 3602
rect 46296 3538 46348 3544
rect 46112 3528 46164 3534
rect 46112 3470 46164 3476
rect 45192 3052 45244 3058
rect 45192 2994 45244 3000
rect 43812 2984 43864 2990
rect 43812 2926 43864 2932
rect 46112 2644 46164 2650
rect 46112 2586 46164 2592
rect 46124 2446 46152 2586
rect 46112 2440 46164 2446
rect 46112 2382 46164 2388
rect 43404 2264 43484 2292
rect 43812 2304 43864 2310
rect 43352 2246 43404 2252
rect 43812 2246 43864 2252
rect 45744 2304 45796 2310
rect 45744 2246 45796 2252
rect 42708 1964 42760 1970
rect 42708 1906 42760 1912
rect 43364 1834 43392 2246
rect 43352 1828 43404 1834
rect 43352 1770 43404 1776
rect 43824 800 43852 2246
rect 45756 800 45784 2246
rect 46492 2038 46520 16546
rect 48688 15972 48740 15978
rect 48688 15914 48740 15920
rect 47308 15904 47360 15910
rect 47308 15846 47360 15852
rect 47320 15570 47348 15846
rect 47308 15564 47360 15570
rect 47308 15506 47360 15512
rect 46848 15496 46900 15502
rect 46848 15438 46900 15444
rect 46860 14822 46888 15438
rect 48700 15366 48728 15914
rect 48688 15360 48740 15366
rect 48688 15302 48740 15308
rect 48700 15026 48728 15302
rect 48688 15020 48740 15026
rect 48688 14962 48740 14968
rect 48780 15020 48832 15026
rect 48780 14962 48832 14968
rect 48792 14890 48820 14962
rect 48780 14884 48832 14890
rect 48780 14826 48832 14832
rect 46848 14816 46900 14822
rect 46848 14758 46900 14764
rect 46756 13388 46808 13394
rect 46756 13330 46808 13336
rect 46662 13288 46718 13297
rect 46662 13223 46718 13232
rect 46676 11354 46704 13223
rect 46768 12850 46796 13330
rect 46860 12850 46888 14758
rect 48792 14346 48820 14826
rect 48780 14340 48832 14346
rect 48780 14282 48832 14288
rect 46940 14272 46992 14278
rect 46940 14214 46992 14220
rect 46952 13326 46980 14214
rect 46940 13320 46992 13326
rect 46940 13262 46992 13268
rect 48320 13320 48372 13326
rect 48320 13262 48372 13268
rect 47952 13252 48004 13258
rect 47952 13194 48004 13200
rect 47964 12850 47992 13194
rect 48332 12986 48360 13262
rect 48320 12980 48372 12986
rect 48320 12922 48372 12928
rect 46756 12844 46808 12850
rect 46756 12786 46808 12792
rect 46848 12844 46900 12850
rect 46848 12786 46900 12792
rect 47952 12844 48004 12850
rect 47952 12786 48004 12792
rect 48596 12232 48648 12238
rect 48596 12174 48648 12180
rect 48608 11694 48636 12174
rect 48596 11688 48648 11694
rect 48596 11630 48648 11636
rect 47952 11552 48004 11558
rect 47952 11494 48004 11500
rect 46664 11348 46716 11354
rect 46664 11290 46716 11296
rect 47676 11348 47728 11354
rect 47676 11290 47728 11296
rect 47688 11218 47716 11290
rect 47676 11212 47728 11218
rect 47676 11154 47728 11160
rect 47688 10810 47716 11154
rect 47676 10804 47728 10810
rect 47676 10746 47728 10752
rect 47766 10160 47822 10169
rect 47766 10095 47822 10104
rect 47780 10062 47808 10095
rect 47768 10056 47820 10062
rect 47768 9998 47820 10004
rect 47964 6866 47992 11494
rect 48608 11286 48636 11630
rect 48596 11280 48648 11286
rect 48596 11222 48648 11228
rect 48596 11144 48648 11150
rect 48424 11092 48596 11098
rect 48424 11086 48648 11092
rect 48424 11070 48636 11086
rect 48688 11076 48740 11082
rect 48424 11014 48452 11070
rect 48688 11018 48740 11024
rect 48412 11008 48464 11014
rect 48412 10950 48464 10956
rect 48412 10056 48464 10062
rect 48412 9998 48464 10004
rect 48320 8628 48372 8634
rect 48320 8570 48372 8576
rect 48332 8362 48360 8570
rect 48424 8362 48452 9998
rect 48700 8974 48728 11018
rect 48688 8968 48740 8974
rect 48688 8910 48740 8916
rect 48688 8492 48740 8498
rect 48688 8434 48740 8440
rect 48320 8356 48372 8362
rect 48320 8298 48372 8304
rect 48412 8356 48464 8362
rect 48412 8298 48464 8304
rect 48332 7954 48360 8298
rect 48320 7948 48372 7954
rect 48320 7890 48372 7896
rect 48700 7886 48728 8434
rect 48688 7880 48740 7886
rect 48688 7822 48740 7828
rect 48700 7002 48728 7822
rect 48688 6996 48740 7002
rect 48688 6938 48740 6944
rect 47676 6860 47728 6866
rect 47676 6802 47728 6808
rect 47952 6860 48004 6866
rect 47952 6802 48004 6808
rect 47688 6322 47716 6802
rect 47964 6322 47992 6802
rect 47676 6316 47728 6322
rect 47676 6258 47728 6264
rect 47952 6316 48004 6322
rect 47952 6258 48004 6264
rect 48884 2774 48912 32864
rect 48964 32846 49016 32852
rect 48976 32570 49004 32846
rect 48964 32564 49016 32570
rect 48964 32506 49016 32512
rect 49068 32026 49096 33866
rect 49332 33516 49384 33522
rect 49332 33458 49384 33464
rect 49344 32978 49372 33458
rect 49332 32972 49384 32978
rect 49332 32914 49384 32920
rect 49056 32020 49108 32026
rect 49056 31962 49108 31968
rect 49528 30122 49556 34478
rect 49792 32428 49844 32434
rect 49792 32370 49844 32376
rect 49804 31482 49832 32370
rect 49792 31476 49844 31482
rect 49792 31418 49844 31424
rect 50080 31210 50108 37062
rect 50172 36922 50200 37182
rect 52196 37126 52224 39200
rect 52552 37256 52604 37262
rect 52552 37198 52604 37204
rect 50712 37120 50764 37126
rect 50712 37062 50764 37068
rect 52184 37120 52236 37126
rect 52184 37062 52236 37068
rect 50294 37020 50602 37040
rect 50294 37018 50300 37020
rect 50356 37018 50380 37020
rect 50436 37018 50460 37020
rect 50516 37018 50540 37020
rect 50596 37018 50602 37020
rect 50356 36966 50358 37018
rect 50538 36966 50540 37018
rect 50294 36964 50300 36966
rect 50356 36964 50380 36966
rect 50436 36964 50460 36966
rect 50516 36964 50540 36966
rect 50596 36964 50602 36966
rect 50294 36944 50602 36964
rect 50160 36916 50212 36922
rect 50160 36858 50212 36864
rect 50294 35932 50602 35952
rect 50294 35930 50300 35932
rect 50356 35930 50380 35932
rect 50436 35930 50460 35932
rect 50516 35930 50540 35932
rect 50596 35930 50602 35932
rect 50356 35878 50358 35930
rect 50538 35878 50540 35930
rect 50294 35876 50300 35878
rect 50356 35876 50380 35878
rect 50436 35876 50460 35878
rect 50516 35876 50540 35878
rect 50596 35876 50602 35878
rect 50294 35856 50602 35876
rect 50724 35766 50752 37062
rect 50712 35760 50764 35766
rect 50712 35702 50764 35708
rect 52184 35148 52236 35154
rect 52184 35090 52236 35096
rect 50294 34844 50602 34864
rect 50294 34842 50300 34844
rect 50356 34842 50380 34844
rect 50436 34842 50460 34844
rect 50516 34842 50540 34844
rect 50596 34842 50602 34844
rect 50356 34790 50358 34842
rect 50538 34790 50540 34842
rect 50294 34788 50300 34790
rect 50356 34788 50380 34790
rect 50436 34788 50460 34790
rect 50516 34788 50540 34790
rect 50596 34788 50602 34790
rect 50294 34768 50602 34788
rect 52196 34746 52224 35090
rect 52184 34740 52236 34746
rect 52184 34682 52236 34688
rect 52460 34672 52512 34678
rect 52460 34614 52512 34620
rect 52184 34468 52236 34474
rect 52184 34410 52236 34416
rect 52196 33998 52224 34410
rect 52472 34066 52500 34614
rect 52460 34060 52512 34066
rect 52460 34002 52512 34008
rect 51264 33992 51316 33998
rect 51264 33934 51316 33940
rect 52184 33992 52236 33998
rect 52184 33934 52236 33940
rect 50294 33756 50602 33776
rect 50294 33754 50300 33756
rect 50356 33754 50380 33756
rect 50436 33754 50460 33756
rect 50516 33754 50540 33756
rect 50596 33754 50602 33756
rect 50356 33702 50358 33754
rect 50538 33702 50540 33754
rect 50294 33700 50300 33702
rect 50356 33700 50380 33702
rect 50436 33700 50460 33702
rect 50516 33700 50540 33702
rect 50596 33700 50602 33702
rect 50294 33680 50602 33700
rect 51276 33522 51304 33934
rect 52184 33856 52236 33862
rect 52184 33798 52236 33804
rect 51264 33516 51316 33522
rect 51264 33458 51316 33464
rect 50294 32668 50602 32688
rect 50294 32666 50300 32668
rect 50356 32666 50380 32668
rect 50436 32666 50460 32668
rect 50516 32666 50540 32668
rect 50596 32666 50602 32668
rect 50356 32614 50358 32666
rect 50538 32614 50540 32666
rect 50294 32612 50300 32614
rect 50356 32612 50380 32614
rect 50436 32612 50460 32614
rect 50516 32612 50540 32614
rect 50596 32612 50602 32614
rect 50294 32592 50602 32612
rect 50294 31580 50602 31600
rect 50294 31578 50300 31580
rect 50356 31578 50380 31580
rect 50436 31578 50460 31580
rect 50516 31578 50540 31580
rect 50596 31578 50602 31580
rect 50356 31526 50358 31578
rect 50538 31526 50540 31578
rect 50294 31524 50300 31526
rect 50356 31524 50380 31526
rect 50436 31524 50460 31526
rect 50516 31524 50540 31526
rect 50596 31524 50602 31526
rect 50294 31504 50602 31524
rect 49976 31204 50028 31210
rect 49976 31146 50028 31152
rect 50068 31204 50120 31210
rect 50068 31146 50120 31152
rect 49988 30734 50016 31146
rect 49976 30728 50028 30734
rect 49976 30670 50028 30676
rect 50896 30728 50948 30734
rect 50896 30670 50948 30676
rect 50294 30492 50602 30512
rect 50294 30490 50300 30492
rect 50356 30490 50380 30492
rect 50436 30490 50460 30492
rect 50516 30490 50540 30492
rect 50596 30490 50602 30492
rect 50356 30438 50358 30490
rect 50538 30438 50540 30490
rect 50294 30436 50300 30438
rect 50356 30436 50380 30438
rect 50436 30436 50460 30438
rect 50516 30436 50540 30438
rect 50596 30436 50602 30438
rect 50294 30416 50602 30436
rect 49516 30116 49568 30122
rect 49516 30058 49568 30064
rect 50294 29404 50602 29424
rect 50294 29402 50300 29404
rect 50356 29402 50380 29404
rect 50436 29402 50460 29404
rect 50516 29402 50540 29404
rect 50596 29402 50602 29404
rect 50356 29350 50358 29402
rect 50538 29350 50540 29402
rect 50294 29348 50300 29350
rect 50356 29348 50380 29350
rect 50436 29348 50460 29350
rect 50516 29348 50540 29350
rect 50596 29348 50602 29350
rect 50294 29328 50602 29348
rect 49608 29300 49660 29306
rect 49608 29242 49660 29248
rect 49148 29164 49200 29170
rect 49148 29106 49200 29112
rect 49160 28540 49188 29106
rect 49620 28558 49648 29242
rect 50908 29170 50936 30670
rect 51080 30660 51132 30666
rect 51080 30602 51132 30608
rect 51092 29238 51120 30602
rect 51080 29232 51132 29238
rect 51080 29174 51132 29180
rect 50896 29164 50948 29170
rect 50896 29106 50948 29112
rect 51276 28762 51304 33458
rect 52196 33318 52224 33798
rect 52472 33590 52500 34002
rect 52460 33584 52512 33590
rect 52460 33526 52512 33532
rect 52184 33312 52236 33318
rect 52184 33254 52236 33260
rect 52196 31754 52224 33254
rect 51920 31726 52224 31754
rect 52276 31748 52328 31754
rect 51356 30864 51408 30870
rect 51356 30806 51408 30812
rect 51264 28756 51316 28762
rect 51264 28698 51316 28704
rect 51368 28626 51396 30806
rect 51632 30592 51684 30598
rect 51632 30534 51684 30540
rect 51644 30258 51672 30534
rect 51632 30252 51684 30258
rect 51632 30194 51684 30200
rect 51724 30116 51776 30122
rect 51724 30058 51776 30064
rect 51540 29572 51592 29578
rect 51540 29514 51592 29520
rect 51356 28620 51408 28626
rect 51356 28562 51408 28568
rect 49332 28552 49384 28558
rect 49160 28512 49332 28540
rect 49332 28494 49384 28500
rect 49608 28552 49660 28558
rect 49608 28494 49660 28500
rect 49148 27668 49200 27674
rect 49148 27610 49200 27616
rect 49160 27470 49188 27610
rect 49344 27470 49372 28494
rect 51264 28484 51316 28490
rect 51264 28426 51316 28432
rect 50294 28316 50602 28336
rect 50294 28314 50300 28316
rect 50356 28314 50380 28316
rect 50436 28314 50460 28316
rect 50516 28314 50540 28316
rect 50596 28314 50602 28316
rect 50356 28262 50358 28314
rect 50538 28262 50540 28314
rect 50294 28260 50300 28262
rect 50356 28260 50380 28262
rect 50436 28260 50460 28262
rect 50516 28260 50540 28262
rect 50596 28260 50602 28262
rect 50294 28240 50602 28260
rect 51080 28076 51132 28082
rect 51080 28018 51132 28024
rect 51092 27554 51120 28018
rect 51276 27674 51304 28426
rect 51368 28218 51396 28562
rect 51356 28212 51408 28218
rect 51356 28154 51408 28160
rect 51356 28076 51408 28082
rect 51356 28018 51408 28024
rect 51264 27668 51316 27674
rect 51264 27610 51316 27616
rect 51092 27526 51304 27554
rect 51276 27470 51304 27526
rect 49148 27464 49200 27470
rect 49148 27406 49200 27412
rect 49332 27464 49384 27470
rect 49332 27406 49384 27412
rect 50712 27464 50764 27470
rect 50712 27406 50764 27412
rect 51264 27464 51316 27470
rect 51264 27406 51316 27412
rect 49344 26042 49372 27406
rect 50294 27228 50602 27248
rect 50294 27226 50300 27228
rect 50356 27226 50380 27228
rect 50436 27226 50460 27228
rect 50516 27226 50540 27228
rect 50596 27226 50602 27228
rect 50356 27174 50358 27226
rect 50538 27174 50540 27226
rect 50294 27172 50300 27174
rect 50356 27172 50380 27174
rect 50436 27172 50460 27174
rect 50516 27172 50540 27174
rect 50596 27172 50602 27174
rect 50294 27152 50602 27172
rect 50724 26586 50752 27406
rect 51172 27328 51224 27334
rect 51172 27270 51224 27276
rect 51184 27062 51212 27270
rect 51276 27130 51304 27406
rect 51368 27402 51396 28018
rect 51448 27872 51500 27878
rect 51448 27814 51500 27820
rect 51356 27396 51408 27402
rect 51356 27338 51408 27344
rect 51460 27282 51488 27814
rect 51368 27254 51488 27282
rect 51264 27124 51316 27130
rect 51264 27066 51316 27072
rect 51368 27062 51396 27254
rect 51172 27056 51224 27062
rect 51172 26998 51224 27004
rect 51356 27056 51408 27062
rect 51356 26998 51408 27004
rect 50896 26988 50948 26994
rect 50896 26930 50948 26936
rect 50712 26580 50764 26586
rect 50712 26522 50764 26528
rect 50908 26450 50936 26930
rect 49976 26444 50028 26450
rect 49976 26386 50028 26392
rect 50896 26444 50948 26450
rect 50896 26386 50948 26392
rect 49332 26036 49384 26042
rect 49332 25978 49384 25984
rect 49240 25832 49292 25838
rect 49240 25774 49292 25780
rect 49252 25362 49280 25774
rect 49240 25356 49292 25362
rect 49240 25298 49292 25304
rect 49252 24274 49280 25298
rect 49988 25276 50016 26386
rect 51368 26382 51396 26998
rect 50068 26376 50120 26382
rect 50068 26318 50120 26324
rect 51356 26376 51408 26382
rect 51356 26318 51408 26324
rect 50080 26042 50108 26318
rect 50294 26140 50602 26160
rect 50294 26138 50300 26140
rect 50356 26138 50380 26140
rect 50436 26138 50460 26140
rect 50516 26138 50540 26140
rect 50596 26138 50602 26140
rect 50356 26086 50358 26138
rect 50538 26086 50540 26138
rect 50294 26084 50300 26086
rect 50356 26084 50380 26086
rect 50436 26084 50460 26086
rect 50516 26084 50540 26086
rect 50596 26084 50602 26086
rect 50294 26064 50602 26084
rect 50068 26036 50120 26042
rect 50068 25978 50120 25984
rect 50160 25900 50212 25906
rect 50160 25842 50212 25848
rect 50172 25498 50200 25842
rect 50160 25492 50212 25498
rect 50160 25434 50212 25440
rect 50160 25288 50212 25294
rect 49988 25248 50160 25276
rect 50160 25230 50212 25236
rect 50172 24954 50200 25230
rect 50294 25052 50602 25072
rect 50294 25050 50300 25052
rect 50356 25050 50380 25052
rect 50436 25050 50460 25052
rect 50516 25050 50540 25052
rect 50596 25050 50602 25052
rect 50356 24998 50358 25050
rect 50538 24998 50540 25050
rect 50294 24996 50300 24998
rect 50356 24996 50380 24998
rect 50436 24996 50460 24998
rect 50516 24996 50540 24998
rect 50596 24996 50602 24998
rect 50294 24976 50602 24996
rect 50160 24948 50212 24954
rect 50160 24890 50212 24896
rect 51080 24812 51132 24818
rect 51080 24754 51132 24760
rect 49516 24608 49568 24614
rect 49516 24550 49568 24556
rect 49240 24268 49292 24274
rect 49240 24210 49292 24216
rect 49528 23798 49556 24550
rect 50294 23964 50602 23984
rect 50294 23962 50300 23964
rect 50356 23962 50380 23964
rect 50436 23962 50460 23964
rect 50516 23962 50540 23964
rect 50596 23962 50602 23964
rect 50356 23910 50358 23962
rect 50538 23910 50540 23962
rect 50294 23908 50300 23910
rect 50356 23908 50380 23910
rect 50436 23908 50460 23910
rect 50516 23908 50540 23910
rect 50596 23908 50602 23910
rect 50294 23888 50602 23908
rect 49516 23792 49568 23798
rect 49516 23734 49568 23740
rect 51092 23730 51120 24754
rect 50252 23724 50304 23730
rect 50252 23666 50304 23672
rect 50620 23724 50672 23730
rect 50620 23666 50672 23672
rect 51080 23724 51132 23730
rect 51080 23666 51132 23672
rect 50264 23118 50292 23666
rect 50632 23118 50660 23666
rect 51092 23186 51120 23666
rect 51080 23180 51132 23186
rect 51080 23122 51132 23128
rect 50252 23112 50304 23118
rect 50252 23054 50304 23060
rect 50620 23112 50672 23118
rect 50620 23054 50672 23060
rect 50294 22876 50602 22896
rect 50294 22874 50300 22876
rect 50356 22874 50380 22876
rect 50436 22874 50460 22876
rect 50516 22874 50540 22876
rect 50596 22874 50602 22876
rect 50356 22822 50358 22874
rect 50538 22822 50540 22874
rect 50294 22820 50300 22822
rect 50356 22820 50380 22822
rect 50436 22820 50460 22822
rect 50516 22820 50540 22822
rect 50596 22820 50602 22822
rect 50294 22800 50602 22820
rect 50632 22710 50660 23054
rect 50620 22704 50672 22710
rect 50620 22646 50672 22652
rect 49332 22636 49384 22642
rect 49332 22578 49384 22584
rect 49700 22636 49752 22642
rect 49700 22578 49752 22584
rect 49344 21690 49372 22578
rect 49332 21684 49384 21690
rect 49332 21626 49384 21632
rect 49712 21554 49740 22578
rect 50294 21788 50602 21808
rect 50294 21786 50300 21788
rect 50356 21786 50380 21788
rect 50436 21786 50460 21788
rect 50516 21786 50540 21788
rect 50596 21786 50602 21788
rect 50356 21734 50358 21786
rect 50538 21734 50540 21786
rect 50294 21732 50300 21734
rect 50356 21732 50380 21734
rect 50436 21732 50460 21734
rect 50516 21732 50540 21734
rect 50596 21732 50602 21734
rect 50294 21712 50602 21732
rect 49700 21548 49752 21554
rect 49700 21490 49752 21496
rect 49240 21412 49292 21418
rect 49240 21354 49292 21360
rect 49252 20942 49280 21354
rect 49712 21146 49740 21490
rect 51080 21344 51132 21350
rect 51080 21286 51132 21292
rect 49700 21140 49752 21146
rect 49700 21082 49752 21088
rect 51092 21010 51120 21286
rect 51080 21004 51132 21010
rect 51080 20946 51132 20952
rect 49240 20936 49292 20942
rect 49240 20878 49292 20884
rect 50294 20700 50602 20720
rect 50294 20698 50300 20700
rect 50356 20698 50380 20700
rect 50436 20698 50460 20700
rect 50516 20698 50540 20700
rect 50596 20698 50602 20700
rect 50356 20646 50358 20698
rect 50538 20646 50540 20698
rect 50294 20644 50300 20646
rect 50356 20644 50380 20646
rect 50436 20644 50460 20646
rect 50516 20644 50540 20646
rect 50596 20644 50602 20646
rect 50294 20624 50602 20644
rect 51092 20466 51120 20946
rect 51356 20936 51408 20942
rect 51356 20878 51408 20884
rect 51368 20466 51396 20878
rect 51080 20460 51132 20466
rect 51080 20402 51132 20408
rect 51356 20460 51408 20466
rect 51356 20402 51408 20408
rect 48964 19916 49016 19922
rect 48964 19858 49016 19864
rect 48976 19378 49004 19858
rect 49884 19848 49936 19854
rect 49884 19790 49936 19796
rect 50620 19848 50672 19854
rect 50620 19790 50672 19796
rect 50712 19848 50764 19854
rect 50712 19790 50764 19796
rect 48964 19372 49016 19378
rect 48964 19314 49016 19320
rect 49516 19372 49568 19378
rect 49516 19314 49568 19320
rect 49700 19372 49752 19378
rect 49700 19314 49752 19320
rect 49528 18970 49556 19314
rect 49608 19304 49660 19310
rect 49608 19246 49660 19252
rect 49516 18964 49568 18970
rect 49516 18906 49568 18912
rect 49620 18834 49648 19246
rect 49608 18828 49660 18834
rect 49608 18770 49660 18776
rect 49712 18698 49740 19314
rect 49896 19242 49924 19790
rect 50294 19612 50602 19632
rect 50294 19610 50300 19612
rect 50356 19610 50380 19612
rect 50436 19610 50460 19612
rect 50516 19610 50540 19612
rect 50596 19610 50602 19612
rect 50356 19558 50358 19610
rect 50538 19558 50540 19610
rect 50294 19556 50300 19558
rect 50356 19556 50380 19558
rect 50436 19556 50460 19558
rect 50516 19556 50540 19558
rect 50596 19556 50602 19558
rect 50294 19536 50602 19556
rect 50632 19514 50660 19790
rect 50620 19508 50672 19514
rect 50620 19450 50672 19456
rect 50160 19372 50212 19378
rect 50160 19314 50212 19320
rect 50436 19372 50488 19378
rect 50436 19314 50488 19320
rect 49884 19236 49936 19242
rect 49884 19178 49936 19184
rect 50172 18766 50200 19314
rect 50448 18970 50476 19314
rect 50620 19304 50672 19310
rect 50620 19246 50672 19252
rect 50436 18964 50488 18970
rect 50436 18906 50488 18912
rect 50160 18760 50212 18766
rect 50160 18702 50212 18708
rect 49700 18692 49752 18698
rect 49700 18634 49752 18640
rect 48964 18284 49016 18290
rect 48964 18226 49016 18232
rect 49148 18284 49200 18290
rect 49148 18226 49200 18232
rect 48976 17678 49004 18226
rect 48964 17672 49016 17678
rect 48964 17614 49016 17620
rect 49160 17610 49188 18226
rect 49712 17882 49740 18634
rect 50172 18426 50200 18702
rect 50632 18698 50660 19246
rect 50724 19174 50752 19790
rect 50988 19780 51040 19786
rect 50988 19722 51040 19728
rect 51000 19514 51028 19722
rect 50988 19508 51040 19514
rect 50988 19450 51040 19456
rect 50712 19168 50764 19174
rect 50712 19110 50764 19116
rect 50620 18692 50672 18698
rect 50620 18634 50672 18640
rect 50294 18524 50602 18544
rect 50294 18522 50300 18524
rect 50356 18522 50380 18524
rect 50436 18522 50460 18524
rect 50516 18522 50540 18524
rect 50596 18522 50602 18524
rect 50356 18470 50358 18522
rect 50538 18470 50540 18522
rect 50294 18468 50300 18470
rect 50356 18468 50380 18470
rect 50436 18468 50460 18470
rect 50516 18468 50540 18470
rect 50596 18468 50602 18470
rect 50294 18448 50602 18468
rect 50160 18420 50212 18426
rect 50160 18362 50212 18368
rect 49700 17876 49752 17882
rect 49700 17818 49752 17824
rect 50158 17640 50214 17649
rect 49148 17604 49200 17610
rect 50158 17575 50214 17584
rect 49148 17546 49200 17552
rect 50172 16794 50200 17575
rect 50294 17436 50602 17456
rect 50294 17434 50300 17436
rect 50356 17434 50380 17436
rect 50436 17434 50460 17436
rect 50516 17434 50540 17436
rect 50596 17434 50602 17436
rect 50356 17382 50358 17434
rect 50538 17382 50540 17434
rect 50294 17380 50300 17382
rect 50356 17380 50380 17382
rect 50436 17380 50460 17382
rect 50516 17380 50540 17382
rect 50596 17380 50602 17382
rect 50294 17360 50602 17380
rect 50804 17196 50856 17202
rect 50804 17138 50856 17144
rect 50252 17128 50304 17134
rect 50252 17070 50304 17076
rect 50160 16788 50212 16794
rect 50160 16730 50212 16736
rect 50264 16726 50292 17070
rect 50816 16794 50844 17138
rect 51172 16992 51224 16998
rect 51172 16934 51224 16940
rect 50804 16788 50856 16794
rect 50804 16730 50856 16736
rect 50252 16720 50304 16726
rect 50252 16662 50304 16668
rect 51184 16658 51212 16934
rect 51172 16652 51224 16658
rect 51172 16594 51224 16600
rect 51552 16574 51580 29514
rect 51736 29306 51764 30058
rect 51724 29300 51776 29306
rect 51724 29242 51776 29248
rect 51632 28416 51684 28422
rect 51632 28358 51684 28364
rect 51644 28082 51672 28358
rect 51632 28076 51684 28082
rect 51632 28018 51684 28024
rect 51724 27872 51776 27878
rect 51724 27814 51776 27820
rect 51736 27470 51764 27814
rect 51920 27606 51948 31726
rect 52276 31690 52328 31696
rect 52288 31278 52316 31690
rect 52368 31340 52420 31346
rect 52368 31282 52420 31288
rect 52276 31272 52328 31278
rect 52276 31214 52328 31220
rect 52000 31136 52052 31142
rect 52000 31078 52052 31084
rect 52012 30546 52040 31078
rect 52288 30734 52316 31214
rect 52380 31210 52408 31282
rect 52368 31204 52420 31210
rect 52368 31146 52420 31152
rect 52380 30734 52408 31146
rect 52276 30728 52328 30734
rect 52276 30670 52328 30676
rect 52368 30728 52420 30734
rect 52368 30670 52420 30676
rect 52184 30660 52236 30666
rect 52184 30602 52236 30608
rect 52012 30518 52132 30546
rect 52104 30190 52132 30518
rect 52092 30184 52144 30190
rect 52092 30126 52144 30132
rect 52104 29646 52132 30126
rect 52092 29640 52144 29646
rect 52092 29582 52144 29588
rect 51908 27600 51960 27606
rect 51908 27542 51960 27548
rect 51724 27464 51776 27470
rect 51724 27406 51776 27412
rect 52092 23520 52144 23526
rect 52092 23462 52144 23468
rect 52104 23186 52132 23462
rect 52092 23180 52144 23186
rect 52092 23122 52144 23128
rect 52104 22642 52132 23122
rect 52092 22636 52144 22642
rect 52092 22578 52144 22584
rect 52196 22094 52224 30602
rect 52368 27600 52420 27606
rect 52368 27542 52420 27548
rect 52276 26308 52328 26314
rect 52276 26250 52328 26256
rect 52288 25838 52316 26250
rect 52380 25906 52408 27542
rect 52460 26308 52512 26314
rect 52460 26250 52512 26256
rect 52472 25945 52500 26250
rect 52458 25936 52514 25945
rect 52368 25900 52420 25906
rect 52458 25871 52514 25880
rect 52368 25842 52420 25848
rect 52276 25832 52328 25838
rect 52276 25774 52328 25780
rect 52380 25362 52408 25842
rect 52564 25430 52592 37198
rect 54128 37126 54156 39200
rect 56060 37262 56088 39200
rect 57886 37496 57942 37505
rect 57886 37431 57942 37440
rect 54208 37256 54260 37262
rect 54208 37198 54260 37204
rect 56048 37256 56100 37262
rect 56048 37198 56100 37204
rect 54116 37120 54168 37126
rect 54116 37062 54168 37068
rect 54220 35222 54248 37198
rect 56692 37188 56744 37194
rect 56692 37130 56744 37136
rect 56600 37120 56652 37126
rect 56600 37062 56652 37068
rect 56612 36718 56640 37062
rect 56600 36712 56652 36718
rect 56600 36654 56652 36660
rect 56600 36576 56652 36582
rect 56600 36518 56652 36524
rect 54208 35216 54260 35222
rect 54208 35158 54260 35164
rect 53564 35080 53616 35086
rect 53564 35022 53616 35028
rect 53576 34746 53604 35022
rect 53564 34740 53616 34746
rect 53564 34682 53616 34688
rect 52644 34604 52696 34610
rect 52644 34546 52696 34552
rect 52828 34604 52880 34610
rect 52828 34546 52880 34552
rect 53472 34604 53524 34610
rect 53472 34546 53524 34552
rect 52656 33522 52684 34546
rect 52644 33516 52696 33522
rect 52644 33458 52696 33464
rect 52840 33318 52868 34546
rect 52920 34400 52972 34406
rect 52920 34342 52972 34348
rect 52932 33998 52960 34342
rect 53484 34066 53512 34546
rect 53472 34060 53524 34066
rect 53472 34002 53524 34008
rect 52920 33992 52972 33998
rect 52920 33934 52972 33940
rect 53484 33386 53512 34002
rect 55588 33924 55640 33930
rect 55588 33866 55640 33872
rect 53472 33380 53524 33386
rect 53472 33322 53524 33328
rect 52828 33312 52880 33318
rect 52828 33254 52880 33260
rect 52920 32836 52972 32842
rect 52920 32778 52972 32784
rect 52932 32434 52960 32778
rect 52920 32428 52972 32434
rect 52920 32370 52972 32376
rect 52736 32224 52788 32230
rect 52736 32166 52788 32172
rect 52748 31414 52776 32166
rect 52932 31822 52960 32370
rect 53288 32360 53340 32366
rect 53288 32302 53340 32308
rect 53300 32026 53328 32302
rect 53288 32020 53340 32026
rect 53288 31962 53340 31968
rect 53300 31822 53328 31962
rect 52920 31816 52972 31822
rect 52920 31758 52972 31764
rect 53288 31816 53340 31822
rect 53288 31758 53340 31764
rect 55496 31816 55548 31822
rect 55496 31758 55548 31764
rect 52736 31408 52788 31414
rect 54944 31408 54996 31414
rect 52736 31350 52788 31356
rect 54942 31376 54944 31385
rect 54996 31376 54998 31385
rect 54942 31311 54998 31320
rect 55404 31340 55456 31346
rect 55404 31282 55456 31288
rect 55312 31272 55364 31278
rect 55312 31214 55364 31220
rect 55324 30802 55352 31214
rect 55312 30796 55364 30802
rect 55312 30738 55364 30744
rect 55324 30394 55352 30738
rect 55416 30394 55444 31282
rect 55508 30938 55536 31758
rect 55496 30932 55548 30938
rect 55496 30874 55548 30880
rect 55312 30388 55364 30394
rect 55312 30330 55364 30336
rect 55404 30388 55456 30394
rect 55404 30330 55456 30336
rect 55312 30252 55364 30258
rect 55312 30194 55364 30200
rect 53012 30048 53064 30054
rect 53012 29990 53064 29996
rect 53024 29646 53052 29990
rect 55220 29708 55272 29714
rect 55220 29650 55272 29656
rect 53012 29640 53064 29646
rect 53012 29582 53064 29588
rect 53932 27464 53984 27470
rect 53932 27406 53984 27412
rect 52644 27396 52696 27402
rect 52644 27338 52696 27344
rect 52552 25424 52604 25430
rect 52552 25366 52604 25372
rect 52368 25356 52420 25362
rect 52368 25298 52420 25304
rect 52276 25152 52328 25158
rect 52276 25094 52328 25100
rect 52288 24206 52316 25094
rect 52276 24200 52328 24206
rect 52276 24142 52328 24148
rect 52288 23730 52316 24142
rect 52276 23724 52328 23730
rect 52276 23666 52328 23672
rect 52276 23588 52328 23594
rect 52276 23530 52328 23536
rect 52288 23118 52316 23530
rect 52276 23112 52328 23118
rect 52276 23054 52328 23060
rect 52288 22710 52316 23054
rect 52276 22704 52328 22710
rect 52276 22646 52328 22652
rect 52196 22066 52408 22094
rect 51724 21480 51776 21486
rect 51724 21422 51776 21428
rect 51736 21146 51764 21422
rect 51816 21344 51868 21350
rect 51816 21286 51868 21292
rect 51724 21140 51776 21146
rect 51724 21082 51776 21088
rect 51724 21004 51776 21010
rect 51724 20946 51776 20952
rect 51736 20466 51764 20946
rect 51828 20602 51856 21286
rect 52000 20936 52052 20942
rect 52000 20878 52052 20884
rect 51816 20596 51868 20602
rect 51816 20538 51868 20544
rect 51724 20460 51776 20466
rect 51724 20402 51776 20408
rect 51736 19174 51764 20402
rect 52012 20398 52040 20878
rect 52000 20392 52052 20398
rect 52000 20334 52052 20340
rect 52012 19718 52040 20334
rect 52000 19712 52052 19718
rect 52000 19654 52052 19660
rect 51724 19168 51776 19174
rect 51724 19110 51776 19116
rect 51736 18970 51764 19110
rect 51724 18964 51776 18970
rect 51724 18906 51776 18912
rect 51632 16992 51684 16998
rect 51632 16934 51684 16940
rect 51816 16992 51868 16998
rect 51816 16934 51868 16940
rect 51644 16658 51672 16934
rect 51632 16652 51684 16658
rect 51632 16594 51684 16600
rect 51828 16590 51856 16934
rect 51368 16546 51580 16574
rect 51816 16584 51868 16590
rect 50294 16348 50602 16368
rect 50294 16346 50300 16348
rect 50356 16346 50380 16348
rect 50436 16346 50460 16348
rect 50516 16346 50540 16348
rect 50596 16346 50602 16348
rect 50356 16294 50358 16346
rect 50538 16294 50540 16346
rect 50294 16292 50300 16294
rect 50356 16292 50380 16294
rect 50436 16292 50460 16294
rect 50516 16292 50540 16294
rect 50596 16292 50602 16294
rect 50294 16272 50602 16292
rect 49976 15496 50028 15502
rect 49976 15438 50028 15444
rect 50068 15496 50120 15502
rect 50068 15438 50120 15444
rect 49700 15360 49752 15366
rect 49700 15302 49752 15308
rect 49712 15026 49740 15302
rect 49988 15026 50016 15438
rect 49700 15020 49752 15026
rect 49700 14962 49752 14968
rect 49976 15020 50028 15026
rect 49976 14962 50028 14968
rect 49790 14920 49846 14929
rect 50080 14890 50108 15438
rect 50160 15360 50212 15366
rect 50160 15302 50212 15308
rect 50172 15162 50200 15302
rect 50294 15260 50602 15280
rect 50294 15258 50300 15260
rect 50356 15258 50380 15260
rect 50436 15258 50460 15260
rect 50516 15258 50540 15260
rect 50596 15258 50602 15260
rect 50356 15206 50358 15258
rect 50538 15206 50540 15258
rect 50294 15204 50300 15206
rect 50356 15204 50380 15206
rect 50436 15204 50460 15206
rect 50516 15204 50540 15206
rect 50596 15204 50602 15206
rect 50294 15184 50602 15204
rect 50160 15156 50212 15162
rect 50160 15098 50212 15104
rect 50252 15088 50304 15094
rect 50252 15030 50304 15036
rect 49790 14855 49846 14864
rect 50068 14884 50120 14890
rect 49804 14074 49832 14855
rect 50068 14826 50120 14832
rect 50160 14816 50212 14822
rect 50160 14758 50212 14764
rect 50172 14414 50200 14758
rect 50264 14414 50292 15030
rect 50436 15020 50488 15026
rect 50436 14962 50488 14968
rect 50448 14414 50476 14962
rect 50160 14408 50212 14414
rect 50160 14350 50212 14356
rect 50252 14408 50304 14414
rect 50252 14350 50304 14356
rect 50436 14408 50488 14414
rect 50436 14350 50488 14356
rect 50294 14172 50602 14192
rect 50294 14170 50300 14172
rect 50356 14170 50380 14172
rect 50436 14170 50460 14172
rect 50516 14170 50540 14172
rect 50596 14170 50602 14172
rect 50356 14118 50358 14170
rect 50538 14118 50540 14170
rect 50294 14116 50300 14118
rect 50356 14116 50380 14118
rect 50436 14116 50460 14118
rect 50516 14116 50540 14118
rect 50596 14116 50602 14118
rect 50294 14096 50602 14116
rect 49792 14068 49844 14074
rect 49792 14010 49844 14016
rect 50712 14068 50764 14074
rect 50712 14010 50764 14016
rect 50724 13394 50752 14010
rect 50712 13388 50764 13394
rect 50712 13330 50764 13336
rect 50294 13084 50602 13104
rect 50294 13082 50300 13084
rect 50356 13082 50380 13084
rect 50436 13082 50460 13084
rect 50516 13082 50540 13084
rect 50596 13082 50602 13084
rect 50356 13030 50358 13082
rect 50538 13030 50540 13082
rect 50294 13028 50300 13030
rect 50356 13028 50380 13030
rect 50436 13028 50460 13030
rect 50516 13028 50540 13030
rect 50596 13028 50602 13030
rect 50294 13008 50602 13028
rect 50724 12986 50752 13330
rect 50804 13320 50856 13326
rect 50804 13262 50856 13268
rect 50712 12980 50764 12986
rect 50712 12922 50764 12928
rect 50816 12850 50844 13262
rect 51172 13184 51224 13190
rect 51172 13126 51224 13132
rect 51184 12850 51212 13126
rect 50804 12844 50856 12850
rect 50804 12786 50856 12792
rect 51172 12844 51224 12850
rect 51172 12786 51224 12792
rect 49056 12640 49108 12646
rect 49056 12582 49108 12588
rect 49068 12238 49096 12582
rect 49056 12232 49108 12238
rect 49056 12174 49108 12180
rect 48964 12164 49016 12170
rect 48964 12106 49016 12112
rect 48976 11694 49004 12106
rect 49068 11762 49096 12174
rect 51172 12164 51224 12170
rect 51172 12106 51224 12112
rect 50294 11996 50602 12016
rect 50294 11994 50300 11996
rect 50356 11994 50380 11996
rect 50436 11994 50460 11996
rect 50516 11994 50540 11996
rect 50596 11994 50602 11996
rect 50356 11942 50358 11994
rect 50538 11942 50540 11994
rect 50294 11940 50300 11942
rect 50356 11940 50380 11942
rect 50436 11940 50460 11942
rect 50516 11940 50540 11942
rect 50596 11940 50602 11942
rect 50294 11920 50602 11940
rect 51184 11898 51212 12106
rect 51172 11892 51224 11898
rect 51172 11834 51224 11840
rect 49056 11756 49108 11762
rect 49056 11698 49108 11704
rect 48964 11688 49016 11694
rect 48964 11630 49016 11636
rect 48964 11008 49016 11014
rect 48964 10950 49016 10956
rect 48976 10674 49004 10950
rect 50294 10908 50602 10928
rect 50294 10906 50300 10908
rect 50356 10906 50380 10908
rect 50436 10906 50460 10908
rect 50516 10906 50540 10908
rect 50596 10906 50602 10908
rect 50356 10854 50358 10906
rect 50538 10854 50540 10906
rect 50294 10852 50300 10854
rect 50356 10852 50380 10854
rect 50436 10852 50460 10854
rect 50516 10852 50540 10854
rect 50596 10852 50602 10854
rect 50294 10832 50602 10852
rect 48964 10668 49016 10674
rect 48964 10610 49016 10616
rect 49516 10600 49568 10606
rect 49516 10542 49568 10548
rect 49148 9036 49200 9042
rect 49148 8978 49200 8984
rect 48964 8968 49016 8974
rect 48964 8910 49016 8916
rect 48976 8498 49004 8910
rect 49160 8498 49188 8978
rect 48964 8492 49016 8498
rect 48964 8434 49016 8440
rect 49148 8492 49200 8498
rect 49148 8434 49200 8440
rect 49160 8022 49188 8434
rect 49148 8016 49200 8022
rect 49148 7958 49200 7964
rect 49528 6798 49556 10542
rect 51170 10024 51226 10033
rect 51170 9959 51172 9968
rect 51224 9959 51226 9968
rect 51172 9930 51224 9936
rect 50294 9820 50602 9840
rect 50294 9818 50300 9820
rect 50356 9818 50380 9820
rect 50436 9818 50460 9820
rect 50516 9818 50540 9820
rect 50596 9818 50602 9820
rect 50356 9766 50358 9818
rect 50538 9766 50540 9818
rect 50294 9764 50300 9766
rect 50356 9764 50380 9766
rect 50436 9764 50460 9766
rect 50516 9764 50540 9766
rect 50596 9764 50602 9766
rect 50294 9744 50602 9764
rect 50294 8732 50602 8752
rect 50294 8730 50300 8732
rect 50356 8730 50380 8732
rect 50436 8730 50460 8732
rect 50516 8730 50540 8732
rect 50596 8730 50602 8732
rect 50356 8678 50358 8730
rect 50538 8678 50540 8730
rect 50294 8676 50300 8678
rect 50356 8676 50380 8678
rect 50436 8676 50460 8678
rect 50516 8676 50540 8678
rect 50596 8676 50602 8678
rect 50294 8656 50602 8676
rect 50294 7644 50602 7664
rect 50294 7642 50300 7644
rect 50356 7642 50380 7644
rect 50436 7642 50460 7644
rect 50516 7642 50540 7644
rect 50596 7642 50602 7644
rect 50356 7590 50358 7642
rect 50538 7590 50540 7642
rect 50294 7588 50300 7590
rect 50356 7588 50380 7590
rect 50436 7588 50460 7590
rect 50516 7588 50540 7590
rect 50596 7588 50602 7590
rect 50294 7568 50602 7588
rect 51264 6996 51316 7002
rect 51264 6938 51316 6944
rect 49516 6792 49568 6798
rect 49516 6734 49568 6740
rect 49056 6656 49108 6662
rect 49056 6598 49108 6604
rect 49068 6322 49096 6598
rect 49528 6322 49556 6734
rect 50294 6556 50602 6576
rect 50294 6554 50300 6556
rect 50356 6554 50380 6556
rect 50436 6554 50460 6556
rect 50516 6554 50540 6556
rect 50596 6554 50602 6556
rect 50356 6502 50358 6554
rect 50538 6502 50540 6554
rect 50294 6500 50300 6502
rect 50356 6500 50380 6502
rect 50436 6500 50460 6502
rect 50516 6500 50540 6502
rect 50596 6500 50602 6502
rect 50294 6480 50602 6500
rect 51276 6322 51304 6938
rect 49056 6316 49108 6322
rect 49056 6258 49108 6264
rect 49516 6316 49568 6322
rect 49516 6258 49568 6264
rect 51264 6316 51316 6322
rect 51264 6258 51316 6264
rect 50294 5468 50602 5488
rect 50294 5466 50300 5468
rect 50356 5466 50380 5468
rect 50436 5466 50460 5468
rect 50516 5466 50540 5468
rect 50596 5466 50602 5468
rect 50356 5414 50358 5466
rect 50538 5414 50540 5466
rect 50294 5412 50300 5414
rect 50356 5412 50380 5414
rect 50436 5412 50460 5414
rect 50516 5412 50540 5414
rect 50596 5412 50602 5414
rect 50294 5392 50602 5412
rect 50294 4380 50602 4400
rect 50294 4378 50300 4380
rect 50356 4378 50380 4380
rect 50436 4378 50460 4380
rect 50516 4378 50540 4380
rect 50596 4378 50602 4380
rect 50356 4326 50358 4378
rect 50538 4326 50540 4378
rect 50294 4324 50300 4326
rect 50356 4324 50380 4326
rect 50436 4324 50460 4326
rect 50516 4324 50540 4326
rect 50596 4324 50602 4326
rect 50294 4304 50602 4324
rect 50294 3292 50602 3312
rect 50294 3290 50300 3292
rect 50356 3290 50380 3292
rect 50436 3290 50460 3292
rect 50516 3290 50540 3292
rect 50596 3290 50602 3292
rect 50356 3238 50358 3290
rect 50538 3238 50540 3290
rect 50294 3236 50300 3238
rect 50356 3236 50380 3238
rect 50436 3236 50460 3238
rect 50516 3236 50540 3238
rect 50596 3236 50602 3238
rect 50294 3216 50602 3236
rect 51368 2802 51396 16546
rect 51816 16526 51868 16532
rect 52276 15632 52328 15638
rect 52276 15574 52328 15580
rect 52288 14958 52316 15574
rect 52276 14952 52328 14958
rect 52276 14894 52328 14900
rect 52288 14482 52316 14894
rect 52276 14476 52328 14482
rect 52276 14418 52328 14424
rect 51448 12844 51500 12850
rect 51448 12786 51500 12792
rect 51460 12238 51488 12786
rect 51632 12776 51684 12782
rect 51632 12718 51684 12724
rect 51644 12238 51672 12718
rect 51724 12640 51776 12646
rect 51724 12582 51776 12588
rect 51736 12306 51764 12582
rect 51724 12300 51776 12306
rect 51724 12242 51776 12248
rect 51448 12232 51500 12238
rect 51448 12174 51500 12180
rect 51632 12232 51684 12238
rect 51632 12174 51684 12180
rect 51908 12164 51960 12170
rect 51908 12106 51960 12112
rect 51540 11144 51592 11150
rect 51540 11086 51592 11092
rect 51552 10606 51580 11086
rect 51816 11008 51868 11014
rect 51816 10950 51868 10956
rect 51828 10742 51856 10950
rect 51816 10736 51868 10742
rect 51722 10704 51778 10713
rect 51816 10678 51868 10684
rect 51722 10639 51724 10648
rect 51776 10639 51778 10648
rect 51724 10610 51776 10616
rect 51540 10600 51592 10606
rect 51540 10542 51592 10548
rect 51448 8968 51500 8974
rect 51448 8910 51500 8916
rect 51460 8498 51488 8910
rect 51552 8634 51580 10542
rect 51736 10266 51764 10610
rect 51724 10260 51776 10266
rect 51724 10202 51776 10208
rect 51828 10062 51856 10678
rect 51816 10056 51868 10062
rect 51816 9998 51868 10004
rect 51816 9036 51868 9042
rect 51816 8978 51868 8984
rect 51540 8628 51592 8634
rect 51540 8570 51592 8576
rect 51828 8498 51856 8978
rect 51448 8492 51500 8498
rect 51448 8434 51500 8440
rect 51816 8492 51868 8498
rect 51816 8434 51868 8440
rect 51920 7886 51948 12106
rect 52092 10668 52144 10674
rect 52092 10610 52144 10616
rect 52104 9994 52132 10610
rect 52092 9988 52144 9994
rect 52092 9930 52144 9936
rect 52092 8492 52144 8498
rect 52092 8434 52144 8440
rect 52104 8022 52132 8434
rect 52092 8016 52144 8022
rect 52092 7958 52144 7964
rect 51632 7880 51684 7886
rect 51632 7822 51684 7828
rect 51908 7880 51960 7886
rect 51908 7822 51960 7828
rect 51644 7410 51672 7822
rect 51632 7404 51684 7410
rect 51632 7346 51684 7352
rect 51644 7002 51672 7346
rect 51920 7342 51948 7822
rect 51908 7336 51960 7342
rect 51908 7278 51960 7284
rect 51632 6996 51684 7002
rect 51632 6938 51684 6944
rect 48792 2746 48912 2774
rect 51092 2774 51396 2802
rect 48504 2576 48556 2582
rect 48504 2518 48556 2524
rect 47676 2304 47728 2310
rect 47676 2246 47728 2252
rect 46480 2032 46532 2038
rect 46480 1974 46532 1980
rect 47688 800 47716 2246
rect 48516 2106 48544 2518
rect 48504 2100 48556 2106
rect 48504 2042 48556 2048
rect 48792 1970 48820 2746
rect 51092 2666 51120 2774
rect 51000 2650 51120 2666
rect 52380 2650 52408 22066
rect 52552 18896 52604 18902
rect 52552 18838 52604 18844
rect 52564 18766 52592 18838
rect 52552 18760 52604 18766
rect 52552 18702 52604 18708
rect 52552 17536 52604 17542
rect 52552 17478 52604 17484
rect 52564 17202 52592 17478
rect 52552 17196 52604 17202
rect 52552 17138 52604 17144
rect 52564 16658 52592 17138
rect 52552 16652 52604 16658
rect 52552 16594 52604 16600
rect 52552 15700 52604 15706
rect 52552 15642 52604 15648
rect 52564 15026 52592 15642
rect 52552 15020 52604 15026
rect 52552 14962 52604 14968
rect 52552 12708 52604 12714
rect 52552 12650 52604 12656
rect 52460 12640 52512 12646
rect 52460 12582 52512 12588
rect 52472 12238 52500 12582
rect 52460 12232 52512 12238
rect 52460 12174 52512 12180
rect 52564 8566 52592 12650
rect 52552 8560 52604 8566
rect 52552 8502 52604 8508
rect 52564 7886 52592 8502
rect 52552 7880 52604 7886
rect 52552 7822 52604 7828
rect 52656 6914 52684 27338
rect 53380 26988 53432 26994
rect 53380 26930 53432 26936
rect 53392 26586 53420 26930
rect 53380 26580 53432 26586
rect 53380 26522 53432 26528
rect 52828 26376 52880 26382
rect 52828 26318 52880 26324
rect 52840 26042 52868 26318
rect 53656 26308 53708 26314
rect 53656 26250 53708 26256
rect 53196 26240 53248 26246
rect 53196 26182 53248 26188
rect 53208 26042 53236 26182
rect 52828 26036 52880 26042
rect 52828 25978 52880 25984
rect 53196 26036 53248 26042
rect 53196 25978 53248 25984
rect 52840 25498 52868 25978
rect 53104 25900 53156 25906
rect 53104 25842 53156 25848
rect 52920 25832 52972 25838
rect 52920 25774 52972 25780
rect 52828 25492 52880 25498
rect 52828 25434 52880 25440
rect 52932 25362 52960 25774
rect 53116 25514 53144 25842
rect 53208 25702 53236 25978
rect 53668 25974 53696 26250
rect 53656 25968 53708 25974
rect 53656 25910 53708 25916
rect 53196 25696 53248 25702
rect 53196 25638 53248 25644
rect 53116 25486 53236 25514
rect 52920 25356 52972 25362
rect 52920 25298 52972 25304
rect 52932 24886 52960 25298
rect 53208 25294 53236 25486
rect 53196 25288 53248 25294
rect 53196 25230 53248 25236
rect 53656 25288 53708 25294
rect 53656 25230 53708 25236
rect 52920 24880 52972 24886
rect 52920 24822 52972 24828
rect 53208 24818 53236 25230
rect 53196 24812 53248 24818
rect 53196 24754 53248 24760
rect 52828 24268 52880 24274
rect 52828 24210 52880 24216
rect 52736 24200 52788 24206
rect 52736 24142 52788 24148
rect 52748 23662 52776 24142
rect 52736 23656 52788 23662
rect 52736 23598 52788 23604
rect 52748 23254 52776 23598
rect 52840 23526 52868 24210
rect 53208 23866 53236 24754
rect 53668 24206 53696 25230
rect 53944 24954 53972 27406
rect 55128 27396 55180 27402
rect 55128 27338 55180 27344
rect 55140 26994 55168 27338
rect 54024 26988 54076 26994
rect 54024 26930 54076 26936
rect 55128 26988 55180 26994
rect 55128 26930 55180 26936
rect 54036 26042 54064 26930
rect 54024 26036 54076 26042
rect 54024 25978 54076 25984
rect 53932 24948 53984 24954
rect 53932 24890 53984 24896
rect 53656 24200 53708 24206
rect 53656 24142 53708 24148
rect 53196 23860 53248 23866
rect 53196 23802 53248 23808
rect 52828 23520 52880 23526
rect 52828 23462 52880 23468
rect 52736 23248 52788 23254
rect 52736 23190 52788 23196
rect 52840 22778 52868 23462
rect 53288 23180 53340 23186
rect 53288 23122 53340 23128
rect 53012 23112 53064 23118
rect 53012 23054 53064 23060
rect 52828 22772 52880 22778
rect 52828 22714 52880 22720
rect 53024 22642 53052 23054
rect 53300 22642 53328 23122
rect 53668 22642 53696 24142
rect 54484 23112 54536 23118
rect 54484 23054 54536 23060
rect 53748 23044 53800 23050
rect 53748 22986 53800 22992
rect 53760 22710 53788 22986
rect 54496 22982 54524 23054
rect 54484 22976 54536 22982
rect 54484 22918 54536 22924
rect 53748 22704 53800 22710
rect 53748 22646 53800 22652
rect 53012 22636 53064 22642
rect 53012 22578 53064 22584
rect 53288 22636 53340 22642
rect 53288 22578 53340 22584
rect 53656 22636 53708 22642
rect 53656 22578 53708 22584
rect 53024 21690 53052 22578
rect 53300 21690 53328 22578
rect 54496 22506 54524 22918
rect 54484 22500 54536 22506
rect 54484 22442 54536 22448
rect 54496 21690 54524 22442
rect 53012 21684 53064 21690
rect 53012 21626 53064 21632
rect 53288 21684 53340 21690
rect 53288 21626 53340 21632
rect 54484 21684 54536 21690
rect 54484 21626 54536 21632
rect 53748 21616 53800 21622
rect 53748 21558 53800 21564
rect 53760 21146 53788 21558
rect 54116 21548 54168 21554
rect 54116 21490 54168 21496
rect 54208 21548 54260 21554
rect 54208 21490 54260 21496
rect 53748 21140 53800 21146
rect 53748 21082 53800 21088
rect 54128 21010 54156 21490
rect 54116 21004 54168 21010
rect 54116 20946 54168 20952
rect 54220 20942 54248 21490
rect 54392 21004 54444 21010
rect 54392 20946 54444 20952
rect 54208 20936 54260 20942
rect 54208 20878 54260 20884
rect 54024 20256 54076 20262
rect 54024 20198 54076 20204
rect 53472 19848 53524 19854
rect 53472 19790 53524 19796
rect 53932 19848 53984 19854
rect 53932 19790 53984 19796
rect 53484 19378 53512 19790
rect 53564 19712 53616 19718
rect 53564 19654 53616 19660
rect 53472 19372 53524 19378
rect 53472 19314 53524 19320
rect 52736 19304 52788 19310
rect 52736 19246 52788 19252
rect 52748 18630 52776 19246
rect 53484 18970 53512 19314
rect 53576 19310 53604 19654
rect 53944 19310 53972 19790
rect 53564 19304 53616 19310
rect 53564 19246 53616 19252
rect 53932 19304 53984 19310
rect 53932 19246 53984 19252
rect 53196 18964 53248 18970
rect 53196 18906 53248 18912
rect 53472 18964 53524 18970
rect 53472 18906 53524 18912
rect 53208 18766 53236 18906
rect 53196 18760 53248 18766
rect 53196 18702 53248 18708
rect 53472 18760 53524 18766
rect 53524 18720 53604 18748
rect 53472 18702 53524 18708
rect 53380 18692 53432 18698
rect 53380 18634 53432 18640
rect 52736 18624 52788 18630
rect 52736 18566 52788 18572
rect 53392 18426 53420 18634
rect 53380 18420 53432 18426
rect 53380 18362 53432 18368
rect 53472 18284 53524 18290
rect 53472 18226 53524 18232
rect 53380 18080 53432 18086
rect 53380 18022 53432 18028
rect 52736 17876 52788 17882
rect 52736 17818 52788 17824
rect 52748 17066 52776 17818
rect 53392 17678 53420 18022
rect 53484 17882 53512 18226
rect 53472 17876 53524 17882
rect 53472 17818 53524 17824
rect 53380 17672 53432 17678
rect 53432 17620 53512 17626
rect 53380 17614 53512 17620
rect 53392 17598 53512 17614
rect 53392 17549 53420 17598
rect 53104 17332 53156 17338
rect 53104 17274 53156 17280
rect 52736 17060 52788 17066
rect 52736 17002 52788 17008
rect 53116 16726 53144 17274
rect 53196 17196 53248 17202
rect 53196 17138 53248 17144
rect 53104 16720 53156 16726
rect 53104 16662 53156 16668
rect 53116 16454 53144 16662
rect 53208 16590 53236 17138
rect 53484 17134 53512 17598
rect 53576 17542 53604 18720
rect 53656 18284 53708 18290
rect 53656 18226 53708 18232
rect 53668 17746 53696 18226
rect 53656 17740 53708 17746
rect 53708 17700 53788 17728
rect 53656 17682 53708 17688
rect 53564 17536 53616 17542
rect 53564 17478 53616 17484
rect 53760 17202 53788 17700
rect 53656 17196 53708 17202
rect 53656 17138 53708 17144
rect 53748 17196 53800 17202
rect 53748 17138 53800 17144
rect 53472 17128 53524 17134
rect 53472 17070 53524 17076
rect 53484 16794 53512 17070
rect 53668 16794 53696 17138
rect 53760 16794 53788 17138
rect 53472 16788 53524 16794
rect 53472 16730 53524 16736
rect 53656 16788 53708 16794
rect 53656 16730 53708 16736
rect 53748 16788 53800 16794
rect 53748 16730 53800 16736
rect 53196 16584 53248 16590
rect 53196 16526 53248 16532
rect 53104 16448 53156 16454
rect 53104 16390 53156 16396
rect 52920 16108 52972 16114
rect 52920 16050 52972 16056
rect 52828 16040 52880 16046
rect 52828 15982 52880 15988
rect 52840 15570 52868 15982
rect 52828 15564 52880 15570
rect 52828 15506 52880 15512
rect 52840 14890 52868 15506
rect 52932 15502 52960 16050
rect 53012 15904 53064 15910
rect 53012 15846 53064 15852
rect 53024 15638 53052 15846
rect 53116 15706 53144 16390
rect 53208 16250 53236 16526
rect 53196 16244 53248 16250
rect 53196 16186 53248 16192
rect 53104 15700 53156 15706
rect 53104 15642 53156 15648
rect 53012 15632 53064 15638
rect 53012 15574 53064 15580
rect 53562 15600 53618 15609
rect 52920 15496 52972 15502
rect 52920 15438 52972 15444
rect 52932 15094 52960 15438
rect 52920 15088 52972 15094
rect 52920 15030 52972 15036
rect 53024 14890 53052 15574
rect 53562 15535 53564 15544
rect 53616 15535 53618 15544
rect 53564 15506 53616 15512
rect 53576 15094 53604 15506
rect 53564 15088 53616 15094
rect 53564 15030 53616 15036
rect 53380 15020 53432 15026
rect 53380 14962 53432 14968
rect 52828 14884 52880 14890
rect 52828 14826 52880 14832
rect 53012 14884 53064 14890
rect 53012 14826 53064 14832
rect 53024 14618 53052 14826
rect 53196 14816 53248 14822
rect 53196 14758 53248 14764
rect 53012 14612 53064 14618
rect 53012 14554 53064 14560
rect 53208 13938 53236 14758
rect 53392 14618 53420 14962
rect 53380 14612 53432 14618
rect 53380 14554 53432 14560
rect 53576 14550 53604 15030
rect 53564 14544 53616 14550
rect 53564 14486 53616 14492
rect 53196 13932 53248 13938
rect 53196 13874 53248 13880
rect 53012 13864 53064 13870
rect 53012 13806 53064 13812
rect 53024 13326 53052 13806
rect 53208 13530 53236 13874
rect 53196 13524 53248 13530
rect 53196 13466 53248 13472
rect 53012 13320 53064 13326
rect 53012 13262 53064 13268
rect 53840 11756 53892 11762
rect 53840 11698 53892 11704
rect 52734 11656 52790 11665
rect 52734 11591 52790 11600
rect 52748 11286 52776 11591
rect 53288 11552 53340 11558
rect 53288 11494 53340 11500
rect 52736 11280 52788 11286
rect 52736 11222 52788 11228
rect 53300 11218 53328 11494
rect 53288 11212 53340 11218
rect 53288 11154 53340 11160
rect 53852 11150 53880 11698
rect 54036 11218 54064 20198
rect 54220 20058 54248 20878
rect 54404 20058 54432 20946
rect 54208 20052 54260 20058
rect 54208 19994 54260 20000
rect 54392 20052 54444 20058
rect 54392 19994 54444 20000
rect 54668 19780 54720 19786
rect 54668 19722 54720 19728
rect 54680 19378 54708 19722
rect 54668 19372 54720 19378
rect 54668 19314 54720 19320
rect 54484 14816 54536 14822
rect 54484 14758 54536 14764
rect 54496 14414 54524 14758
rect 54484 14408 54536 14414
rect 54484 14350 54536 14356
rect 54496 13870 54524 14350
rect 55128 14340 55180 14346
rect 55128 14282 55180 14288
rect 55140 13938 55168 14282
rect 55128 13932 55180 13938
rect 55128 13874 55180 13880
rect 54484 13864 54536 13870
rect 54484 13806 54536 13812
rect 54484 13184 54536 13190
rect 54484 13126 54536 13132
rect 54496 12986 54524 13126
rect 54484 12980 54536 12986
rect 54484 12922 54536 12928
rect 55036 12980 55088 12986
rect 55036 12922 55088 12928
rect 54496 12782 54524 12922
rect 55048 12850 55076 12922
rect 55036 12844 55088 12850
rect 55036 12786 55088 12792
rect 54484 12776 54536 12782
rect 54484 12718 54536 12724
rect 54668 11824 54720 11830
rect 54668 11766 54720 11772
rect 54024 11212 54076 11218
rect 54024 11154 54076 11160
rect 53012 11144 53064 11150
rect 53012 11086 53064 11092
rect 53840 11144 53892 11150
rect 53840 11086 53892 11092
rect 53024 10810 53052 11086
rect 53852 10810 53880 11086
rect 53012 10804 53064 10810
rect 53012 10746 53064 10752
rect 53840 10804 53892 10810
rect 53840 10746 53892 10752
rect 54036 10690 54064 11154
rect 54680 11150 54708 11766
rect 54668 11144 54720 11150
rect 54668 11086 54720 11092
rect 54036 10674 54156 10690
rect 54680 10674 54708 11086
rect 55128 10736 55180 10742
rect 55128 10678 55180 10684
rect 53656 10668 53708 10674
rect 54036 10668 54168 10674
rect 54036 10662 54116 10668
rect 53656 10610 53708 10616
rect 54116 10610 54168 10616
rect 54668 10668 54720 10674
rect 54668 10610 54720 10616
rect 53668 10266 53696 10610
rect 54024 10600 54076 10606
rect 54024 10542 54076 10548
rect 53656 10260 53708 10266
rect 53656 10202 53708 10208
rect 54036 9586 54064 10542
rect 54576 10464 54628 10470
rect 54576 10406 54628 10412
rect 54024 9580 54076 9586
rect 54024 9522 54076 9528
rect 54036 9178 54064 9522
rect 54484 9376 54536 9382
rect 54484 9318 54536 9324
rect 54024 9172 54076 9178
rect 54024 9114 54076 9120
rect 54496 8498 54524 9318
rect 52828 8492 52880 8498
rect 52828 8434 52880 8440
rect 54484 8492 54536 8498
rect 54484 8434 54536 8440
rect 52840 7954 52868 8434
rect 54588 8430 54616 10406
rect 55140 9722 55168 10678
rect 55128 9716 55180 9722
rect 55128 9658 55180 9664
rect 54576 8424 54628 8430
rect 54576 8366 54628 8372
rect 54668 8356 54720 8362
rect 54668 8298 54720 8304
rect 52828 7948 52880 7954
rect 52828 7890 52880 7896
rect 52840 7478 52868 7890
rect 52828 7472 52880 7478
rect 52828 7414 52880 7420
rect 54680 6914 54708 8298
rect 52564 6886 52684 6914
rect 54588 6886 54708 6914
rect 55232 6914 55260 29650
rect 55324 29646 55352 30194
rect 55312 29640 55364 29646
rect 55312 29582 55364 29588
rect 55324 29306 55352 29582
rect 55312 29300 55364 29306
rect 55312 29242 55364 29248
rect 55600 28082 55628 33866
rect 56324 31816 56376 31822
rect 56324 31758 56376 31764
rect 55772 30728 55824 30734
rect 55772 30670 55824 30676
rect 55680 30252 55732 30258
rect 55680 30194 55732 30200
rect 55692 29646 55720 30194
rect 55680 29640 55732 29646
rect 55680 29582 55732 29588
rect 55692 28218 55720 29582
rect 55784 29102 55812 30670
rect 56048 30592 56100 30598
rect 56048 30534 56100 30540
rect 56060 30054 56088 30534
rect 56048 30048 56100 30054
rect 56048 29990 56100 29996
rect 56060 29578 56088 29990
rect 56336 29646 56364 31758
rect 56324 29640 56376 29646
rect 56324 29582 56376 29588
rect 56048 29572 56100 29578
rect 56048 29514 56100 29520
rect 56060 29170 56088 29514
rect 56336 29306 56364 29582
rect 56324 29300 56376 29306
rect 56324 29242 56376 29248
rect 56048 29164 56100 29170
rect 56048 29106 56100 29112
rect 55772 29096 55824 29102
rect 55772 29038 55824 29044
rect 56060 28422 56088 29106
rect 56048 28416 56100 28422
rect 56048 28358 56100 28364
rect 55680 28212 55732 28218
rect 55680 28154 55732 28160
rect 55312 28076 55364 28082
rect 55312 28018 55364 28024
rect 55588 28076 55640 28082
rect 55588 28018 55640 28024
rect 55864 28076 55916 28082
rect 55864 28018 55916 28024
rect 55324 27470 55352 28018
rect 55600 27470 55628 28018
rect 55772 28008 55824 28014
rect 55772 27950 55824 27956
rect 55312 27464 55364 27470
rect 55312 27406 55364 27412
rect 55588 27464 55640 27470
rect 55588 27406 55640 27412
rect 55324 27062 55352 27406
rect 55312 27056 55364 27062
rect 55312 26998 55364 27004
rect 55784 26586 55812 27950
rect 55876 26858 55904 28018
rect 55956 27532 56008 27538
rect 55956 27474 56008 27480
rect 55968 26994 55996 27474
rect 55956 26988 56008 26994
rect 55956 26930 56008 26936
rect 55864 26852 55916 26858
rect 55864 26794 55916 26800
rect 55772 26580 55824 26586
rect 55772 26522 55824 26528
rect 55968 26382 55996 26930
rect 55956 26376 56008 26382
rect 55956 26318 56008 26324
rect 55968 26042 55996 26318
rect 55956 26036 56008 26042
rect 55956 25978 56008 25984
rect 55956 25900 56008 25906
rect 55956 25842 56008 25848
rect 55772 25832 55824 25838
rect 55772 25774 55824 25780
rect 55588 25356 55640 25362
rect 55588 25298 55640 25304
rect 55404 25288 55456 25294
rect 55404 25230 55456 25236
rect 55416 24818 55444 25230
rect 55600 24886 55628 25298
rect 55680 25152 55732 25158
rect 55680 25094 55732 25100
rect 55588 24880 55640 24886
rect 55588 24822 55640 24828
rect 55404 24812 55456 24818
rect 55404 24754 55456 24760
rect 55496 24812 55548 24818
rect 55496 24754 55548 24760
rect 55416 24206 55444 24754
rect 55508 24410 55536 24754
rect 55496 24404 55548 24410
rect 55496 24346 55548 24352
rect 55600 24206 55628 24822
rect 55692 24750 55720 25094
rect 55680 24744 55732 24750
rect 55680 24686 55732 24692
rect 55692 24206 55720 24686
rect 55312 24200 55364 24206
rect 55312 24142 55364 24148
rect 55404 24200 55456 24206
rect 55404 24142 55456 24148
rect 55588 24200 55640 24206
rect 55588 24142 55640 24148
rect 55680 24200 55732 24206
rect 55680 24142 55732 24148
rect 55324 23798 55352 24142
rect 55784 23866 55812 25774
rect 55968 25498 55996 25842
rect 55956 25492 56008 25498
rect 55956 25434 56008 25440
rect 55864 25356 55916 25362
rect 55864 25298 55916 25304
rect 55876 24818 55904 25298
rect 55864 24812 55916 24818
rect 55864 24754 55916 24760
rect 55772 23860 55824 23866
rect 55772 23802 55824 23808
rect 55312 23792 55364 23798
rect 55312 23734 55364 23740
rect 55324 23322 55352 23734
rect 55680 23724 55732 23730
rect 55680 23666 55732 23672
rect 55312 23316 55364 23322
rect 55312 23258 55364 23264
rect 55496 23316 55548 23322
rect 55496 23258 55548 23264
rect 55508 23118 55536 23258
rect 55496 23112 55548 23118
rect 55496 23054 55548 23060
rect 55508 22574 55536 23054
rect 55692 22982 55720 23666
rect 55680 22976 55732 22982
rect 55680 22918 55732 22924
rect 55496 22568 55548 22574
rect 55496 22510 55548 22516
rect 55508 20874 55536 22510
rect 55692 21894 55720 22918
rect 55680 21888 55732 21894
rect 55680 21830 55732 21836
rect 55680 21480 55732 21486
rect 55680 21422 55732 21428
rect 55692 20942 55720 21422
rect 55680 20936 55732 20942
rect 55680 20878 55732 20884
rect 55496 20868 55548 20874
rect 55496 20810 55548 20816
rect 56060 16574 56088 28358
rect 56612 27470 56640 36518
rect 56704 32502 56732 37130
rect 57900 36854 57928 37431
rect 57992 37262 58020 39200
rect 57980 37256 58032 37262
rect 57980 37198 58032 37204
rect 57992 36922 58020 37198
rect 59924 37126 59952 39200
rect 58164 37120 58216 37126
rect 58164 37062 58216 37068
rect 59912 37120 59964 37126
rect 59912 37062 59964 37068
rect 57980 36916 58032 36922
rect 57980 36858 58032 36864
rect 57888 36848 57940 36854
rect 57888 36790 57940 36796
rect 58176 36174 58204 37062
rect 58164 36168 58216 36174
rect 58164 36110 58216 36116
rect 57796 36100 57848 36106
rect 57796 36042 57848 36048
rect 56692 32496 56744 32502
rect 56692 32438 56744 32444
rect 56968 29640 57020 29646
rect 56968 29582 57020 29588
rect 57704 29640 57756 29646
rect 57704 29582 57756 29588
rect 56980 28966 57008 29582
rect 57612 29232 57664 29238
rect 57612 29174 57664 29180
rect 57428 29028 57480 29034
rect 57428 28970 57480 28976
rect 56968 28960 57020 28966
rect 56968 28902 57020 28908
rect 56980 28218 57008 28902
rect 57440 28558 57468 28970
rect 57244 28552 57296 28558
rect 57244 28494 57296 28500
rect 57428 28552 57480 28558
rect 57428 28494 57480 28500
rect 56968 28212 57020 28218
rect 56968 28154 57020 28160
rect 57256 28150 57284 28494
rect 57440 28150 57468 28494
rect 57244 28144 57296 28150
rect 57244 28086 57296 28092
rect 57428 28144 57480 28150
rect 57428 28086 57480 28092
rect 56968 27940 57020 27946
rect 56968 27882 57020 27888
rect 56980 27606 57008 27882
rect 56968 27600 57020 27606
rect 56968 27542 57020 27548
rect 56600 27464 56652 27470
rect 56600 27406 56652 27412
rect 56612 27130 56640 27406
rect 56876 27328 56928 27334
rect 56876 27270 56928 27276
rect 56600 27124 56652 27130
rect 56600 27066 56652 27072
rect 56612 26382 56640 27066
rect 56888 26926 56916 27270
rect 56980 26994 57008 27542
rect 56968 26988 57020 26994
rect 56968 26930 57020 26936
rect 56876 26920 56928 26926
rect 56876 26862 56928 26868
rect 56600 26376 56652 26382
rect 56600 26318 56652 26324
rect 57256 24818 57284 28086
rect 56968 24812 57020 24818
rect 56968 24754 57020 24760
rect 57244 24812 57296 24818
rect 57244 24754 57296 24760
rect 56980 24682 57008 24754
rect 57060 24744 57112 24750
rect 57112 24692 57192 24698
rect 57060 24686 57192 24692
rect 56968 24676 57020 24682
rect 57072 24670 57192 24686
rect 56968 24618 57020 24624
rect 56782 24168 56838 24177
rect 56692 24132 56744 24138
rect 56782 24103 56784 24112
rect 56692 24074 56744 24080
rect 56836 24103 56838 24112
rect 56784 24074 56836 24080
rect 56324 24064 56376 24070
rect 56324 24006 56376 24012
rect 56336 22642 56364 24006
rect 56508 23112 56560 23118
rect 56508 23054 56560 23060
rect 56520 22710 56548 23054
rect 56508 22704 56560 22710
rect 56508 22646 56560 22652
rect 56704 22642 56732 24074
rect 56232 22636 56284 22642
rect 56232 22578 56284 22584
rect 56324 22636 56376 22642
rect 56324 22578 56376 22584
rect 56692 22636 56744 22642
rect 56692 22578 56744 22584
rect 56244 20942 56272 22578
rect 56336 21078 56364 22578
rect 56704 21690 56732 22578
rect 56980 22094 57008 24618
rect 57164 24614 57192 24670
rect 57152 24608 57204 24614
rect 57152 24550 57204 24556
rect 57060 23112 57112 23118
rect 57060 23054 57112 23060
rect 57072 22778 57100 23054
rect 57164 22930 57192 24550
rect 57164 22902 57284 22930
rect 57060 22772 57112 22778
rect 57060 22714 57112 22720
rect 57152 22636 57204 22642
rect 57152 22578 57204 22584
rect 57060 22094 57112 22098
rect 56980 22092 57112 22094
rect 56980 22066 57060 22092
rect 57060 22034 57112 22040
rect 56692 21684 56744 21690
rect 56692 21626 56744 21632
rect 56704 21078 56732 21626
rect 56968 21548 57020 21554
rect 56968 21490 57020 21496
rect 56324 21072 56376 21078
rect 56324 21014 56376 21020
rect 56692 21072 56744 21078
rect 56692 21014 56744 21020
rect 56232 20936 56284 20942
rect 56232 20878 56284 20884
rect 56784 20936 56836 20942
rect 56836 20884 56916 20890
rect 56784 20878 56916 20884
rect 56600 20868 56652 20874
rect 56600 20810 56652 20816
rect 56692 20868 56744 20874
rect 56796 20862 56916 20878
rect 56980 20874 57008 21490
rect 56692 20810 56744 20816
rect 56232 20800 56284 20806
rect 56232 20742 56284 20748
rect 56244 19514 56272 20742
rect 56508 19712 56560 19718
rect 56508 19654 56560 19660
rect 56232 19508 56284 19514
rect 56232 19450 56284 19456
rect 56324 17604 56376 17610
rect 56324 17546 56376 17552
rect 56336 17270 56364 17546
rect 56324 17264 56376 17270
rect 56324 17206 56376 17212
rect 56140 17128 56192 17134
rect 56140 17070 56192 17076
rect 56152 16998 56180 17070
rect 56324 17060 56376 17066
rect 56324 17002 56376 17008
rect 56140 16992 56192 16998
rect 56140 16934 56192 16940
rect 55876 16546 56088 16574
rect 55496 14408 55548 14414
rect 55496 14350 55548 14356
rect 55508 13938 55536 14350
rect 55496 13932 55548 13938
rect 55496 13874 55548 13880
rect 55404 13728 55456 13734
rect 55404 13670 55456 13676
rect 55416 12986 55444 13670
rect 55404 12980 55456 12986
rect 55404 12922 55456 12928
rect 55588 10124 55640 10130
rect 55588 10066 55640 10072
rect 55312 9580 55364 9586
rect 55312 9522 55364 9528
rect 55324 8974 55352 9522
rect 55600 9518 55628 10066
rect 55588 9512 55640 9518
rect 55588 9454 55640 9460
rect 55600 9042 55628 9454
rect 55588 9036 55640 9042
rect 55588 8978 55640 8984
rect 55312 8968 55364 8974
rect 55312 8910 55364 8916
rect 55772 7200 55824 7206
rect 55772 7142 55824 7148
rect 55232 6886 55444 6914
rect 50988 2644 51120 2650
rect 51040 2638 51120 2644
rect 51172 2644 51224 2650
rect 50988 2586 51040 2592
rect 51172 2586 51224 2592
rect 52368 2644 52420 2650
rect 52368 2586 52420 2592
rect 51184 2446 51212 2586
rect 52564 2582 52592 6886
rect 54588 6798 54616 6886
rect 54576 6792 54628 6798
rect 54576 6734 54628 6740
rect 54944 6792 54996 6798
rect 54944 6734 54996 6740
rect 54588 6322 54616 6734
rect 53564 6316 53616 6322
rect 53564 6258 53616 6264
rect 54576 6316 54628 6322
rect 54576 6258 54628 6264
rect 53576 6118 53604 6258
rect 54956 6254 54984 6734
rect 55416 6730 55444 6886
rect 55496 6792 55548 6798
rect 55496 6734 55548 6740
rect 55404 6724 55456 6730
rect 55404 6666 55456 6672
rect 55508 6458 55536 6734
rect 55496 6452 55548 6458
rect 55496 6394 55548 6400
rect 55784 6254 55812 7142
rect 54944 6248 54996 6254
rect 54944 6190 54996 6196
rect 55772 6248 55824 6254
rect 55772 6190 55824 6196
rect 53564 6112 53616 6118
rect 53564 6054 53616 6060
rect 53576 5710 53604 6054
rect 54956 5914 54984 6190
rect 55784 5914 55812 6190
rect 54944 5908 54996 5914
rect 54944 5850 54996 5856
rect 55772 5908 55824 5914
rect 55772 5850 55824 5856
rect 55784 5710 55812 5850
rect 53564 5704 53616 5710
rect 53564 5646 53616 5652
rect 55772 5704 55824 5710
rect 55772 5646 55824 5652
rect 53576 5574 53604 5646
rect 53564 5568 53616 5574
rect 53564 5510 53616 5516
rect 53576 4758 53604 5510
rect 55784 5030 55812 5646
rect 54576 5024 54628 5030
rect 54576 4966 54628 4972
rect 55772 5024 55824 5030
rect 55772 4966 55824 4972
rect 53564 4752 53616 4758
rect 53564 4694 53616 4700
rect 52736 2916 52788 2922
rect 52736 2858 52788 2864
rect 52552 2576 52604 2582
rect 52552 2518 52604 2524
rect 52748 2446 52776 2858
rect 51172 2440 51224 2446
rect 51172 2382 51224 2388
rect 52736 2440 52788 2446
rect 54208 2440 54260 2446
rect 52736 2382 52788 2388
rect 54128 2388 54208 2394
rect 54128 2382 54260 2388
rect 49792 2372 49844 2378
rect 49792 2314 49844 2320
rect 54128 2366 54248 2382
rect 48780 1964 48832 1970
rect 48780 1906 48832 1912
rect 49804 1766 49832 2314
rect 50160 2304 50212 2310
rect 50160 2246 50212 2252
rect 52184 2304 52236 2310
rect 52184 2246 52236 2252
rect 49792 1760 49844 1766
rect 49792 1702 49844 1708
rect 50172 1170 50200 2246
rect 50294 2204 50602 2224
rect 50294 2202 50300 2204
rect 50356 2202 50380 2204
rect 50436 2202 50460 2204
rect 50516 2202 50540 2204
rect 50596 2202 50602 2204
rect 50356 2150 50358 2202
rect 50538 2150 50540 2202
rect 50294 2148 50300 2150
rect 50356 2148 50380 2150
rect 50436 2148 50460 2150
rect 50516 2148 50540 2150
rect 50596 2148 50602 2150
rect 50294 2128 50602 2148
rect 50172 1142 50292 1170
rect 50264 800 50292 1142
rect 52196 800 52224 2246
rect 54128 800 54156 2366
rect 54588 2106 54616 4966
rect 55876 2650 55904 16546
rect 56152 16182 56180 16934
rect 56336 16590 56364 17002
rect 56232 16584 56284 16590
rect 56232 16526 56284 16532
rect 56324 16584 56376 16590
rect 56324 16526 56376 16532
rect 56140 16176 56192 16182
rect 56140 16118 56192 16124
rect 56244 15994 56272 16526
rect 56336 16114 56364 16526
rect 56324 16108 56376 16114
rect 56324 16050 56376 16056
rect 56244 15966 56364 15994
rect 56336 15910 56364 15966
rect 56324 15904 56376 15910
rect 56324 15846 56376 15852
rect 56336 14482 56364 15846
rect 56324 14476 56376 14482
rect 56324 14418 56376 14424
rect 56140 12776 56192 12782
rect 56140 12718 56192 12724
rect 56046 11792 56102 11801
rect 56046 11727 56048 11736
rect 56100 11727 56102 11736
rect 56048 11698 56100 11704
rect 55956 10056 56008 10062
rect 55956 9998 56008 10004
rect 55968 9586 55996 9998
rect 55956 9580 56008 9586
rect 55956 9522 56008 9528
rect 56152 9450 56180 12718
rect 56520 12238 56548 19654
rect 56612 19446 56640 20810
rect 56704 19854 56732 20810
rect 56888 19854 56916 20862
rect 56968 20868 57020 20874
rect 56968 20810 57020 20816
rect 57072 20602 57100 22034
rect 57164 22030 57192 22578
rect 57152 22024 57204 22030
rect 57152 21966 57204 21972
rect 57164 21690 57192 21966
rect 57152 21684 57204 21690
rect 57152 21626 57204 21632
rect 57060 20596 57112 20602
rect 57060 20538 57112 20544
rect 57256 20534 57284 22902
rect 57624 22094 57652 29174
rect 57716 29102 57744 29582
rect 57704 29096 57756 29102
rect 57704 29038 57756 29044
rect 57716 23050 57744 29038
rect 57808 28694 57836 36042
rect 58176 35834 58204 36110
rect 58164 35828 58216 35834
rect 58164 35770 58216 35776
rect 57886 35728 57942 35737
rect 57886 35663 57942 35672
rect 57900 35154 57928 35663
rect 58162 35456 58218 35465
rect 58162 35391 58218 35400
rect 57888 35148 57940 35154
rect 57888 35090 57940 35096
rect 58176 35086 58204 35391
rect 58164 35080 58216 35086
rect 58164 35022 58216 35028
rect 58176 34746 58204 35022
rect 58164 34740 58216 34746
rect 58164 34682 58216 34688
rect 58164 33516 58216 33522
rect 58164 33458 58216 33464
rect 58176 33425 58204 33458
rect 58162 33416 58218 33425
rect 58162 33351 58218 33360
rect 58176 33114 58204 33351
rect 58164 33108 58216 33114
rect 58164 33050 58216 33056
rect 57888 31816 57940 31822
rect 57888 31758 57940 31764
rect 57900 31385 57928 31758
rect 57886 31376 57942 31385
rect 57886 31311 57942 31320
rect 57888 29640 57940 29646
rect 57888 29582 57940 29588
rect 57900 29170 57928 29582
rect 58162 29336 58218 29345
rect 58162 29271 58218 29280
rect 58176 29170 58204 29271
rect 57888 29164 57940 29170
rect 57888 29106 57940 29112
rect 58164 29164 58216 29170
rect 58164 29106 58216 29112
rect 57900 28762 57928 29106
rect 58176 28762 58204 29106
rect 57888 28756 57940 28762
rect 57888 28698 57940 28704
rect 58164 28756 58216 28762
rect 58164 28698 58216 28704
rect 57796 28688 57848 28694
rect 57796 28630 57848 28636
rect 57980 28416 58032 28422
rect 57980 28358 58032 28364
rect 57992 27878 58020 28358
rect 57980 27872 58032 27878
rect 57980 27814 58032 27820
rect 57888 26784 57940 26790
rect 57888 26726 57940 26732
rect 57900 25294 57928 26726
rect 57888 25288 57940 25294
rect 57888 25230 57940 25236
rect 57992 24954 58020 27814
rect 58164 27464 58216 27470
rect 58164 27406 58216 27412
rect 58176 27305 58204 27406
rect 58162 27296 58218 27305
rect 58162 27231 58218 27240
rect 58176 27130 58204 27231
rect 58164 27124 58216 27130
rect 58164 27066 58216 27072
rect 58070 25256 58126 25265
rect 58070 25191 58126 25200
rect 58084 25158 58112 25191
rect 58072 25152 58124 25158
rect 58072 25094 58124 25100
rect 57980 24948 58032 24954
rect 57980 24890 58032 24896
rect 57900 24818 58112 24834
rect 57888 24812 58112 24818
rect 57940 24806 58112 24812
rect 57888 24754 57940 24760
rect 57888 24268 57940 24274
rect 57888 24210 57940 24216
rect 57900 23526 57928 24210
rect 57888 23520 57940 23526
rect 57888 23462 57940 23468
rect 57900 23225 57928 23462
rect 57886 23216 57942 23225
rect 57886 23151 57942 23160
rect 57704 23044 57756 23050
rect 57704 22986 57756 22992
rect 57624 22066 57744 22094
rect 57336 21548 57388 21554
rect 57336 21490 57388 21496
rect 57244 20528 57296 20534
rect 57244 20470 57296 20476
rect 56968 20460 57020 20466
rect 56968 20402 57020 20408
rect 56692 19848 56744 19854
rect 56692 19790 56744 19796
rect 56876 19848 56928 19854
rect 56876 19790 56928 19796
rect 56600 19440 56652 19446
rect 56600 19382 56652 19388
rect 56612 19258 56640 19382
rect 56888 19378 56916 19790
rect 56876 19372 56928 19378
rect 56876 19314 56928 19320
rect 56612 19230 56732 19258
rect 56600 19168 56652 19174
rect 56600 19110 56652 19116
rect 56612 18766 56640 19110
rect 56600 18760 56652 18766
rect 56600 18702 56652 18708
rect 56612 18290 56640 18702
rect 56704 18698 56732 19230
rect 56784 18828 56836 18834
rect 56784 18770 56836 18776
rect 56692 18692 56744 18698
rect 56692 18634 56744 18640
rect 56704 18426 56732 18634
rect 56692 18420 56744 18426
rect 56692 18362 56744 18368
rect 56796 18290 56824 18770
rect 56600 18284 56652 18290
rect 56600 18226 56652 18232
rect 56784 18284 56836 18290
rect 56784 18226 56836 18232
rect 56692 17672 56744 17678
rect 56692 17614 56744 17620
rect 56704 15162 56732 17614
rect 56796 17270 56824 18226
rect 56980 17882 57008 20402
rect 57348 19922 57376 21490
rect 57716 21010 57744 22066
rect 57980 21956 58032 21962
rect 57980 21898 58032 21904
rect 57992 21690 58020 21898
rect 57980 21684 58032 21690
rect 57980 21626 58032 21632
rect 58084 21570 58112 24806
rect 57992 21542 58112 21570
rect 57704 21004 57756 21010
rect 57704 20946 57756 20952
rect 57336 19916 57388 19922
rect 57336 19858 57388 19864
rect 57152 19848 57204 19854
rect 57152 19790 57204 19796
rect 57164 19174 57192 19790
rect 57244 19508 57296 19514
rect 57244 19450 57296 19456
rect 57152 19168 57204 19174
rect 57152 19110 57204 19116
rect 57060 18216 57112 18222
rect 57060 18158 57112 18164
rect 56968 17876 57020 17882
rect 56968 17818 57020 17824
rect 57072 17746 57100 18158
rect 57060 17740 57112 17746
rect 57060 17682 57112 17688
rect 56968 17672 57020 17678
rect 56968 17614 57020 17620
rect 56784 17264 56836 17270
rect 56784 17206 56836 17212
rect 56784 15904 56836 15910
rect 56784 15846 56836 15852
rect 56796 15570 56824 15846
rect 56784 15564 56836 15570
rect 56784 15506 56836 15512
rect 56692 15156 56744 15162
rect 56692 15098 56744 15104
rect 56796 15026 56824 15506
rect 56784 15020 56836 15026
rect 56784 14962 56836 14968
rect 56600 13932 56652 13938
rect 56600 13874 56652 13880
rect 56612 13530 56640 13874
rect 56876 13864 56928 13870
rect 56876 13806 56928 13812
rect 56784 13728 56836 13734
rect 56784 13670 56836 13676
rect 56600 13524 56652 13530
rect 56600 13466 56652 13472
rect 56612 12850 56640 13466
rect 56796 13326 56824 13670
rect 56888 13394 56916 13806
rect 56876 13388 56928 13394
rect 56876 13330 56928 13336
rect 56784 13320 56836 13326
rect 56784 13262 56836 13268
rect 56796 12918 56824 13262
rect 56784 12912 56836 12918
rect 56784 12854 56836 12860
rect 56888 12850 56916 13330
rect 56600 12844 56652 12850
rect 56600 12786 56652 12792
rect 56876 12844 56928 12850
rect 56876 12786 56928 12792
rect 56508 12232 56560 12238
rect 56508 12174 56560 12180
rect 56232 12164 56284 12170
rect 56232 12106 56284 12112
rect 56244 11830 56272 12106
rect 56600 12096 56652 12102
rect 56600 12038 56652 12044
rect 56232 11824 56284 11830
rect 56232 11766 56284 11772
rect 56244 10810 56272 11766
rect 56612 11694 56640 12038
rect 56692 11756 56744 11762
rect 56692 11698 56744 11704
rect 56600 11688 56652 11694
rect 56600 11630 56652 11636
rect 56508 11144 56560 11150
rect 56508 11086 56560 11092
rect 56232 10804 56284 10810
rect 56232 10746 56284 10752
rect 56520 10470 56548 11086
rect 56508 10464 56560 10470
rect 56508 10406 56560 10412
rect 56520 10130 56548 10406
rect 56704 10266 56732 11698
rect 56980 11286 57008 17614
rect 57152 17196 57204 17202
rect 57152 17138 57204 17144
rect 57164 16658 57192 17138
rect 57152 16652 57204 16658
rect 57152 16594 57204 16600
rect 57164 16114 57192 16594
rect 57152 16108 57204 16114
rect 57152 16050 57204 16056
rect 57060 15496 57112 15502
rect 57060 15438 57112 15444
rect 57072 15026 57100 15438
rect 57060 15020 57112 15026
rect 57060 14962 57112 14968
rect 57256 12458 57284 19450
rect 57348 18834 57376 19858
rect 57888 19372 57940 19378
rect 57888 19314 57940 19320
rect 57704 19168 57756 19174
rect 57704 19110 57756 19116
rect 57336 18828 57388 18834
rect 57336 18770 57388 18776
rect 57716 18290 57744 19110
rect 57900 18766 57928 19314
rect 57888 18760 57940 18766
rect 57888 18702 57940 18708
rect 57796 18624 57848 18630
rect 57796 18566 57848 18572
rect 57704 18284 57756 18290
rect 57704 18226 57756 18232
rect 57716 16574 57744 18226
rect 57808 18222 57836 18566
rect 57796 18216 57848 18222
rect 57796 18158 57848 18164
rect 57624 16546 57744 16574
rect 57428 15156 57480 15162
rect 57428 15098 57480 15104
rect 57336 14408 57388 14414
rect 57336 14350 57388 14356
rect 57164 12430 57284 12458
rect 57164 12238 57192 12430
rect 57152 12232 57204 12238
rect 57152 12174 57204 12180
rect 57060 12096 57112 12102
rect 57060 12038 57112 12044
rect 56968 11280 57020 11286
rect 56968 11222 57020 11228
rect 56980 11098 57008 11222
rect 56796 11070 57008 11098
rect 56796 10674 56824 11070
rect 56968 11008 57020 11014
rect 56968 10950 57020 10956
rect 56876 10736 56928 10742
rect 56980 10724 57008 10950
rect 56928 10696 57008 10724
rect 56876 10678 56928 10684
rect 56784 10668 56836 10674
rect 56784 10610 56836 10616
rect 56692 10260 56744 10266
rect 56692 10202 56744 10208
rect 56508 10124 56560 10130
rect 56508 10066 56560 10072
rect 56232 9512 56284 9518
rect 56232 9454 56284 9460
rect 56140 9444 56192 9450
rect 56140 9386 56192 9392
rect 56152 9042 56180 9386
rect 56140 9036 56192 9042
rect 56140 8978 56192 8984
rect 56244 8974 56272 9454
rect 56796 9042 56824 10610
rect 56980 10062 57008 10696
rect 56968 10056 57020 10062
rect 56968 9998 57020 10004
rect 56784 9036 56836 9042
rect 56784 8978 56836 8984
rect 56232 8968 56284 8974
rect 56232 8910 56284 8916
rect 56244 8634 56272 8910
rect 56232 8628 56284 8634
rect 56232 8570 56284 8576
rect 57072 8498 57100 12038
rect 57164 11762 57192 12174
rect 57152 11756 57204 11762
rect 57152 11698 57204 11704
rect 57152 9920 57204 9926
rect 57152 9862 57204 9868
rect 57060 8492 57112 8498
rect 57060 8434 57112 8440
rect 57164 8430 57192 9862
rect 56140 8424 56192 8430
rect 56140 8366 56192 8372
rect 57152 8424 57204 8430
rect 57152 8366 57204 8372
rect 56152 6322 56180 8366
rect 56232 7404 56284 7410
rect 56232 7346 56284 7352
rect 56244 6798 56272 7346
rect 57348 7342 57376 14350
rect 57440 11150 57468 15098
rect 57624 11218 57652 16546
rect 57704 16448 57756 16454
rect 57704 16390 57756 16396
rect 57612 11212 57664 11218
rect 57612 11154 57664 11160
rect 57428 11144 57480 11150
rect 57428 11086 57480 11092
rect 57440 10674 57468 11086
rect 57428 10668 57480 10674
rect 57428 10610 57480 10616
rect 57612 10668 57664 10674
rect 57612 10610 57664 10616
rect 57624 9926 57652 10610
rect 57612 9920 57664 9926
rect 57612 9862 57664 9868
rect 57518 7848 57574 7857
rect 57518 7783 57520 7792
rect 57572 7783 57574 7792
rect 57520 7754 57572 7760
rect 57060 7336 57112 7342
rect 57060 7278 57112 7284
rect 57336 7336 57388 7342
rect 57336 7278 57388 7284
rect 56692 6860 56744 6866
rect 56692 6802 56744 6808
rect 56232 6792 56284 6798
rect 56232 6734 56284 6740
rect 56140 6316 56192 6322
rect 56140 6258 56192 6264
rect 56152 5710 56180 6258
rect 56244 6186 56272 6734
rect 56704 6322 56732 6802
rect 56784 6792 56836 6798
rect 56782 6760 56784 6769
rect 56836 6760 56838 6769
rect 56782 6695 56838 6704
rect 56876 6724 56928 6730
rect 56876 6666 56928 6672
rect 56888 6458 56916 6666
rect 57072 6458 57100 7278
rect 56876 6452 56928 6458
rect 56876 6394 56928 6400
rect 57060 6452 57112 6458
rect 57060 6394 57112 6400
rect 56692 6316 56744 6322
rect 56692 6258 56744 6264
rect 56232 6180 56284 6186
rect 56232 6122 56284 6128
rect 56140 5704 56192 5710
rect 56140 5646 56192 5652
rect 56704 5370 56732 6258
rect 56888 5778 56916 6394
rect 56876 5772 56928 5778
rect 56876 5714 56928 5720
rect 56692 5364 56744 5370
rect 56692 5306 56744 5312
rect 56704 5166 56732 5306
rect 56888 5234 56916 5714
rect 56876 5228 56928 5234
rect 56876 5170 56928 5176
rect 56692 5160 56744 5166
rect 56692 5102 56744 5108
rect 57624 3466 57652 9862
rect 57716 5302 57744 16390
rect 57900 15570 57928 18702
rect 57992 18426 58020 21542
rect 58164 20936 58216 20942
rect 58164 20878 58216 20884
rect 58176 20534 58204 20878
rect 58164 20528 58216 20534
rect 58162 20496 58164 20505
rect 58216 20496 58218 20505
rect 58162 20431 58218 20440
rect 58070 18456 58126 18465
rect 57980 18420 58032 18426
rect 58070 18391 58126 18400
rect 57980 18362 58032 18368
rect 58084 17678 58112 18391
rect 58072 17672 58124 17678
rect 58072 17614 58124 17620
rect 58084 17338 58112 17614
rect 58072 17332 58124 17338
rect 58072 17274 58124 17280
rect 58164 16584 58216 16590
rect 58164 16526 58216 16532
rect 58176 16425 58204 16526
rect 58162 16416 58218 16425
rect 58162 16351 58218 16360
rect 58176 16250 58204 16351
rect 58164 16244 58216 16250
rect 58164 16186 58216 16192
rect 57888 15564 57940 15570
rect 57888 15506 57940 15512
rect 57888 15020 57940 15026
rect 57888 14962 57940 14968
rect 57900 14074 57928 14962
rect 58070 14376 58126 14385
rect 58070 14311 58126 14320
rect 58084 14278 58112 14311
rect 58072 14272 58124 14278
rect 58072 14214 58124 14220
rect 57888 14068 57940 14074
rect 57888 14010 57940 14016
rect 57888 13932 57940 13938
rect 57888 13874 57940 13880
rect 57900 13530 57928 13874
rect 57888 13524 57940 13530
rect 57888 13466 57940 13472
rect 57796 13456 57848 13462
rect 57796 13398 57848 13404
rect 57808 12306 57836 13398
rect 58162 12336 58218 12345
rect 57796 12300 57848 12306
rect 58162 12271 58218 12280
rect 57796 12242 57848 12248
rect 58176 12238 58204 12271
rect 58164 12232 58216 12238
rect 58164 12174 58216 12180
rect 58176 11898 58204 12174
rect 58164 11892 58216 11898
rect 58164 11834 58216 11840
rect 58072 10464 58124 10470
rect 58072 10406 58124 10412
rect 58084 10305 58112 10406
rect 58070 10296 58126 10305
rect 58070 10231 58126 10240
rect 58070 8256 58126 8265
rect 58070 8191 58126 8200
rect 58084 7886 58112 8191
rect 58072 7880 58124 7886
rect 58072 7822 58124 7828
rect 58084 7546 58112 7822
rect 58072 7540 58124 7546
rect 58072 7482 58124 7488
rect 57796 6316 57848 6322
rect 57796 6258 57848 6264
rect 57808 5914 57836 6258
rect 58070 6216 58126 6225
rect 58070 6151 58072 6160
rect 58124 6151 58126 6160
rect 58072 6122 58124 6128
rect 57796 5908 57848 5914
rect 57796 5850 57848 5856
rect 57704 5296 57756 5302
rect 57704 5238 57756 5244
rect 57888 5024 57940 5030
rect 57888 4966 57940 4972
rect 57612 3460 57664 3466
rect 57612 3402 57664 3408
rect 57152 3392 57204 3398
rect 57152 3334 57204 3340
rect 57164 3194 57192 3334
rect 57152 3188 57204 3194
rect 57152 3130 57204 3136
rect 56048 2848 56100 2854
rect 56048 2790 56100 2796
rect 57244 2848 57296 2854
rect 57244 2790 57296 2796
rect 55864 2644 55916 2650
rect 55864 2586 55916 2592
rect 56060 2446 56088 2790
rect 56048 2440 56100 2446
rect 56048 2382 56100 2388
rect 54576 2100 54628 2106
rect 54576 2042 54628 2048
rect 56060 800 56088 2382
rect 57256 2378 57284 2790
rect 57900 2446 57928 4966
rect 58072 3936 58124 3942
rect 58072 3878 58124 3884
rect 58084 3534 58112 3878
rect 58072 3528 58124 3534
rect 58070 3496 58072 3505
rect 58124 3496 58126 3505
rect 58070 3431 58126 3440
rect 59912 2848 59964 2854
rect 59912 2790 59964 2796
rect 57888 2440 57940 2446
rect 57888 2382 57940 2388
rect 57244 2372 57296 2378
rect 57244 2314 57296 2320
rect 57256 1465 57284 2314
rect 57980 2304 58032 2310
rect 57980 2246 58032 2252
rect 57242 1456 57298 1465
rect 57242 1391 57298 1400
rect 57992 800 58020 2246
rect 59924 800 59952 2790
rect 25884 734 26188 762
rect 27710 0 27766 800
rect 29642 0 29698 800
rect 31574 0 31630 800
rect 34150 0 34206 800
rect 36082 0 36138 800
rect 38014 0 38070 800
rect 39946 0 40002 800
rect 41878 0 41934 800
rect 43810 0 43866 800
rect 45742 0 45798 800
rect 47674 0 47730 800
rect 50250 0 50306 800
rect 52182 0 52238 800
rect 54114 0 54170 800
rect 56046 0 56102 800
rect 57978 0 58034 800
rect 59910 0 59966 800
<< via2 >>
rect 1490 38120 1546 38176
rect 4220 37562 4276 37564
rect 4300 37562 4356 37564
rect 4380 37562 4436 37564
rect 4460 37562 4516 37564
rect 4220 37510 4266 37562
rect 4266 37510 4276 37562
rect 4300 37510 4330 37562
rect 4330 37510 4342 37562
rect 4342 37510 4356 37562
rect 4380 37510 4394 37562
rect 4394 37510 4406 37562
rect 4406 37510 4436 37562
rect 4460 37510 4470 37562
rect 4470 37510 4516 37562
rect 4220 37508 4276 37510
rect 4300 37508 4356 37510
rect 4380 37508 4436 37510
rect 4460 37508 4516 37510
rect 1490 36080 1546 36136
rect 1582 33360 1638 33416
rect 1582 31356 1584 31376
rect 1584 31356 1636 31376
rect 1636 31356 1638 31376
rect 1582 31320 1638 31356
rect 1490 29280 1546 29336
rect 1398 21140 1454 21176
rect 1398 21120 1400 21140
rect 1400 21120 1452 21140
rect 1452 21120 1454 21140
rect 1398 19080 1454 19136
rect 1398 14356 1400 14376
rect 1400 14356 1452 14376
rect 1452 14356 1454 14376
rect 1398 14320 1454 14356
rect 1858 27240 1914 27296
rect 1858 25220 1914 25256
rect 1858 25200 1860 25220
rect 1860 25200 1912 25220
rect 1912 25200 1914 25220
rect 1858 23160 1914 23216
rect 2042 23044 2098 23080
rect 2042 23024 2044 23044
rect 2044 23024 2096 23044
rect 2096 23024 2098 23044
rect 3238 31320 3294 31376
rect 1858 16360 1914 16416
rect 2686 18808 2742 18864
rect 1398 12316 1400 12336
rect 1400 12316 1452 12336
rect 1452 12316 1454 12336
rect 1398 12280 1454 12316
rect 1398 10260 1454 10296
rect 1398 10240 1400 10260
rect 1400 10240 1452 10260
rect 1452 10240 1454 10260
rect 4220 36474 4276 36476
rect 4300 36474 4356 36476
rect 4380 36474 4436 36476
rect 4460 36474 4516 36476
rect 4220 36422 4266 36474
rect 4266 36422 4276 36474
rect 4300 36422 4330 36474
rect 4330 36422 4342 36474
rect 4342 36422 4356 36474
rect 4380 36422 4394 36474
rect 4394 36422 4406 36474
rect 4406 36422 4436 36474
rect 4460 36422 4470 36474
rect 4470 36422 4516 36474
rect 4220 36420 4276 36422
rect 4300 36420 4356 36422
rect 4380 36420 4436 36422
rect 4460 36420 4516 36422
rect 4220 35386 4276 35388
rect 4300 35386 4356 35388
rect 4380 35386 4436 35388
rect 4460 35386 4516 35388
rect 4220 35334 4266 35386
rect 4266 35334 4276 35386
rect 4300 35334 4330 35386
rect 4330 35334 4342 35386
rect 4342 35334 4356 35386
rect 4380 35334 4394 35386
rect 4394 35334 4406 35386
rect 4406 35334 4436 35386
rect 4460 35334 4470 35386
rect 4470 35334 4516 35386
rect 4220 35332 4276 35334
rect 4300 35332 4356 35334
rect 4380 35332 4436 35334
rect 4460 35332 4516 35334
rect 4220 34298 4276 34300
rect 4300 34298 4356 34300
rect 4380 34298 4436 34300
rect 4460 34298 4516 34300
rect 4220 34246 4266 34298
rect 4266 34246 4276 34298
rect 4300 34246 4330 34298
rect 4330 34246 4342 34298
rect 4342 34246 4356 34298
rect 4380 34246 4394 34298
rect 4394 34246 4406 34298
rect 4406 34246 4436 34298
rect 4460 34246 4470 34298
rect 4470 34246 4516 34298
rect 4220 34244 4276 34246
rect 4300 34244 4356 34246
rect 4380 34244 4436 34246
rect 4460 34244 4516 34246
rect 4220 33210 4276 33212
rect 4300 33210 4356 33212
rect 4380 33210 4436 33212
rect 4460 33210 4516 33212
rect 4220 33158 4266 33210
rect 4266 33158 4276 33210
rect 4300 33158 4330 33210
rect 4330 33158 4342 33210
rect 4342 33158 4356 33210
rect 4380 33158 4394 33210
rect 4394 33158 4406 33210
rect 4406 33158 4436 33210
rect 4460 33158 4470 33210
rect 4470 33158 4516 33210
rect 4220 33156 4276 33158
rect 4300 33156 4356 33158
rect 4380 33156 4436 33158
rect 4460 33156 4516 33158
rect 4220 32122 4276 32124
rect 4300 32122 4356 32124
rect 4380 32122 4436 32124
rect 4460 32122 4516 32124
rect 4220 32070 4266 32122
rect 4266 32070 4276 32122
rect 4300 32070 4330 32122
rect 4330 32070 4342 32122
rect 4342 32070 4356 32122
rect 4380 32070 4394 32122
rect 4394 32070 4406 32122
rect 4406 32070 4436 32122
rect 4460 32070 4470 32122
rect 4470 32070 4516 32122
rect 4220 32068 4276 32070
rect 4300 32068 4356 32070
rect 4380 32068 4436 32070
rect 4460 32068 4516 32070
rect 4220 31034 4276 31036
rect 4300 31034 4356 31036
rect 4380 31034 4436 31036
rect 4460 31034 4516 31036
rect 4220 30982 4266 31034
rect 4266 30982 4276 31034
rect 4300 30982 4330 31034
rect 4330 30982 4342 31034
rect 4342 30982 4356 31034
rect 4380 30982 4394 31034
rect 4394 30982 4406 31034
rect 4406 30982 4436 31034
rect 4460 30982 4470 31034
rect 4470 30982 4516 31034
rect 4220 30980 4276 30982
rect 4300 30980 4356 30982
rect 4380 30980 4436 30982
rect 4460 30980 4516 30982
rect 4220 29946 4276 29948
rect 4300 29946 4356 29948
rect 4380 29946 4436 29948
rect 4460 29946 4516 29948
rect 4220 29894 4266 29946
rect 4266 29894 4276 29946
rect 4300 29894 4330 29946
rect 4330 29894 4342 29946
rect 4342 29894 4356 29946
rect 4380 29894 4394 29946
rect 4394 29894 4406 29946
rect 4406 29894 4436 29946
rect 4460 29894 4470 29946
rect 4470 29894 4516 29946
rect 4220 29892 4276 29894
rect 4300 29892 4356 29894
rect 4380 29892 4436 29894
rect 4460 29892 4516 29894
rect 4220 28858 4276 28860
rect 4300 28858 4356 28860
rect 4380 28858 4436 28860
rect 4460 28858 4516 28860
rect 4220 28806 4266 28858
rect 4266 28806 4276 28858
rect 4300 28806 4330 28858
rect 4330 28806 4342 28858
rect 4342 28806 4356 28858
rect 4380 28806 4394 28858
rect 4394 28806 4406 28858
rect 4406 28806 4436 28858
rect 4460 28806 4470 28858
rect 4470 28806 4516 28858
rect 4220 28804 4276 28806
rect 4300 28804 4356 28806
rect 4380 28804 4436 28806
rect 4460 28804 4516 28806
rect 4220 27770 4276 27772
rect 4300 27770 4356 27772
rect 4380 27770 4436 27772
rect 4460 27770 4516 27772
rect 4220 27718 4266 27770
rect 4266 27718 4276 27770
rect 4300 27718 4330 27770
rect 4330 27718 4342 27770
rect 4342 27718 4356 27770
rect 4380 27718 4394 27770
rect 4394 27718 4406 27770
rect 4406 27718 4436 27770
rect 4460 27718 4470 27770
rect 4470 27718 4516 27770
rect 4220 27716 4276 27718
rect 4300 27716 4356 27718
rect 4380 27716 4436 27718
rect 4460 27716 4516 27718
rect 4220 26682 4276 26684
rect 4300 26682 4356 26684
rect 4380 26682 4436 26684
rect 4460 26682 4516 26684
rect 4220 26630 4266 26682
rect 4266 26630 4276 26682
rect 4300 26630 4330 26682
rect 4330 26630 4342 26682
rect 4342 26630 4356 26682
rect 4380 26630 4394 26682
rect 4394 26630 4406 26682
rect 4406 26630 4436 26682
rect 4460 26630 4470 26682
rect 4470 26630 4516 26682
rect 4220 26628 4276 26630
rect 4300 26628 4356 26630
rect 4380 26628 4436 26630
rect 4460 26628 4516 26630
rect 4220 25594 4276 25596
rect 4300 25594 4356 25596
rect 4380 25594 4436 25596
rect 4460 25594 4516 25596
rect 4220 25542 4266 25594
rect 4266 25542 4276 25594
rect 4300 25542 4330 25594
rect 4330 25542 4342 25594
rect 4342 25542 4356 25594
rect 4380 25542 4394 25594
rect 4394 25542 4406 25594
rect 4406 25542 4436 25594
rect 4460 25542 4470 25594
rect 4470 25542 4516 25594
rect 4220 25540 4276 25542
rect 4300 25540 4356 25542
rect 4380 25540 4436 25542
rect 4460 25540 4516 25542
rect 4220 24506 4276 24508
rect 4300 24506 4356 24508
rect 4380 24506 4436 24508
rect 4460 24506 4516 24508
rect 4220 24454 4266 24506
rect 4266 24454 4276 24506
rect 4300 24454 4330 24506
rect 4330 24454 4342 24506
rect 4342 24454 4356 24506
rect 4380 24454 4394 24506
rect 4394 24454 4406 24506
rect 4406 24454 4436 24506
rect 4460 24454 4470 24506
rect 4470 24454 4516 24506
rect 4220 24452 4276 24454
rect 4300 24452 4356 24454
rect 4380 24452 4436 24454
rect 4460 24452 4516 24454
rect 4220 23418 4276 23420
rect 4300 23418 4356 23420
rect 4380 23418 4436 23420
rect 4460 23418 4516 23420
rect 4220 23366 4266 23418
rect 4266 23366 4276 23418
rect 4300 23366 4330 23418
rect 4330 23366 4342 23418
rect 4342 23366 4356 23418
rect 4380 23366 4394 23418
rect 4394 23366 4406 23418
rect 4406 23366 4436 23418
rect 4460 23366 4470 23418
rect 4470 23366 4516 23418
rect 4220 23364 4276 23366
rect 4300 23364 4356 23366
rect 4380 23364 4436 23366
rect 4460 23364 4516 23366
rect 7470 25472 7526 25528
rect 4220 22330 4276 22332
rect 4300 22330 4356 22332
rect 4380 22330 4436 22332
rect 4460 22330 4516 22332
rect 4220 22278 4266 22330
rect 4266 22278 4276 22330
rect 4300 22278 4330 22330
rect 4330 22278 4342 22330
rect 4342 22278 4356 22330
rect 4380 22278 4394 22330
rect 4394 22278 4406 22330
rect 4406 22278 4436 22330
rect 4460 22278 4470 22330
rect 4470 22278 4516 22330
rect 4220 22276 4276 22278
rect 4300 22276 4356 22278
rect 4380 22276 4436 22278
rect 4460 22276 4516 22278
rect 4220 21242 4276 21244
rect 4300 21242 4356 21244
rect 4380 21242 4436 21244
rect 4460 21242 4516 21244
rect 4220 21190 4266 21242
rect 4266 21190 4276 21242
rect 4300 21190 4330 21242
rect 4330 21190 4342 21242
rect 4342 21190 4356 21242
rect 4380 21190 4394 21242
rect 4394 21190 4406 21242
rect 4406 21190 4436 21242
rect 4460 21190 4470 21242
rect 4470 21190 4516 21242
rect 4220 21188 4276 21190
rect 4300 21188 4356 21190
rect 4380 21188 4436 21190
rect 4460 21188 4516 21190
rect 4220 20154 4276 20156
rect 4300 20154 4356 20156
rect 4380 20154 4436 20156
rect 4460 20154 4516 20156
rect 4220 20102 4266 20154
rect 4266 20102 4276 20154
rect 4300 20102 4330 20154
rect 4330 20102 4342 20154
rect 4342 20102 4356 20154
rect 4380 20102 4394 20154
rect 4394 20102 4406 20154
rect 4406 20102 4436 20154
rect 4460 20102 4470 20154
rect 4470 20102 4516 20154
rect 4220 20100 4276 20102
rect 4300 20100 4356 20102
rect 4380 20100 4436 20102
rect 4460 20100 4516 20102
rect 4220 19066 4276 19068
rect 4300 19066 4356 19068
rect 4380 19066 4436 19068
rect 4460 19066 4516 19068
rect 4220 19014 4266 19066
rect 4266 19014 4276 19066
rect 4300 19014 4330 19066
rect 4330 19014 4342 19066
rect 4342 19014 4356 19066
rect 4380 19014 4394 19066
rect 4394 19014 4406 19066
rect 4406 19014 4436 19066
rect 4460 19014 4470 19066
rect 4470 19014 4516 19066
rect 4220 19012 4276 19014
rect 4300 19012 4356 19014
rect 4380 19012 4436 19014
rect 4460 19012 4516 19014
rect 4220 17978 4276 17980
rect 4300 17978 4356 17980
rect 4380 17978 4436 17980
rect 4460 17978 4516 17980
rect 4220 17926 4266 17978
rect 4266 17926 4276 17978
rect 4300 17926 4330 17978
rect 4330 17926 4342 17978
rect 4342 17926 4356 17978
rect 4380 17926 4394 17978
rect 4394 17926 4406 17978
rect 4406 17926 4436 17978
rect 4460 17926 4470 17978
rect 4470 17926 4516 17978
rect 4220 17924 4276 17926
rect 4300 17924 4356 17926
rect 4380 17924 4436 17926
rect 4460 17924 4516 17926
rect 4220 16890 4276 16892
rect 4300 16890 4356 16892
rect 4380 16890 4436 16892
rect 4460 16890 4516 16892
rect 4220 16838 4266 16890
rect 4266 16838 4276 16890
rect 4300 16838 4330 16890
rect 4330 16838 4342 16890
rect 4342 16838 4356 16890
rect 4380 16838 4394 16890
rect 4394 16838 4406 16890
rect 4406 16838 4436 16890
rect 4460 16838 4470 16890
rect 4470 16838 4516 16890
rect 4220 16836 4276 16838
rect 4300 16836 4356 16838
rect 4380 16836 4436 16838
rect 4460 16836 4516 16838
rect 4220 15802 4276 15804
rect 4300 15802 4356 15804
rect 4380 15802 4436 15804
rect 4460 15802 4516 15804
rect 4220 15750 4266 15802
rect 4266 15750 4276 15802
rect 4300 15750 4330 15802
rect 4330 15750 4342 15802
rect 4342 15750 4356 15802
rect 4380 15750 4394 15802
rect 4394 15750 4406 15802
rect 4406 15750 4436 15802
rect 4460 15750 4470 15802
rect 4470 15750 4516 15802
rect 4220 15748 4276 15750
rect 4300 15748 4356 15750
rect 4380 15748 4436 15750
rect 4460 15748 4516 15750
rect 4220 14714 4276 14716
rect 4300 14714 4356 14716
rect 4380 14714 4436 14716
rect 4460 14714 4516 14716
rect 4220 14662 4266 14714
rect 4266 14662 4276 14714
rect 4300 14662 4330 14714
rect 4330 14662 4342 14714
rect 4342 14662 4356 14714
rect 4380 14662 4394 14714
rect 4394 14662 4406 14714
rect 4406 14662 4436 14714
rect 4460 14662 4470 14714
rect 4470 14662 4516 14714
rect 4220 14660 4276 14662
rect 4300 14660 4356 14662
rect 4380 14660 4436 14662
rect 4460 14660 4516 14662
rect 1490 8200 1546 8256
rect 1582 6160 1638 6216
rect 1490 4120 1546 4176
rect 4220 13626 4276 13628
rect 4300 13626 4356 13628
rect 4380 13626 4436 13628
rect 4460 13626 4516 13628
rect 4220 13574 4266 13626
rect 4266 13574 4276 13626
rect 4300 13574 4330 13626
rect 4330 13574 4342 13626
rect 4342 13574 4356 13626
rect 4380 13574 4394 13626
rect 4394 13574 4406 13626
rect 4406 13574 4436 13626
rect 4460 13574 4470 13626
rect 4470 13574 4516 13626
rect 4220 13572 4276 13574
rect 4300 13572 4356 13574
rect 4380 13572 4436 13574
rect 4460 13572 4516 13574
rect 4220 12538 4276 12540
rect 4300 12538 4356 12540
rect 4380 12538 4436 12540
rect 4460 12538 4516 12540
rect 4220 12486 4266 12538
rect 4266 12486 4276 12538
rect 4300 12486 4330 12538
rect 4330 12486 4342 12538
rect 4342 12486 4356 12538
rect 4380 12486 4394 12538
rect 4394 12486 4406 12538
rect 4406 12486 4436 12538
rect 4460 12486 4470 12538
rect 4470 12486 4516 12538
rect 4220 12484 4276 12486
rect 4300 12484 4356 12486
rect 4380 12484 4436 12486
rect 4460 12484 4516 12486
rect 4220 11450 4276 11452
rect 4300 11450 4356 11452
rect 4380 11450 4436 11452
rect 4460 11450 4516 11452
rect 4220 11398 4266 11450
rect 4266 11398 4276 11450
rect 4300 11398 4330 11450
rect 4330 11398 4342 11450
rect 4342 11398 4356 11450
rect 4380 11398 4394 11450
rect 4394 11398 4406 11450
rect 4406 11398 4436 11450
rect 4460 11398 4470 11450
rect 4470 11398 4516 11450
rect 4220 11396 4276 11398
rect 4300 11396 4356 11398
rect 4380 11396 4436 11398
rect 4460 11396 4516 11398
rect 4220 10362 4276 10364
rect 4300 10362 4356 10364
rect 4380 10362 4436 10364
rect 4460 10362 4516 10364
rect 4220 10310 4266 10362
rect 4266 10310 4276 10362
rect 4300 10310 4330 10362
rect 4330 10310 4342 10362
rect 4342 10310 4356 10362
rect 4380 10310 4394 10362
rect 4394 10310 4406 10362
rect 4406 10310 4436 10362
rect 4460 10310 4470 10362
rect 4470 10310 4516 10362
rect 4220 10308 4276 10310
rect 4300 10308 4356 10310
rect 4380 10308 4436 10310
rect 4460 10308 4516 10310
rect 4220 9274 4276 9276
rect 4300 9274 4356 9276
rect 4380 9274 4436 9276
rect 4460 9274 4516 9276
rect 4220 9222 4266 9274
rect 4266 9222 4276 9274
rect 4300 9222 4330 9274
rect 4330 9222 4342 9274
rect 4342 9222 4356 9274
rect 4380 9222 4394 9274
rect 4394 9222 4406 9274
rect 4406 9222 4436 9274
rect 4460 9222 4470 9274
rect 4470 9222 4516 9274
rect 4220 9220 4276 9222
rect 4300 9220 4356 9222
rect 4380 9220 4436 9222
rect 4460 9220 4516 9222
rect 4220 8186 4276 8188
rect 4300 8186 4356 8188
rect 4380 8186 4436 8188
rect 4460 8186 4516 8188
rect 4220 8134 4266 8186
rect 4266 8134 4276 8186
rect 4300 8134 4330 8186
rect 4330 8134 4342 8186
rect 4342 8134 4356 8186
rect 4380 8134 4394 8186
rect 4394 8134 4406 8186
rect 4406 8134 4436 8186
rect 4460 8134 4470 8186
rect 4470 8134 4516 8186
rect 4220 8132 4276 8134
rect 4300 8132 4356 8134
rect 4380 8132 4436 8134
rect 4460 8132 4516 8134
rect 4220 7098 4276 7100
rect 4300 7098 4356 7100
rect 4380 7098 4436 7100
rect 4460 7098 4516 7100
rect 4220 7046 4266 7098
rect 4266 7046 4276 7098
rect 4300 7046 4330 7098
rect 4330 7046 4342 7098
rect 4342 7046 4356 7098
rect 4380 7046 4394 7098
rect 4394 7046 4406 7098
rect 4406 7046 4436 7098
rect 4460 7046 4470 7098
rect 4470 7046 4516 7098
rect 4220 7044 4276 7046
rect 4300 7044 4356 7046
rect 4380 7044 4436 7046
rect 4460 7044 4516 7046
rect 4220 6010 4276 6012
rect 4300 6010 4356 6012
rect 4380 6010 4436 6012
rect 4460 6010 4516 6012
rect 4220 5958 4266 6010
rect 4266 5958 4276 6010
rect 4300 5958 4330 6010
rect 4330 5958 4342 6010
rect 4342 5958 4356 6010
rect 4380 5958 4394 6010
rect 4394 5958 4406 6010
rect 4406 5958 4436 6010
rect 4460 5958 4470 6010
rect 4470 5958 4516 6010
rect 4220 5956 4276 5958
rect 4300 5956 4356 5958
rect 4380 5956 4436 5958
rect 4460 5956 4516 5958
rect 4220 4922 4276 4924
rect 4300 4922 4356 4924
rect 4380 4922 4436 4924
rect 4460 4922 4516 4924
rect 4220 4870 4266 4922
rect 4266 4870 4276 4922
rect 4300 4870 4330 4922
rect 4330 4870 4342 4922
rect 4342 4870 4356 4922
rect 4380 4870 4394 4922
rect 4394 4870 4406 4922
rect 4406 4870 4436 4922
rect 4460 4870 4470 4922
rect 4470 4870 4516 4922
rect 4220 4868 4276 4870
rect 4300 4868 4356 4870
rect 4380 4868 4436 4870
rect 4460 4868 4516 4870
rect 4220 3834 4276 3836
rect 4300 3834 4356 3836
rect 4380 3834 4436 3836
rect 4460 3834 4516 3836
rect 4220 3782 4266 3834
rect 4266 3782 4276 3834
rect 4300 3782 4330 3834
rect 4330 3782 4342 3834
rect 4342 3782 4356 3834
rect 4380 3782 4394 3834
rect 4394 3782 4406 3834
rect 4406 3782 4436 3834
rect 4460 3782 4470 3834
rect 4470 3782 4516 3834
rect 4220 3780 4276 3782
rect 4300 3780 4356 3782
rect 4380 3780 4436 3782
rect 4460 3780 4516 3782
rect 4220 2746 4276 2748
rect 4300 2746 4356 2748
rect 4380 2746 4436 2748
rect 4460 2746 4516 2748
rect 4220 2694 4266 2746
rect 4266 2694 4276 2746
rect 4300 2694 4330 2746
rect 4330 2694 4342 2746
rect 4342 2694 4356 2746
rect 4380 2694 4394 2746
rect 4394 2694 4406 2746
rect 4406 2694 4436 2746
rect 4460 2694 4470 2746
rect 4470 2694 4516 2746
rect 4220 2692 4276 2694
rect 4300 2692 4356 2694
rect 4380 2692 4436 2694
rect 4460 2692 4516 2694
rect 1398 2080 1454 2136
rect 7562 16108 7618 16144
rect 7562 16088 7564 16108
rect 7564 16088 7616 16108
rect 7616 16088 7618 16108
rect 5354 7792 5410 7848
rect 8390 24148 8392 24168
rect 8392 24148 8444 24168
rect 8444 24148 8446 24168
rect 8390 24112 8446 24148
rect 7102 11620 7158 11656
rect 7102 11600 7104 11620
rect 7104 11600 7156 11620
rect 7156 11600 7158 11620
rect 9586 35672 9642 35728
rect 8666 6704 8722 6760
rect 8942 24112 8998 24168
rect 10782 29008 10838 29064
rect 9770 21548 9826 21584
rect 9770 21528 9772 21548
rect 9772 21528 9824 21548
rect 9824 21528 9826 21548
rect 11058 29996 11060 30016
rect 11060 29996 11112 30016
rect 11112 29996 11114 30016
rect 11058 29960 11114 29996
rect 13082 29300 13138 29336
rect 13082 29280 13084 29300
rect 13084 29280 13136 29300
rect 13136 29280 13138 29300
rect 13634 29144 13690 29200
rect 10782 23432 10838 23488
rect 13910 29280 13966 29336
rect 14002 29008 14058 29064
rect 14922 29164 14978 29200
rect 14922 29144 14924 29164
rect 14924 29144 14976 29164
rect 14976 29144 14978 29164
rect 14646 29008 14702 29064
rect 10506 21392 10562 21448
rect 11058 21256 11114 21312
rect 10414 20476 10416 20496
rect 10416 20476 10468 20496
rect 10468 20476 10470 20496
rect 10414 20440 10470 20476
rect 16026 29280 16082 29336
rect 15658 27376 15714 27432
rect 14738 25200 14794 25256
rect 14738 24284 14740 24304
rect 14740 24284 14792 24304
rect 14792 24284 14794 24304
rect 14738 24248 14794 24284
rect 16210 29008 16266 29064
rect 15198 24812 15254 24848
rect 15198 24792 15200 24812
rect 15200 24792 15252 24812
rect 15252 24792 15254 24812
rect 15106 23432 15162 23488
rect 14462 22500 14518 22536
rect 14462 22480 14464 22500
rect 14464 22480 14516 22500
rect 14516 22480 14518 22500
rect 14186 22344 14242 22400
rect 15198 22616 15254 22672
rect 14094 21256 14150 21312
rect 10230 10104 10286 10160
rect 9862 9968 9918 10024
rect 9586 9424 9642 9480
rect 10046 8900 10102 8936
rect 10046 8880 10048 8900
rect 10048 8880 10100 8900
rect 10100 8880 10102 8900
rect 11886 16088 11942 16144
rect 12070 14728 12126 14784
rect 12622 14728 12678 14784
rect 10966 12552 11022 12608
rect 13082 20324 13138 20360
rect 13082 20304 13084 20324
rect 13084 20304 13136 20324
rect 13136 20304 13138 20324
rect 10874 10648 10930 10704
rect 10690 10548 10692 10568
rect 10692 10548 10744 10568
rect 10744 10548 10746 10568
rect 10690 10512 10746 10548
rect 13542 16768 13598 16824
rect 13726 15816 13782 15872
rect 13542 12416 13598 12472
rect 15474 22072 15530 22128
rect 15014 20984 15070 21040
rect 14922 18708 14924 18728
rect 14924 18708 14976 18728
rect 14976 18708 14978 18728
rect 14922 18672 14978 18708
rect 15566 17604 15622 17640
rect 15566 17584 15568 17604
rect 15568 17584 15620 17604
rect 15620 17584 15622 17604
rect 13726 7248 13782 7304
rect 15198 15408 15254 15464
rect 15566 14864 15622 14920
rect 19580 37018 19636 37020
rect 19660 37018 19716 37020
rect 19740 37018 19796 37020
rect 19820 37018 19876 37020
rect 19580 36966 19626 37018
rect 19626 36966 19636 37018
rect 19660 36966 19690 37018
rect 19690 36966 19702 37018
rect 19702 36966 19716 37018
rect 19740 36966 19754 37018
rect 19754 36966 19766 37018
rect 19766 36966 19796 37018
rect 19820 36966 19830 37018
rect 19830 36966 19876 37018
rect 19580 36964 19636 36966
rect 19660 36964 19716 36966
rect 19740 36964 19796 36966
rect 19820 36964 19876 36966
rect 19580 35930 19636 35932
rect 19660 35930 19716 35932
rect 19740 35930 19796 35932
rect 19820 35930 19876 35932
rect 19580 35878 19626 35930
rect 19626 35878 19636 35930
rect 19660 35878 19690 35930
rect 19690 35878 19702 35930
rect 19702 35878 19716 35930
rect 19740 35878 19754 35930
rect 19754 35878 19766 35930
rect 19766 35878 19796 35930
rect 19820 35878 19830 35930
rect 19830 35878 19876 35930
rect 19580 35876 19636 35878
rect 19660 35876 19716 35878
rect 19740 35876 19796 35878
rect 19820 35876 19876 35878
rect 19580 34842 19636 34844
rect 19660 34842 19716 34844
rect 19740 34842 19796 34844
rect 19820 34842 19876 34844
rect 19580 34790 19626 34842
rect 19626 34790 19636 34842
rect 19660 34790 19690 34842
rect 19690 34790 19702 34842
rect 19702 34790 19716 34842
rect 19740 34790 19754 34842
rect 19754 34790 19766 34842
rect 19766 34790 19796 34842
rect 19820 34790 19830 34842
rect 19830 34790 19876 34842
rect 19580 34788 19636 34790
rect 19660 34788 19716 34790
rect 19740 34788 19796 34790
rect 19820 34788 19876 34790
rect 19580 33754 19636 33756
rect 19660 33754 19716 33756
rect 19740 33754 19796 33756
rect 19820 33754 19876 33756
rect 19580 33702 19626 33754
rect 19626 33702 19636 33754
rect 19660 33702 19690 33754
rect 19690 33702 19702 33754
rect 19702 33702 19716 33754
rect 19740 33702 19754 33754
rect 19754 33702 19766 33754
rect 19766 33702 19796 33754
rect 19820 33702 19830 33754
rect 19830 33702 19876 33754
rect 19580 33700 19636 33702
rect 19660 33700 19716 33702
rect 19740 33700 19796 33702
rect 19820 33700 19876 33702
rect 18050 29960 18106 30016
rect 17038 22344 17094 22400
rect 16118 21256 16174 21312
rect 15750 20204 15752 20224
rect 15752 20204 15804 20224
rect 15804 20204 15806 20224
rect 15750 20168 15806 20204
rect 15934 19388 15936 19408
rect 15936 19388 15988 19408
rect 15988 19388 15990 19408
rect 15934 19352 15990 19388
rect 15842 15036 15844 15056
rect 15844 15036 15896 15056
rect 15896 15036 15898 15056
rect 15842 15000 15898 15036
rect 16302 20168 16358 20224
rect 16486 20848 16542 20904
rect 19580 32666 19636 32668
rect 19660 32666 19716 32668
rect 19740 32666 19796 32668
rect 19820 32666 19876 32668
rect 19580 32614 19626 32666
rect 19626 32614 19636 32666
rect 19660 32614 19690 32666
rect 19690 32614 19702 32666
rect 19702 32614 19716 32666
rect 19740 32614 19754 32666
rect 19754 32614 19766 32666
rect 19766 32614 19796 32666
rect 19820 32614 19830 32666
rect 19830 32614 19876 32666
rect 19580 32612 19636 32614
rect 19660 32612 19716 32614
rect 19740 32612 19796 32614
rect 19820 32612 19876 32614
rect 19580 31578 19636 31580
rect 19660 31578 19716 31580
rect 19740 31578 19796 31580
rect 19820 31578 19876 31580
rect 19580 31526 19626 31578
rect 19626 31526 19636 31578
rect 19660 31526 19690 31578
rect 19690 31526 19702 31578
rect 19702 31526 19716 31578
rect 19740 31526 19754 31578
rect 19754 31526 19766 31578
rect 19766 31526 19796 31578
rect 19820 31526 19830 31578
rect 19830 31526 19876 31578
rect 19580 31524 19636 31526
rect 19660 31524 19716 31526
rect 19740 31524 19796 31526
rect 19820 31524 19876 31526
rect 19580 30490 19636 30492
rect 19660 30490 19716 30492
rect 19740 30490 19796 30492
rect 19820 30490 19876 30492
rect 19580 30438 19626 30490
rect 19626 30438 19636 30490
rect 19660 30438 19690 30490
rect 19690 30438 19702 30490
rect 19702 30438 19716 30490
rect 19740 30438 19754 30490
rect 19754 30438 19766 30490
rect 19766 30438 19796 30490
rect 19820 30438 19830 30490
rect 19830 30438 19876 30490
rect 19580 30436 19636 30438
rect 19660 30436 19716 30438
rect 19740 30436 19796 30438
rect 19820 30436 19876 30438
rect 18694 26324 18696 26344
rect 18696 26324 18748 26344
rect 18748 26324 18750 26344
rect 18694 26288 18750 26324
rect 19580 29402 19636 29404
rect 19660 29402 19716 29404
rect 19740 29402 19796 29404
rect 19820 29402 19876 29404
rect 19580 29350 19626 29402
rect 19626 29350 19636 29402
rect 19660 29350 19690 29402
rect 19690 29350 19702 29402
rect 19702 29350 19716 29402
rect 19740 29350 19754 29402
rect 19754 29350 19766 29402
rect 19766 29350 19796 29402
rect 19820 29350 19830 29402
rect 19830 29350 19876 29402
rect 19580 29348 19636 29350
rect 19660 29348 19716 29350
rect 19740 29348 19796 29350
rect 19820 29348 19876 29350
rect 19338 29028 19394 29064
rect 19338 29008 19340 29028
rect 19340 29008 19392 29028
rect 19392 29008 19394 29028
rect 19338 27376 19394 27432
rect 15842 13932 15898 13968
rect 15842 13912 15844 13932
rect 15844 13912 15896 13932
rect 15896 13912 15898 13932
rect 16302 13948 16304 13968
rect 16304 13948 16356 13968
rect 16356 13948 16358 13968
rect 16302 13912 16358 13948
rect 16854 14900 16856 14920
rect 16856 14900 16908 14920
rect 16908 14900 16910 14920
rect 16854 14864 16910 14900
rect 16486 12688 16542 12744
rect 17222 12280 17278 12336
rect 17682 14884 17738 14920
rect 17682 14864 17684 14884
rect 17684 14864 17736 14884
rect 17736 14864 17738 14884
rect 17774 9152 17830 9208
rect 17498 9036 17554 9072
rect 17498 9016 17500 9036
rect 17500 9016 17552 9036
rect 17552 9016 17554 9036
rect 18050 3052 18106 3088
rect 18050 3032 18052 3052
rect 18052 3032 18104 3052
rect 18104 3032 18106 3052
rect 19580 28314 19636 28316
rect 19660 28314 19716 28316
rect 19740 28314 19796 28316
rect 19820 28314 19876 28316
rect 19580 28262 19626 28314
rect 19626 28262 19636 28314
rect 19660 28262 19690 28314
rect 19690 28262 19702 28314
rect 19702 28262 19716 28314
rect 19740 28262 19754 28314
rect 19754 28262 19766 28314
rect 19766 28262 19796 28314
rect 19820 28262 19830 28314
rect 19830 28262 19876 28314
rect 19580 28260 19636 28262
rect 19660 28260 19716 28262
rect 19740 28260 19796 28262
rect 19820 28260 19876 28262
rect 19580 27226 19636 27228
rect 19660 27226 19716 27228
rect 19740 27226 19796 27228
rect 19820 27226 19876 27228
rect 19580 27174 19626 27226
rect 19626 27174 19636 27226
rect 19660 27174 19690 27226
rect 19690 27174 19702 27226
rect 19702 27174 19716 27226
rect 19740 27174 19754 27226
rect 19754 27174 19766 27226
rect 19766 27174 19796 27226
rect 19820 27174 19830 27226
rect 19830 27174 19876 27226
rect 19580 27172 19636 27174
rect 19660 27172 19716 27174
rect 19740 27172 19796 27174
rect 19820 27172 19876 27174
rect 19706 26324 19708 26344
rect 19708 26324 19760 26344
rect 19760 26324 19762 26344
rect 19706 26288 19762 26324
rect 19580 26138 19636 26140
rect 19660 26138 19716 26140
rect 19740 26138 19796 26140
rect 19820 26138 19876 26140
rect 19580 26086 19626 26138
rect 19626 26086 19636 26138
rect 19660 26086 19690 26138
rect 19690 26086 19702 26138
rect 19702 26086 19716 26138
rect 19740 26086 19754 26138
rect 19754 26086 19766 26138
rect 19766 26086 19796 26138
rect 19820 26086 19830 26138
rect 19830 26086 19876 26138
rect 19580 26084 19636 26086
rect 19660 26084 19716 26086
rect 19740 26084 19796 26086
rect 19820 26084 19876 26086
rect 19580 25050 19636 25052
rect 19660 25050 19716 25052
rect 19740 25050 19796 25052
rect 19820 25050 19876 25052
rect 19580 24998 19626 25050
rect 19626 24998 19636 25050
rect 19660 24998 19690 25050
rect 19690 24998 19702 25050
rect 19702 24998 19716 25050
rect 19740 24998 19754 25050
rect 19754 24998 19766 25050
rect 19766 24998 19796 25050
rect 19820 24998 19830 25050
rect 19830 24998 19876 25050
rect 19580 24996 19636 24998
rect 19660 24996 19716 24998
rect 19740 24996 19796 24998
rect 19820 24996 19876 24998
rect 22006 27956 22008 27976
rect 22008 27956 22060 27976
rect 22060 27956 22062 27976
rect 22006 27920 22062 27956
rect 20810 26560 20866 26616
rect 19982 24792 20038 24848
rect 20350 24792 20406 24848
rect 19580 23962 19636 23964
rect 19660 23962 19716 23964
rect 19740 23962 19796 23964
rect 19820 23962 19876 23964
rect 19580 23910 19626 23962
rect 19626 23910 19636 23962
rect 19660 23910 19690 23962
rect 19690 23910 19702 23962
rect 19702 23910 19716 23962
rect 19740 23910 19754 23962
rect 19754 23910 19766 23962
rect 19766 23910 19796 23962
rect 19820 23910 19830 23962
rect 19830 23910 19876 23962
rect 19580 23908 19636 23910
rect 19660 23908 19716 23910
rect 19740 23908 19796 23910
rect 19820 23908 19876 23910
rect 19580 22874 19636 22876
rect 19660 22874 19716 22876
rect 19740 22874 19796 22876
rect 19820 22874 19876 22876
rect 19580 22822 19626 22874
rect 19626 22822 19636 22874
rect 19660 22822 19690 22874
rect 19690 22822 19702 22874
rect 19702 22822 19716 22874
rect 19740 22822 19754 22874
rect 19754 22822 19766 22874
rect 19766 22822 19796 22874
rect 19820 22822 19830 22874
rect 19830 22822 19876 22874
rect 19580 22820 19636 22822
rect 19660 22820 19716 22822
rect 19740 22820 19796 22822
rect 19820 22820 19876 22822
rect 20166 23976 20222 24032
rect 19338 21256 19394 21312
rect 19982 21800 20038 21856
rect 19580 21786 19636 21788
rect 19660 21786 19716 21788
rect 19740 21786 19796 21788
rect 19820 21786 19876 21788
rect 19580 21734 19626 21786
rect 19626 21734 19636 21786
rect 19660 21734 19690 21786
rect 19690 21734 19702 21786
rect 19702 21734 19716 21786
rect 19740 21734 19754 21786
rect 19754 21734 19766 21786
rect 19766 21734 19796 21786
rect 19820 21734 19830 21786
rect 19830 21734 19876 21786
rect 19580 21732 19636 21734
rect 19660 21732 19716 21734
rect 19740 21732 19796 21734
rect 19820 21732 19876 21734
rect 19580 20698 19636 20700
rect 19660 20698 19716 20700
rect 19740 20698 19796 20700
rect 19820 20698 19876 20700
rect 19580 20646 19626 20698
rect 19626 20646 19636 20698
rect 19660 20646 19690 20698
rect 19690 20646 19702 20698
rect 19702 20646 19716 20698
rect 19740 20646 19754 20698
rect 19754 20646 19766 20698
rect 19766 20646 19796 20698
rect 19820 20646 19830 20698
rect 19830 20646 19876 20698
rect 19580 20644 19636 20646
rect 19660 20644 19716 20646
rect 19740 20644 19796 20646
rect 19820 20644 19876 20646
rect 19580 19610 19636 19612
rect 19660 19610 19716 19612
rect 19740 19610 19796 19612
rect 19820 19610 19876 19612
rect 19580 19558 19626 19610
rect 19626 19558 19636 19610
rect 19660 19558 19690 19610
rect 19690 19558 19702 19610
rect 19702 19558 19716 19610
rect 19740 19558 19754 19610
rect 19754 19558 19766 19610
rect 19766 19558 19796 19610
rect 19820 19558 19830 19610
rect 19830 19558 19876 19610
rect 19580 19556 19636 19558
rect 19660 19556 19716 19558
rect 19740 19556 19796 19558
rect 19820 19556 19876 19558
rect 19580 18522 19636 18524
rect 19660 18522 19716 18524
rect 19740 18522 19796 18524
rect 19820 18522 19876 18524
rect 19580 18470 19626 18522
rect 19626 18470 19636 18522
rect 19660 18470 19690 18522
rect 19690 18470 19702 18522
rect 19702 18470 19716 18522
rect 19740 18470 19754 18522
rect 19754 18470 19766 18522
rect 19766 18470 19796 18522
rect 19820 18470 19830 18522
rect 19830 18470 19876 18522
rect 19580 18468 19636 18470
rect 19660 18468 19716 18470
rect 19740 18468 19796 18470
rect 19820 18468 19876 18470
rect 20350 21256 20406 21312
rect 20258 21120 20314 21176
rect 19580 17434 19636 17436
rect 19660 17434 19716 17436
rect 19740 17434 19796 17436
rect 19820 17434 19876 17436
rect 19580 17382 19626 17434
rect 19626 17382 19636 17434
rect 19660 17382 19690 17434
rect 19690 17382 19702 17434
rect 19702 17382 19716 17434
rect 19740 17382 19754 17434
rect 19754 17382 19766 17434
rect 19766 17382 19796 17434
rect 19820 17382 19830 17434
rect 19830 17382 19876 17434
rect 19580 17380 19636 17382
rect 19660 17380 19716 17382
rect 19740 17380 19796 17382
rect 19820 17380 19876 17382
rect 19706 16652 19762 16688
rect 19706 16632 19708 16652
rect 19708 16632 19760 16652
rect 19760 16632 19762 16652
rect 19580 16346 19636 16348
rect 19660 16346 19716 16348
rect 19740 16346 19796 16348
rect 19820 16346 19876 16348
rect 19580 16294 19626 16346
rect 19626 16294 19636 16346
rect 19660 16294 19690 16346
rect 19690 16294 19702 16346
rect 19702 16294 19716 16346
rect 19740 16294 19754 16346
rect 19754 16294 19766 16346
rect 19766 16294 19796 16346
rect 19820 16294 19830 16346
rect 19830 16294 19876 16346
rect 19580 16292 19636 16294
rect 19660 16292 19716 16294
rect 19740 16292 19796 16294
rect 19820 16292 19876 16294
rect 19338 14320 19394 14376
rect 19580 15258 19636 15260
rect 19660 15258 19716 15260
rect 19740 15258 19796 15260
rect 19820 15258 19876 15260
rect 19580 15206 19626 15258
rect 19626 15206 19636 15258
rect 19660 15206 19690 15258
rect 19690 15206 19702 15258
rect 19702 15206 19716 15258
rect 19740 15206 19754 15258
rect 19754 15206 19766 15258
rect 19766 15206 19796 15258
rect 19820 15206 19830 15258
rect 19830 15206 19876 15258
rect 19580 15204 19636 15206
rect 19660 15204 19716 15206
rect 19740 15204 19796 15206
rect 19820 15204 19876 15206
rect 19522 15000 19578 15056
rect 19580 14170 19636 14172
rect 19660 14170 19716 14172
rect 19740 14170 19796 14172
rect 19820 14170 19876 14172
rect 19580 14118 19626 14170
rect 19626 14118 19636 14170
rect 19660 14118 19690 14170
rect 19690 14118 19702 14170
rect 19702 14118 19716 14170
rect 19740 14118 19754 14170
rect 19754 14118 19766 14170
rect 19766 14118 19796 14170
rect 19820 14118 19830 14170
rect 19830 14118 19876 14170
rect 19580 14116 19636 14118
rect 19660 14116 19716 14118
rect 19740 14116 19796 14118
rect 19820 14116 19876 14118
rect 20810 17484 20812 17504
rect 20812 17484 20864 17504
rect 20864 17484 20866 17504
rect 20810 17448 20866 17484
rect 20626 15952 20682 16008
rect 21822 21256 21878 21312
rect 19982 13252 20038 13288
rect 19982 13232 19984 13252
rect 19984 13232 20036 13252
rect 20036 13232 20038 13252
rect 19580 13082 19636 13084
rect 19660 13082 19716 13084
rect 19740 13082 19796 13084
rect 19820 13082 19876 13084
rect 19580 13030 19626 13082
rect 19626 13030 19636 13082
rect 19660 13030 19690 13082
rect 19690 13030 19702 13082
rect 19702 13030 19716 13082
rect 19740 13030 19754 13082
rect 19754 13030 19766 13082
rect 19766 13030 19796 13082
rect 19820 13030 19830 13082
rect 19830 13030 19876 13082
rect 19580 13028 19636 13030
rect 19660 13028 19716 13030
rect 19740 13028 19796 13030
rect 19820 13028 19876 13030
rect 19580 11994 19636 11996
rect 19660 11994 19716 11996
rect 19740 11994 19796 11996
rect 19820 11994 19876 11996
rect 19580 11942 19626 11994
rect 19626 11942 19636 11994
rect 19660 11942 19690 11994
rect 19690 11942 19702 11994
rect 19702 11942 19716 11994
rect 19740 11942 19754 11994
rect 19754 11942 19766 11994
rect 19766 11942 19796 11994
rect 19820 11942 19830 11994
rect 19830 11942 19876 11994
rect 19580 11940 19636 11942
rect 19660 11940 19716 11942
rect 19740 11940 19796 11942
rect 19820 11940 19876 11942
rect 19580 10906 19636 10908
rect 19660 10906 19716 10908
rect 19740 10906 19796 10908
rect 19820 10906 19876 10908
rect 19580 10854 19626 10906
rect 19626 10854 19636 10906
rect 19660 10854 19690 10906
rect 19690 10854 19702 10906
rect 19702 10854 19716 10906
rect 19740 10854 19754 10906
rect 19754 10854 19766 10906
rect 19766 10854 19796 10906
rect 19820 10854 19830 10906
rect 19830 10854 19876 10906
rect 19580 10852 19636 10854
rect 19660 10852 19716 10854
rect 19740 10852 19796 10854
rect 19820 10852 19876 10854
rect 20718 15156 20774 15192
rect 20718 15136 20720 15156
rect 20720 15136 20772 15156
rect 20772 15136 20774 15156
rect 22098 21836 22100 21856
rect 22100 21836 22152 21856
rect 22152 21836 22154 21856
rect 22098 21800 22154 21836
rect 23294 29008 23350 29064
rect 22190 21256 22246 21312
rect 21086 15680 21142 15736
rect 20718 14728 20774 14784
rect 20902 13776 20958 13832
rect 20626 12164 20682 12200
rect 21822 13776 21878 13832
rect 21454 12280 21510 12336
rect 20626 12144 20628 12164
rect 20628 12144 20680 12164
rect 20680 12144 20682 12164
rect 19580 9818 19636 9820
rect 19660 9818 19716 9820
rect 19740 9818 19796 9820
rect 19820 9818 19876 9820
rect 19580 9766 19626 9818
rect 19626 9766 19636 9818
rect 19660 9766 19690 9818
rect 19690 9766 19702 9818
rect 19702 9766 19716 9818
rect 19740 9766 19754 9818
rect 19754 9766 19766 9818
rect 19766 9766 19796 9818
rect 19820 9766 19830 9818
rect 19830 9766 19876 9818
rect 19580 9764 19636 9766
rect 19660 9764 19716 9766
rect 19740 9764 19796 9766
rect 19820 9764 19876 9766
rect 19338 9560 19394 9616
rect 19580 8730 19636 8732
rect 19660 8730 19716 8732
rect 19740 8730 19796 8732
rect 19820 8730 19876 8732
rect 19580 8678 19626 8730
rect 19626 8678 19636 8730
rect 19660 8678 19690 8730
rect 19690 8678 19702 8730
rect 19702 8678 19716 8730
rect 19740 8678 19754 8730
rect 19754 8678 19766 8730
rect 19766 8678 19796 8730
rect 19820 8678 19830 8730
rect 19830 8678 19876 8730
rect 19580 8676 19636 8678
rect 19660 8676 19716 8678
rect 19740 8676 19796 8678
rect 19820 8676 19876 8678
rect 21914 10920 21970 10976
rect 20718 9288 20774 9344
rect 19580 7642 19636 7644
rect 19660 7642 19716 7644
rect 19740 7642 19796 7644
rect 19820 7642 19876 7644
rect 19580 7590 19626 7642
rect 19626 7590 19636 7642
rect 19660 7590 19690 7642
rect 19690 7590 19702 7642
rect 19702 7590 19716 7642
rect 19740 7590 19754 7642
rect 19754 7590 19766 7642
rect 19766 7590 19796 7642
rect 19820 7590 19830 7642
rect 19830 7590 19876 7642
rect 19580 7588 19636 7590
rect 19660 7588 19716 7590
rect 19740 7588 19796 7590
rect 19820 7588 19876 7590
rect 19580 6554 19636 6556
rect 19660 6554 19716 6556
rect 19740 6554 19796 6556
rect 19820 6554 19876 6556
rect 19580 6502 19626 6554
rect 19626 6502 19636 6554
rect 19660 6502 19690 6554
rect 19690 6502 19702 6554
rect 19702 6502 19716 6554
rect 19740 6502 19754 6554
rect 19754 6502 19766 6554
rect 19766 6502 19796 6554
rect 19820 6502 19830 6554
rect 19830 6502 19876 6554
rect 19580 6500 19636 6502
rect 19660 6500 19716 6502
rect 19740 6500 19796 6502
rect 19820 6500 19876 6502
rect 19580 5466 19636 5468
rect 19660 5466 19716 5468
rect 19740 5466 19796 5468
rect 19820 5466 19876 5468
rect 19580 5414 19626 5466
rect 19626 5414 19636 5466
rect 19660 5414 19690 5466
rect 19690 5414 19702 5466
rect 19702 5414 19716 5466
rect 19740 5414 19754 5466
rect 19754 5414 19766 5466
rect 19766 5414 19796 5466
rect 19820 5414 19830 5466
rect 19830 5414 19876 5466
rect 19580 5412 19636 5414
rect 19660 5412 19716 5414
rect 19740 5412 19796 5414
rect 19820 5412 19876 5414
rect 19580 4378 19636 4380
rect 19660 4378 19716 4380
rect 19740 4378 19796 4380
rect 19820 4378 19876 4380
rect 19580 4326 19626 4378
rect 19626 4326 19636 4378
rect 19660 4326 19690 4378
rect 19690 4326 19702 4378
rect 19702 4326 19716 4378
rect 19740 4326 19754 4378
rect 19754 4326 19766 4378
rect 19766 4326 19796 4378
rect 19820 4326 19830 4378
rect 19830 4326 19876 4378
rect 19580 4324 19636 4326
rect 19660 4324 19716 4326
rect 19740 4324 19796 4326
rect 19820 4324 19876 4326
rect 19580 3290 19636 3292
rect 19660 3290 19716 3292
rect 19740 3290 19796 3292
rect 19820 3290 19876 3292
rect 19580 3238 19626 3290
rect 19626 3238 19636 3290
rect 19660 3238 19690 3290
rect 19690 3238 19702 3290
rect 19702 3238 19716 3290
rect 19740 3238 19754 3290
rect 19754 3238 19766 3290
rect 19766 3238 19796 3290
rect 19820 3238 19830 3290
rect 19830 3238 19876 3290
rect 19580 3236 19636 3238
rect 19660 3236 19716 3238
rect 19740 3236 19796 3238
rect 19820 3236 19876 3238
rect 22466 13096 22522 13152
rect 23386 23024 23442 23080
rect 23110 22072 23166 22128
rect 28078 36796 28080 36816
rect 28080 36796 28132 36816
rect 28132 36796 28134 36816
rect 28078 36760 28134 36796
rect 34940 37562 34996 37564
rect 35020 37562 35076 37564
rect 35100 37562 35156 37564
rect 35180 37562 35236 37564
rect 34940 37510 34986 37562
rect 34986 37510 34996 37562
rect 35020 37510 35050 37562
rect 35050 37510 35062 37562
rect 35062 37510 35076 37562
rect 35100 37510 35114 37562
rect 35114 37510 35126 37562
rect 35126 37510 35156 37562
rect 35180 37510 35190 37562
rect 35190 37510 35236 37562
rect 34940 37508 34996 37510
rect 35020 37508 35076 37510
rect 35100 37508 35156 37510
rect 35180 37508 35236 37510
rect 23386 19216 23442 19272
rect 24858 23976 24914 24032
rect 24122 18300 24124 18320
rect 24124 18300 24176 18320
rect 24176 18300 24178 18320
rect 24122 18264 24178 18300
rect 23386 15272 23442 15328
rect 25042 18300 25044 18320
rect 25044 18300 25096 18320
rect 25096 18300 25098 18320
rect 25042 18264 25098 18300
rect 26514 20168 26570 20224
rect 26238 17040 26294 17096
rect 24766 15680 24822 15736
rect 23478 12552 23534 12608
rect 23018 12416 23074 12472
rect 23478 11736 23534 11792
rect 23018 11192 23074 11248
rect 22650 9580 22706 9616
rect 22650 9560 22652 9580
rect 22652 9560 22704 9580
rect 22704 9560 22706 9580
rect 24398 10920 24454 10976
rect 25226 12280 25282 12336
rect 24030 9832 24086 9888
rect 24030 9288 24086 9344
rect 26330 9560 26386 9616
rect 23938 3032 23994 3088
rect 24306 3052 24362 3088
rect 24306 3032 24308 3052
rect 24308 3032 24360 3052
rect 24360 3032 24362 3052
rect 19580 2202 19636 2204
rect 19660 2202 19716 2204
rect 19740 2202 19796 2204
rect 19820 2202 19876 2204
rect 19580 2150 19626 2202
rect 19626 2150 19636 2202
rect 19660 2150 19690 2202
rect 19690 2150 19702 2202
rect 19702 2150 19716 2202
rect 19740 2150 19754 2202
rect 19754 2150 19766 2202
rect 19766 2150 19796 2202
rect 19820 2150 19830 2202
rect 19830 2150 19876 2202
rect 19580 2148 19636 2150
rect 19660 2148 19716 2150
rect 19740 2148 19796 2150
rect 19820 2148 19876 2150
rect 27618 21528 27674 21584
rect 27342 20984 27398 21040
rect 26882 10512 26938 10568
rect 26882 3068 26884 3088
rect 26884 3068 26936 3088
rect 26936 3068 26938 3088
rect 26882 3032 26938 3068
rect 27802 9016 27858 9072
rect 28354 9288 28410 9344
rect 34940 36474 34996 36476
rect 35020 36474 35076 36476
rect 35100 36474 35156 36476
rect 35180 36474 35236 36476
rect 34940 36422 34986 36474
rect 34986 36422 34996 36474
rect 35020 36422 35050 36474
rect 35050 36422 35062 36474
rect 35062 36422 35076 36474
rect 35100 36422 35114 36474
rect 35114 36422 35126 36474
rect 35126 36422 35156 36474
rect 35180 36422 35190 36474
rect 35190 36422 35236 36474
rect 34940 36420 34996 36422
rect 35020 36420 35076 36422
rect 35100 36420 35156 36422
rect 35180 36420 35236 36422
rect 34940 35386 34996 35388
rect 35020 35386 35076 35388
rect 35100 35386 35156 35388
rect 35180 35386 35236 35388
rect 34940 35334 34986 35386
rect 34986 35334 34996 35386
rect 35020 35334 35050 35386
rect 35050 35334 35062 35386
rect 35062 35334 35076 35386
rect 35100 35334 35114 35386
rect 35114 35334 35126 35386
rect 35126 35334 35156 35386
rect 35180 35334 35190 35386
rect 35190 35334 35236 35386
rect 34940 35332 34996 35334
rect 35020 35332 35076 35334
rect 35100 35332 35156 35334
rect 35180 35332 35236 35334
rect 34940 34298 34996 34300
rect 35020 34298 35076 34300
rect 35100 34298 35156 34300
rect 35180 34298 35236 34300
rect 34940 34246 34986 34298
rect 34986 34246 34996 34298
rect 35020 34246 35050 34298
rect 35050 34246 35062 34298
rect 35062 34246 35076 34298
rect 35100 34246 35114 34298
rect 35114 34246 35126 34298
rect 35126 34246 35156 34298
rect 35180 34246 35190 34298
rect 35190 34246 35236 34298
rect 34940 34244 34996 34246
rect 35020 34244 35076 34246
rect 35100 34244 35156 34246
rect 35180 34244 35236 34246
rect 28906 9288 28962 9344
rect 30378 25472 30434 25528
rect 29642 23468 29644 23488
rect 29644 23468 29696 23488
rect 29696 23468 29698 23488
rect 29642 23432 29698 23468
rect 34940 33210 34996 33212
rect 35020 33210 35076 33212
rect 35100 33210 35156 33212
rect 35180 33210 35236 33212
rect 34940 33158 34986 33210
rect 34986 33158 34996 33210
rect 35020 33158 35050 33210
rect 35050 33158 35062 33210
rect 35062 33158 35076 33210
rect 35100 33158 35114 33210
rect 35114 33158 35126 33210
rect 35126 33158 35156 33210
rect 35180 33158 35190 33210
rect 35190 33158 35236 33210
rect 34940 33156 34996 33158
rect 35020 33156 35076 33158
rect 35100 33156 35156 33158
rect 35180 33156 35236 33158
rect 34940 32122 34996 32124
rect 35020 32122 35076 32124
rect 35100 32122 35156 32124
rect 35180 32122 35236 32124
rect 34940 32070 34986 32122
rect 34986 32070 34996 32122
rect 35020 32070 35050 32122
rect 35050 32070 35062 32122
rect 35062 32070 35076 32122
rect 35100 32070 35114 32122
rect 35114 32070 35126 32122
rect 35126 32070 35156 32122
rect 35180 32070 35190 32122
rect 35190 32070 35236 32122
rect 34940 32068 34996 32070
rect 35020 32068 35076 32070
rect 35100 32068 35156 32070
rect 35180 32068 35236 32070
rect 34940 31034 34996 31036
rect 35020 31034 35076 31036
rect 35100 31034 35156 31036
rect 35180 31034 35236 31036
rect 34940 30982 34986 31034
rect 34986 30982 34996 31034
rect 35020 30982 35050 31034
rect 35050 30982 35062 31034
rect 35062 30982 35076 31034
rect 35100 30982 35114 31034
rect 35114 30982 35126 31034
rect 35126 30982 35156 31034
rect 35180 30982 35190 31034
rect 35190 30982 35236 31034
rect 34940 30980 34996 30982
rect 35020 30980 35076 30982
rect 35100 30980 35156 30982
rect 35180 30980 35236 30982
rect 34940 29946 34996 29948
rect 35020 29946 35076 29948
rect 35100 29946 35156 29948
rect 35180 29946 35236 29948
rect 34940 29894 34986 29946
rect 34986 29894 34996 29946
rect 35020 29894 35050 29946
rect 35050 29894 35062 29946
rect 35062 29894 35076 29946
rect 35100 29894 35114 29946
rect 35114 29894 35126 29946
rect 35126 29894 35156 29946
rect 35180 29894 35190 29946
rect 35190 29894 35236 29946
rect 34940 29892 34996 29894
rect 35020 29892 35076 29894
rect 35100 29892 35156 29894
rect 35180 29892 35236 29894
rect 34940 28858 34996 28860
rect 35020 28858 35076 28860
rect 35100 28858 35156 28860
rect 35180 28858 35236 28860
rect 34940 28806 34986 28858
rect 34986 28806 34996 28858
rect 35020 28806 35050 28858
rect 35050 28806 35062 28858
rect 35062 28806 35076 28858
rect 35100 28806 35114 28858
rect 35114 28806 35126 28858
rect 35126 28806 35156 28858
rect 35180 28806 35190 28858
rect 35190 28806 35236 28858
rect 34940 28804 34996 28806
rect 35020 28804 35076 28806
rect 35100 28804 35156 28806
rect 35180 28804 35236 28806
rect 31298 25200 31354 25256
rect 33230 24248 33286 24304
rect 30562 21120 30618 21176
rect 33506 22652 33508 22672
rect 33508 22652 33560 22672
rect 33560 22652 33562 22672
rect 33506 22616 33562 22652
rect 34940 27770 34996 27772
rect 35020 27770 35076 27772
rect 35100 27770 35156 27772
rect 35180 27770 35236 27772
rect 34940 27718 34986 27770
rect 34986 27718 34996 27770
rect 35020 27718 35050 27770
rect 35050 27718 35062 27770
rect 35062 27718 35076 27770
rect 35100 27718 35114 27770
rect 35114 27718 35126 27770
rect 35126 27718 35156 27770
rect 35180 27718 35190 27770
rect 35190 27718 35236 27770
rect 34940 27716 34996 27718
rect 35020 27716 35076 27718
rect 35100 27716 35156 27718
rect 35180 27716 35236 27718
rect 37278 27920 37334 27976
rect 34940 26682 34996 26684
rect 35020 26682 35076 26684
rect 35100 26682 35156 26684
rect 35180 26682 35236 26684
rect 34940 26630 34986 26682
rect 34986 26630 34996 26682
rect 35020 26630 35050 26682
rect 35050 26630 35062 26682
rect 35062 26630 35076 26682
rect 35100 26630 35114 26682
rect 35114 26630 35126 26682
rect 35126 26630 35156 26682
rect 35180 26630 35190 26682
rect 35190 26630 35236 26682
rect 34940 26628 34996 26630
rect 35020 26628 35076 26630
rect 35100 26628 35156 26630
rect 35180 26628 35236 26630
rect 34940 25594 34996 25596
rect 35020 25594 35076 25596
rect 35100 25594 35156 25596
rect 35180 25594 35236 25596
rect 34940 25542 34986 25594
rect 34986 25542 34996 25594
rect 35020 25542 35050 25594
rect 35050 25542 35062 25594
rect 35062 25542 35076 25594
rect 35100 25542 35114 25594
rect 35114 25542 35126 25594
rect 35126 25542 35156 25594
rect 35180 25542 35190 25594
rect 35190 25542 35236 25594
rect 34940 25540 34996 25542
rect 35020 25540 35076 25542
rect 35100 25540 35156 25542
rect 35180 25540 35236 25542
rect 30378 20340 30380 20360
rect 30380 20340 30432 20360
rect 30432 20340 30434 20360
rect 30378 20304 30434 20340
rect 31022 15816 31078 15872
rect 30286 13096 30342 13152
rect 33322 21392 33378 21448
rect 31390 14320 31446 14376
rect 29826 9580 29882 9616
rect 29826 9560 29828 9580
rect 29828 9560 29880 9580
rect 29880 9560 29882 9580
rect 30746 9560 30802 9616
rect 31574 12416 31630 12472
rect 31022 9152 31078 9208
rect 33046 15544 33102 15600
rect 32954 14320 33010 14376
rect 34940 24506 34996 24508
rect 35020 24506 35076 24508
rect 35100 24506 35156 24508
rect 35180 24506 35236 24508
rect 34940 24454 34986 24506
rect 34986 24454 34996 24506
rect 35020 24454 35050 24506
rect 35050 24454 35062 24506
rect 35062 24454 35076 24506
rect 35100 24454 35114 24506
rect 35114 24454 35126 24506
rect 35126 24454 35156 24506
rect 35180 24454 35190 24506
rect 35190 24454 35236 24506
rect 34940 24452 34996 24454
rect 35020 24452 35076 24454
rect 35100 24452 35156 24454
rect 35180 24452 35236 24454
rect 34940 23418 34996 23420
rect 35020 23418 35076 23420
rect 35100 23418 35156 23420
rect 35180 23418 35236 23420
rect 34940 23366 34986 23418
rect 34986 23366 34996 23418
rect 35020 23366 35050 23418
rect 35050 23366 35062 23418
rect 35062 23366 35076 23418
rect 35100 23366 35114 23418
rect 35114 23366 35126 23418
rect 35126 23366 35156 23418
rect 35180 23366 35190 23418
rect 35190 23366 35236 23418
rect 34940 23364 34996 23366
rect 35020 23364 35076 23366
rect 35100 23364 35156 23366
rect 35180 23364 35236 23366
rect 34940 22330 34996 22332
rect 35020 22330 35076 22332
rect 35100 22330 35156 22332
rect 35180 22330 35236 22332
rect 34940 22278 34986 22330
rect 34986 22278 34996 22330
rect 35020 22278 35050 22330
rect 35050 22278 35062 22330
rect 35062 22278 35076 22330
rect 35100 22278 35114 22330
rect 35114 22278 35126 22330
rect 35126 22278 35156 22330
rect 35180 22278 35190 22330
rect 35190 22278 35236 22330
rect 34940 22276 34996 22278
rect 35020 22276 35076 22278
rect 35100 22276 35156 22278
rect 35180 22276 35236 22278
rect 36634 22500 36690 22536
rect 36634 22480 36636 22500
rect 36636 22480 36688 22500
rect 36688 22480 36690 22500
rect 42522 36760 42578 36816
rect 34940 21242 34996 21244
rect 35020 21242 35076 21244
rect 35100 21242 35156 21244
rect 35180 21242 35236 21244
rect 34940 21190 34986 21242
rect 34986 21190 34996 21242
rect 35020 21190 35050 21242
rect 35050 21190 35062 21242
rect 35062 21190 35076 21242
rect 35100 21190 35114 21242
rect 35114 21190 35126 21242
rect 35126 21190 35156 21242
rect 35180 21190 35190 21242
rect 35190 21190 35236 21242
rect 34940 21188 34996 21190
rect 35020 21188 35076 21190
rect 35100 21188 35156 21190
rect 35180 21188 35236 21190
rect 34610 20440 34666 20496
rect 34940 20154 34996 20156
rect 35020 20154 35076 20156
rect 35100 20154 35156 20156
rect 35180 20154 35236 20156
rect 34940 20102 34986 20154
rect 34986 20102 34996 20154
rect 35020 20102 35050 20154
rect 35050 20102 35062 20154
rect 35062 20102 35076 20154
rect 35100 20102 35114 20154
rect 35114 20102 35126 20154
rect 35126 20102 35156 20154
rect 35180 20102 35190 20154
rect 35190 20102 35236 20154
rect 34940 20100 34996 20102
rect 35020 20100 35076 20102
rect 35100 20100 35156 20102
rect 35180 20100 35236 20102
rect 38198 20848 38254 20904
rect 34940 19066 34996 19068
rect 35020 19066 35076 19068
rect 35100 19066 35156 19068
rect 35180 19066 35236 19068
rect 34940 19014 34986 19066
rect 34986 19014 34996 19066
rect 35020 19014 35050 19066
rect 35050 19014 35062 19066
rect 35062 19014 35076 19066
rect 35100 19014 35114 19066
rect 35114 19014 35126 19066
rect 35126 19014 35156 19066
rect 35180 19014 35190 19066
rect 35190 19014 35236 19066
rect 34940 19012 34996 19014
rect 35020 19012 35076 19014
rect 35100 19012 35156 19014
rect 35180 19012 35236 19014
rect 34940 17978 34996 17980
rect 35020 17978 35076 17980
rect 35100 17978 35156 17980
rect 35180 17978 35236 17980
rect 34940 17926 34986 17978
rect 34986 17926 34996 17978
rect 35020 17926 35050 17978
rect 35050 17926 35062 17978
rect 35062 17926 35076 17978
rect 35100 17926 35114 17978
rect 35114 17926 35126 17978
rect 35126 17926 35156 17978
rect 35180 17926 35190 17978
rect 35190 17926 35236 17978
rect 34940 17924 34996 17926
rect 35020 17924 35076 17926
rect 35100 17924 35156 17926
rect 35180 17924 35236 17926
rect 34940 16890 34996 16892
rect 35020 16890 35076 16892
rect 35100 16890 35156 16892
rect 35180 16890 35236 16892
rect 34940 16838 34986 16890
rect 34986 16838 34996 16890
rect 35020 16838 35050 16890
rect 35050 16838 35062 16890
rect 35062 16838 35076 16890
rect 35100 16838 35114 16890
rect 35114 16838 35126 16890
rect 35126 16838 35156 16890
rect 35180 16838 35190 16890
rect 35190 16838 35236 16890
rect 34940 16836 34996 16838
rect 35020 16836 35076 16838
rect 35100 16836 35156 16838
rect 35180 16836 35236 16838
rect 34940 15802 34996 15804
rect 35020 15802 35076 15804
rect 35100 15802 35156 15804
rect 35180 15802 35236 15804
rect 34940 15750 34986 15802
rect 34986 15750 34996 15802
rect 35020 15750 35050 15802
rect 35050 15750 35062 15802
rect 35062 15750 35076 15802
rect 35100 15750 35114 15802
rect 35114 15750 35126 15802
rect 35126 15750 35156 15802
rect 35180 15750 35190 15802
rect 35190 15750 35236 15802
rect 34940 15748 34996 15750
rect 35020 15748 35076 15750
rect 35100 15748 35156 15750
rect 35180 15748 35236 15750
rect 34940 14714 34996 14716
rect 35020 14714 35076 14716
rect 35100 14714 35156 14716
rect 35180 14714 35236 14716
rect 34940 14662 34986 14714
rect 34986 14662 34996 14714
rect 35020 14662 35050 14714
rect 35050 14662 35062 14714
rect 35062 14662 35076 14714
rect 35100 14662 35114 14714
rect 35114 14662 35126 14714
rect 35126 14662 35156 14714
rect 35180 14662 35190 14714
rect 35190 14662 35236 14714
rect 34940 14660 34996 14662
rect 35020 14660 35076 14662
rect 35100 14660 35156 14662
rect 35180 14660 35236 14662
rect 34940 13626 34996 13628
rect 35020 13626 35076 13628
rect 35100 13626 35156 13628
rect 35180 13626 35236 13628
rect 34940 13574 34986 13626
rect 34986 13574 34996 13626
rect 35020 13574 35050 13626
rect 35050 13574 35062 13626
rect 35062 13574 35076 13626
rect 35100 13574 35114 13626
rect 35114 13574 35126 13626
rect 35126 13574 35156 13626
rect 35180 13574 35190 13626
rect 35190 13574 35236 13626
rect 34940 13572 34996 13574
rect 35020 13572 35076 13574
rect 35100 13572 35156 13574
rect 35180 13572 35236 13574
rect 34940 12538 34996 12540
rect 35020 12538 35076 12540
rect 35100 12538 35156 12540
rect 35180 12538 35236 12540
rect 34940 12486 34986 12538
rect 34986 12486 34996 12538
rect 35020 12486 35050 12538
rect 35050 12486 35062 12538
rect 35062 12486 35076 12538
rect 35100 12486 35114 12538
rect 35114 12486 35126 12538
rect 35126 12486 35156 12538
rect 35180 12486 35190 12538
rect 35190 12486 35236 12538
rect 34940 12484 34996 12486
rect 35020 12484 35076 12486
rect 35100 12484 35156 12486
rect 35180 12484 35236 12486
rect 34940 11450 34996 11452
rect 35020 11450 35076 11452
rect 35100 11450 35156 11452
rect 35180 11450 35236 11452
rect 34940 11398 34986 11450
rect 34986 11398 34996 11450
rect 35020 11398 35050 11450
rect 35050 11398 35062 11450
rect 35062 11398 35076 11450
rect 35100 11398 35114 11450
rect 35114 11398 35126 11450
rect 35126 11398 35156 11450
rect 35180 11398 35190 11450
rect 35190 11398 35236 11450
rect 34940 11396 34996 11398
rect 35020 11396 35076 11398
rect 35100 11396 35156 11398
rect 35180 11396 35236 11398
rect 34940 10362 34996 10364
rect 35020 10362 35076 10364
rect 35100 10362 35156 10364
rect 35180 10362 35236 10364
rect 34940 10310 34986 10362
rect 34986 10310 34996 10362
rect 35020 10310 35050 10362
rect 35050 10310 35062 10362
rect 35062 10310 35076 10362
rect 35100 10310 35114 10362
rect 35114 10310 35126 10362
rect 35126 10310 35156 10362
rect 35180 10310 35190 10362
rect 35190 10310 35236 10362
rect 34940 10308 34996 10310
rect 35020 10308 35076 10310
rect 35100 10308 35156 10310
rect 35180 10308 35236 10310
rect 35346 9868 35348 9888
rect 35348 9868 35400 9888
rect 35400 9868 35402 9888
rect 35346 9832 35402 9868
rect 34940 9274 34996 9276
rect 35020 9274 35076 9276
rect 35100 9274 35156 9276
rect 35180 9274 35236 9276
rect 34940 9222 34986 9274
rect 34986 9222 34996 9274
rect 35020 9222 35050 9274
rect 35050 9222 35062 9274
rect 35062 9222 35076 9274
rect 35100 9222 35114 9274
rect 35114 9222 35126 9274
rect 35126 9222 35156 9274
rect 35180 9222 35190 9274
rect 35190 9222 35236 9274
rect 34940 9220 34996 9222
rect 35020 9220 35076 9222
rect 35100 9220 35156 9222
rect 35180 9220 35236 9222
rect 34940 8186 34996 8188
rect 35020 8186 35076 8188
rect 35100 8186 35156 8188
rect 35180 8186 35236 8188
rect 34940 8134 34986 8186
rect 34986 8134 34996 8186
rect 35020 8134 35050 8186
rect 35050 8134 35062 8186
rect 35062 8134 35076 8186
rect 35100 8134 35114 8186
rect 35114 8134 35126 8186
rect 35126 8134 35156 8186
rect 35180 8134 35190 8186
rect 35190 8134 35236 8186
rect 34940 8132 34996 8134
rect 35020 8132 35076 8134
rect 35100 8132 35156 8134
rect 35180 8132 35236 8134
rect 34940 7098 34996 7100
rect 35020 7098 35076 7100
rect 35100 7098 35156 7100
rect 35180 7098 35236 7100
rect 34940 7046 34986 7098
rect 34986 7046 34996 7098
rect 35020 7046 35050 7098
rect 35050 7046 35062 7098
rect 35062 7046 35076 7098
rect 35100 7046 35114 7098
rect 35114 7046 35126 7098
rect 35126 7046 35156 7098
rect 35180 7046 35190 7098
rect 35190 7046 35236 7098
rect 34940 7044 34996 7046
rect 35020 7044 35076 7046
rect 35100 7044 35156 7046
rect 35180 7044 35236 7046
rect 38014 19252 38016 19272
rect 38016 19252 38068 19272
rect 38068 19252 38070 19272
rect 38014 19216 38070 19252
rect 38750 17040 38806 17096
rect 37554 12688 37610 12744
rect 37370 11192 37426 11248
rect 40222 17484 40224 17504
rect 40224 17484 40276 17504
rect 40276 17484 40278 17504
rect 40222 17448 40278 17484
rect 40038 16632 40094 16688
rect 39854 15952 39910 16008
rect 42706 36780 42762 36816
rect 42706 36760 42708 36780
rect 42708 36760 42760 36780
rect 42760 36760 42762 36780
rect 41786 18672 41842 18728
rect 40038 15136 40094 15192
rect 40314 12144 40370 12200
rect 35898 9424 35954 9480
rect 34940 6010 34996 6012
rect 35020 6010 35076 6012
rect 35100 6010 35156 6012
rect 35180 6010 35236 6012
rect 34940 5958 34986 6010
rect 34986 5958 34996 6010
rect 35020 5958 35050 6010
rect 35050 5958 35062 6010
rect 35062 5958 35076 6010
rect 35100 5958 35114 6010
rect 35114 5958 35126 6010
rect 35126 5958 35156 6010
rect 35180 5958 35190 6010
rect 35190 5958 35236 6010
rect 34940 5956 34996 5958
rect 35020 5956 35076 5958
rect 35100 5956 35156 5958
rect 35180 5956 35236 5958
rect 34940 4922 34996 4924
rect 35020 4922 35076 4924
rect 35100 4922 35156 4924
rect 35180 4922 35236 4924
rect 34940 4870 34986 4922
rect 34986 4870 34996 4922
rect 35020 4870 35050 4922
rect 35050 4870 35062 4922
rect 35062 4870 35076 4922
rect 35100 4870 35114 4922
rect 35114 4870 35126 4922
rect 35126 4870 35156 4922
rect 35180 4870 35190 4922
rect 35190 4870 35236 4922
rect 34940 4868 34996 4870
rect 35020 4868 35076 4870
rect 35100 4868 35156 4870
rect 35180 4868 35236 4870
rect 34940 3834 34996 3836
rect 35020 3834 35076 3836
rect 35100 3834 35156 3836
rect 35180 3834 35236 3836
rect 34940 3782 34986 3834
rect 34986 3782 34996 3834
rect 35020 3782 35050 3834
rect 35050 3782 35062 3834
rect 35062 3782 35076 3834
rect 35100 3782 35114 3834
rect 35114 3782 35126 3834
rect 35126 3782 35156 3834
rect 35180 3782 35190 3834
rect 35190 3782 35236 3834
rect 34940 3780 34996 3782
rect 35020 3780 35076 3782
rect 35100 3780 35156 3782
rect 35180 3780 35236 3782
rect 39118 8880 39174 8936
rect 39670 7284 39672 7304
rect 39672 7284 39724 7304
rect 39724 7284 39726 7304
rect 39670 7248 39726 7284
rect 41970 15444 41972 15464
rect 41972 15444 42024 15464
rect 42024 15444 42026 15464
rect 41970 15408 42026 15444
rect 43350 19352 43406 19408
rect 44362 14320 44418 14376
rect 34940 2746 34996 2748
rect 35020 2746 35076 2748
rect 35100 2746 35156 2748
rect 35180 2746 35236 2748
rect 34940 2694 34986 2746
rect 34986 2694 34996 2746
rect 35020 2694 35050 2746
rect 35050 2694 35062 2746
rect 35062 2694 35076 2746
rect 35100 2694 35114 2746
rect 35114 2694 35126 2746
rect 35126 2694 35156 2746
rect 35180 2694 35190 2746
rect 35190 2694 35236 2746
rect 34940 2692 34996 2694
rect 35020 2692 35076 2694
rect 35100 2692 35156 2694
rect 35180 2692 35236 2694
rect 46662 13232 46718 13288
rect 47766 10104 47822 10160
rect 50300 37018 50356 37020
rect 50380 37018 50436 37020
rect 50460 37018 50516 37020
rect 50540 37018 50596 37020
rect 50300 36966 50346 37018
rect 50346 36966 50356 37018
rect 50380 36966 50410 37018
rect 50410 36966 50422 37018
rect 50422 36966 50436 37018
rect 50460 36966 50474 37018
rect 50474 36966 50486 37018
rect 50486 36966 50516 37018
rect 50540 36966 50550 37018
rect 50550 36966 50596 37018
rect 50300 36964 50356 36966
rect 50380 36964 50436 36966
rect 50460 36964 50516 36966
rect 50540 36964 50596 36966
rect 50300 35930 50356 35932
rect 50380 35930 50436 35932
rect 50460 35930 50516 35932
rect 50540 35930 50596 35932
rect 50300 35878 50346 35930
rect 50346 35878 50356 35930
rect 50380 35878 50410 35930
rect 50410 35878 50422 35930
rect 50422 35878 50436 35930
rect 50460 35878 50474 35930
rect 50474 35878 50486 35930
rect 50486 35878 50516 35930
rect 50540 35878 50550 35930
rect 50550 35878 50596 35930
rect 50300 35876 50356 35878
rect 50380 35876 50436 35878
rect 50460 35876 50516 35878
rect 50540 35876 50596 35878
rect 50300 34842 50356 34844
rect 50380 34842 50436 34844
rect 50460 34842 50516 34844
rect 50540 34842 50596 34844
rect 50300 34790 50346 34842
rect 50346 34790 50356 34842
rect 50380 34790 50410 34842
rect 50410 34790 50422 34842
rect 50422 34790 50436 34842
rect 50460 34790 50474 34842
rect 50474 34790 50486 34842
rect 50486 34790 50516 34842
rect 50540 34790 50550 34842
rect 50550 34790 50596 34842
rect 50300 34788 50356 34790
rect 50380 34788 50436 34790
rect 50460 34788 50516 34790
rect 50540 34788 50596 34790
rect 50300 33754 50356 33756
rect 50380 33754 50436 33756
rect 50460 33754 50516 33756
rect 50540 33754 50596 33756
rect 50300 33702 50346 33754
rect 50346 33702 50356 33754
rect 50380 33702 50410 33754
rect 50410 33702 50422 33754
rect 50422 33702 50436 33754
rect 50460 33702 50474 33754
rect 50474 33702 50486 33754
rect 50486 33702 50516 33754
rect 50540 33702 50550 33754
rect 50550 33702 50596 33754
rect 50300 33700 50356 33702
rect 50380 33700 50436 33702
rect 50460 33700 50516 33702
rect 50540 33700 50596 33702
rect 50300 32666 50356 32668
rect 50380 32666 50436 32668
rect 50460 32666 50516 32668
rect 50540 32666 50596 32668
rect 50300 32614 50346 32666
rect 50346 32614 50356 32666
rect 50380 32614 50410 32666
rect 50410 32614 50422 32666
rect 50422 32614 50436 32666
rect 50460 32614 50474 32666
rect 50474 32614 50486 32666
rect 50486 32614 50516 32666
rect 50540 32614 50550 32666
rect 50550 32614 50596 32666
rect 50300 32612 50356 32614
rect 50380 32612 50436 32614
rect 50460 32612 50516 32614
rect 50540 32612 50596 32614
rect 50300 31578 50356 31580
rect 50380 31578 50436 31580
rect 50460 31578 50516 31580
rect 50540 31578 50596 31580
rect 50300 31526 50346 31578
rect 50346 31526 50356 31578
rect 50380 31526 50410 31578
rect 50410 31526 50422 31578
rect 50422 31526 50436 31578
rect 50460 31526 50474 31578
rect 50474 31526 50486 31578
rect 50486 31526 50516 31578
rect 50540 31526 50550 31578
rect 50550 31526 50596 31578
rect 50300 31524 50356 31526
rect 50380 31524 50436 31526
rect 50460 31524 50516 31526
rect 50540 31524 50596 31526
rect 50300 30490 50356 30492
rect 50380 30490 50436 30492
rect 50460 30490 50516 30492
rect 50540 30490 50596 30492
rect 50300 30438 50346 30490
rect 50346 30438 50356 30490
rect 50380 30438 50410 30490
rect 50410 30438 50422 30490
rect 50422 30438 50436 30490
rect 50460 30438 50474 30490
rect 50474 30438 50486 30490
rect 50486 30438 50516 30490
rect 50540 30438 50550 30490
rect 50550 30438 50596 30490
rect 50300 30436 50356 30438
rect 50380 30436 50436 30438
rect 50460 30436 50516 30438
rect 50540 30436 50596 30438
rect 50300 29402 50356 29404
rect 50380 29402 50436 29404
rect 50460 29402 50516 29404
rect 50540 29402 50596 29404
rect 50300 29350 50346 29402
rect 50346 29350 50356 29402
rect 50380 29350 50410 29402
rect 50410 29350 50422 29402
rect 50422 29350 50436 29402
rect 50460 29350 50474 29402
rect 50474 29350 50486 29402
rect 50486 29350 50516 29402
rect 50540 29350 50550 29402
rect 50550 29350 50596 29402
rect 50300 29348 50356 29350
rect 50380 29348 50436 29350
rect 50460 29348 50516 29350
rect 50540 29348 50596 29350
rect 50300 28314 50356 28316
rect 50380 28314 50436 28316
rect 50460 28314 50516 28316
rect 50540 28314 50596 28316
rect 50300 28262 50346 28314
rect 50346 28262 50356 28314
rect 50380 28262 50410 28314
rect 50410 28262 50422 28314
rect 50422 28262 50436 28314
rect 50460 28262 50474 28314
rect 50474 28262 50486 28314
rect 50486 28262 50516 28314
rect 50540 28262 50550 28314
rect 50550 28262 50596 28314
rect 50300 28260 50356 28262
rect 50380 28260 50436 28262
rect 50460 28260 50516 28262
rect 50540 28260 50596 28262
rect 50300 27226 50356 27228
rect 50380 27226 50436 27228
rect 50460 27226 50516 27228
rect 50540 27226 50596 27228
rect 50300 27174 50346 27226
rect 50346 27174 50356 27226
rect 50380 27174 50410 27226
rect 50410 27174 50422 27226
rect 50422 27174 50436 27226
rect 50460 27174 50474 27226
rect 50474 27174 50486 27226
rect 50486 27174 50516 27226
rect 50540 27174 50550 27226
rect 50550 27174 50596 27226
rect 50300 27172 50356 27174
rect 50380 27172 50436 27174
rect 50460 27172 50516 27174
rect 50540 27172 50596 27174
rect 50300 26138 50356 26140
rect 50380 26138 50436 26140
rect 50460 26138 50516 26140
rect 50540 26138 50596 26140
rect 50300 26086 50346 26138
rect 50346 26086 50356 26138
rect 50380 26086 50410 26138
rect 50410 26086 50422 26138
rect 50422 26086 50436 26138
rect 50460 26086 50474 26138
rect 50474 26086 50486 26138
rect 50486 26086 50516 26138
rect 50540 26086 50550 26138
rect 50550 26086 50596 26138
rect 50300 26084 50356 26086
rect 50380 26084 50436 26086
rect 50460 26084 50516 26086
rect 50540 26084 50596 26086
rect 50300 25050 50356 25052
rect 50380 25050 50436 25052
rect 50460 25050 50516 25052
rect 50540 25050 50596 25052
rect 50300 24998 50346 25050
rect 50346 24998 50356 25050
rect 50380 24998 50410 25050
rect 50410 24998 50422 25050
rect 50422 24998 50436 25050
rect 50460 24998 50474 25050
rect 50474 24998 50486 25050
rect 50486 24998 50516 25050
rect 50540 24998 50550 25050
rect 50550 24998 50596 25050
rect 50300 24996 50356 24998
rect 50380 24996 50436 24998
rect 50460 24996 50516 24998
rect 50540 24996 50596 24998
rect 50300 23962 50356 23964
rect 50380 23962 50436 23964
rect 50460 23962 50516 23964
rect 50540 23962 50596 23964
rect 50300 23910 50346 23962
rect 50346 23910 50356 23962
rect 50380 23910 50410 23962
rect 50410 23910 50422 23962
rect 50422 23910 50436 23962
rect 50460 23910 50474 23962
rect 50474 23910 50486 23962
rect 50486 23910 50516 23962
rect 50540 23910 50550 23962
rect 50550 23910 50596 23962
rect 50300 23908 50356 23910
rect 50380 23908 50436 23910
rect 50460 23908 50516 23910
rect 50540 23908 50596 23910
rect 50300 22874 50356 22876
rect 50380 22874 50436 22876
rect 50460 22874 50516 22876
rect 50540 22874 50596 22876
rect 50300 22822 50346 22874
rect 50346 22822 50356 22874
rect 50380 22822 50410 22874
rect 50410 22822 50422 22874
rect 50422 22822 50436 22874
rect 50460 22822 50474 22874
rect 50474 22822 50486 22874
rect 50486 22822 50516 22874
rect 50540 22822 50550 22874
rect 50550 22822 50596 22874
rect 50300 22820 50356 22822
rect 50380 22820 50436 22822
rect 50460 22820 50516 22822
rect 50540 22820 50596 22822
rect 50300 21786 50356 21788
rect 50380 21786 50436 21788
rect 50460 21786 50516 21788
rect 50540 21786 50596 21788
rect 50300 21734 50346 21786
rect 50346 21734 50356 21786
rect 50380 21734 50410 21786
rect 50410 21734 50422 21786
rect 50422 21734 50436 21786
rect 50460 21734 50474 21786
rect 50474 21734 50486 21786
rect 50486 21734 50516 21786
rect 50540 21734 50550 21786
rect 50550 21734 50596 21786
rect 50300 21732 50356 21734
rect 50380 21732 50436 21734
rect 50460 21732 50516 21734
rect 50540 21732 50596 21734
rect 50300 20698 50356 20700
rect 50380 20698 50436 20700
rect 50460 20698 50516 20700
rect 50540 20698 50596 20700
rect 50300 20646 50346 20698
rect 50346 20646 50356 20698
rect 50380 20646 50410 20698
rect 50410 20646 50422 20698
rect 50422 20646 50436 20698
rect 50460 20646 50474 20698
rect 50474 20646 50486 20698
rect 50486 20646 50516 20698
rect 50540 20646 50550 20698
rect 50550 20646 50596 20698
rect 50300 20644 50356 20646
rect 50380 20644 50436 20646
rect 50460 20644 50516 20646
rect 50540 20644 50596 20646
rect 50300 19610 50356 19612
rect 50380 19610 50436 19612
rect 50460 19610 50516 19612
rect 50540 19610 50596 19612
rect 50300 19558 50346 19610
rect 50346 19558 50356 19610
rect 50380 19558 50410 19610
rect 50410 19558 50422 19610
rect 50422 19558 50436 19610
rect 50460 19558 50474 19610
rect 50474 19558 50486 19610
rect 50486 19558 50516 19610
rect 50540 19558 50550 19610
rect 50550 19558 50596 19610
rect 50300 19556 50356 19558
rect 50380 19556 50436 19558
rect 50460 19556 50516 19558
rect 50540 19556 50596 19558
rect 50300 18522 50356 18524
rect 50380 18522 50436 18524
rect 50460 18522 50516 18524
rect 50540 18522 50596 18524
rect 50300 18470 50346 18522
rect 50346 18470 50356 18522
rect 50380 18470 50410 18522
rect 50410 18470 50422 18522
rect 50422 18470 50436 18522
rect 50460 18470 50474 18522
rect 50474 18470 50486 18522
rect 50486 18470 50516 18522
rect 50540 18470 50550 18522
rect 50550 18470 50596 18522
rect 50300 18468 50356 18470
rect 50380 18468 50436 18470
rect 50460 18468 50516 18470
rect 50540 18468 50596 18470
rect 50158 17584 50214 17640
rect 50300 17434 50356 17436
rect 50380 17434 50436 17436
rect 50460 17434 50516 17436
rect 50540 17434 50596 17436
rect 50300 17382 50346 17434
rect 50346 17382 50356 17434
rect 50380 17382 50410 17434
rect 50410 17382 50422 17434
rect 50422 17382 50436 17434
rect 50460 17382 50474 17434
rect 50474 17382 50486 17434
rect 50486 17382 50516 17434
rect 50540 17382 50550 17434
rect 50550 17382 50596 17434
rect 50300 17380 50356 17382
rect 50380 17380 50436 17382
rect 50460 17380 50516 17382
rect 50540 17380 50596 17382
rect 52458 25880 52514 25936
rect 57886 37440 57942 37496
rect 54942 31356 54944 31376
rect 54944 31356 54996 31376
rect 54996 31356 54998 31376
rect 54942 31320 54998 31356
rect 50300 16346 50356 16348
rect 50380 16346 50436 16348
rect 50460 16346 50516 16348
rect 50540 16346 50596 16348
rect 50300 16294 50346 16346
rect 50346 16294 50356 16346
rect 50380 16294 50410 16346
rect 50410 16294 50422 16346
rect 50422 16294 50436 16346
rect 50460 16294 50474 16346
rect 50474 16294 50486 16346
rect 50486 16294 50516 16346
rect 50540 16294 50550 16346
rect 50550 16294 50596 16346
rect 50300 16292 50356 16294
rect 50380 16292 50436 16294
rect 50460 16292 50516 16294
rect 50540 16292 50596 16294
rect 49790 14864 49846 14920
rect 50300 15258 50356 15260
rect 50380 15258 50436 15260
rect 50460 15258 50516 15260
rect 50540 15258 50596 15260
rect 50300 15206 50346 15258
rect 50346 15206 50356 15258
rect 50380 15206 50410 15258
rect 50410 15206 50422 15258
rect 50422 15206 50436 15258
rect 50460 15206 50474 15258
rect 50474 15206 50486 15258
rect 50486 15206 50516 15258
rect 50540 15206 50550 15258
rect 50550 15206 50596 15258
rect 50300 15204 50356 15206
rect 50380 15204 50436 15206
rect 50460 15204 50516 15206
rect 50540 15204 50596 15206
rect 50300 14170 50356 14172
rect 50380 14170 50436 14172
rect 50460 14170 50516 14172
rect 50540 14170 50596 14172
rect 50300 14118 50346 14170
rect 50346 14118 50356 14170
rect 50380 14118 50410 14170
rect 50410 14118 50422 14170
rect 50422 14118 50436 14170
rect 50460 14118 50474 14170
rect 50474 14118 50486 14170
rect 50486 14118 50516 14170
rect 50540 14118 50550 14170
rect 50550 14118 50596 14170
rect 50300 14116 50356 14118
rect 50380 14116 50436 14118
rect 50460 14116 50516 14118
rect 50540 14116 50596 14118
rect 50300 13082 50356 13084
rect 50380 13082 50436 13084
rect 50460 13082 50516 13084
rect 50540 13082 50596 13084
rect 50300 13030 50346 13082
rect 50346 13030 50356 13082
rect 50380 13030 50410 13082
rect 50410 13030 50422 13082
rect 50422 13030 50436 13082
rect 50460 13030 50474 13082
rect 50474 13030 50486 13082
rect 50486 13030 50516 13082
rect 50540 13030 50550 13082
rect 50550 13030 50596 13082
rect 50300 13028 50356 13030
rect 50380 13028 50436 13030
rect 50460 13028 50516 13030
rect 50540 13028 50596 13030
rect 50300 11994 50356 11996
rect 50380 11994 50436 11996
rect 50460 11994 50516 11996
rect 50540 11994 50596 11996
rect 50300 11942 50346 11994
rect 50346 11942 50356 11994
rect 50380 11942 50410 11994
rect 50410 11942 50422 11994
rect 50422 11942 50436 11994
rect 50460 11942 50474 11994
rect 50474 11942 50486 11994
rect 50486 11942 50516 11994
rect 50540 11942 50550 11994
rect 50550 11942 50596 11994
rect 50300 11940 50356 11942
rect 50380 11940 50436 11942
rect 50460 11940 50516 11942
rect 50540 11940 50596 11942
rect 50300 10906 50356 10908
rect 50380 10906 50436 10908
rect 50460 10906 50516 10908
rect 50540 10906 50596 10908
rect 50300 10854 50346 10906
rect 50346 10854 50356 10906
rect 50380 10854 50410 10906
rect 50410 10854 50422 10906
rect 50422 10854 50436 10906
rect 50460 10854 50474 10906
rect 50474 10854 50486 10906
rect 50486 10854 50516 10906
rect 50540 10854 50550 10906
rect 50550 10854 50596 10906
rect 50300 10852 50356 10854
rect 50380 10852 50436 10854
rect 50460 10852 50516 10854
rect 50540 10852 50596 10854
rect 51170 9988 51226 10024
rect 51170 9968 51172 9988
rect 51172 9968 51224 9988
rect 51224 9968 51226 9988
rect 50300 9818 50356 9820
rect 50380 9818 50436 9820
rect 50460 9818 50516 9820
rect 50540 9818 50596 9820
rect 50300 9766 50346 9818
rect 50346 9766 50356 9818
rect 50380 9766 50410 9818
rect 50410 9766 50422 9818
rect 50422 9766 50436 9818
rect 50460 9766 50474 9818
rect 50474 9766 50486 9818
rect 50486 9766 50516 9818
rect 50540 9766 50550 9818
rect 50550 9766 50596 9818
rect 50300 9764 50356 9766
rect 50380 9764 50436 9766
rect 50460 9764 50516 9766
rect 50540 9764 50596 9766
rect 50300 8730 50356 8732
rect 50380 8730 50436 8732
rect 50460 8730 50516 8732
rect 50540 8730 50596 8732
rect 50300 8678 50346 8730
rect 50346 8678 50356 8730
rect 50380 8678 50410 8730
rect 50410 8678 50422 8730
rect 50422 8678 50436 8730
rect 50460 8678 50474 8730
rect 50474 8678 50486 8730
rect 50486 8678 50516 8730
rect 50540 8678 50550 8730
rect 50550 8678 50596 8730
rect 50300 8676 50356 8678
rect 50380 8676 50436 8678
rect 50460 8676 50516 8678
rect 50540 8676 50596 8678
rect 50300 7642 50356 7644
rect 50380 7642 50436 7644
rect 50460 7642 50516 7644
rect 50540 7642 50596 7644
rect 50300 7590 50346 7642
rect 50346 7590 50356 7642
rect 50380 7590 50410 7642
rect 50410 7590 50422 7642
rect 50422 7590 50436 7642
rect 50460 7590 50474 7642
rect 50474 7590 50486 7642
rect 50486 7590 50516 7642
rect 50540 7590 50550 7642
rect 50550 7590 50596 7642
rect 50300 7588 50356 7590
rect 50380 7588 50436 7590
rect 50460 7588 50516 7590
rect 50540 7588 50596 7590
rect 50300 6554 50356 6556
rect 50380 6554 50436 6556
rect 50460 6554 50516 6556
rect 50540 6554 50596 6556
rect 50300 6502 50346 6554
rect 50346 6502 50356 6554
rect 50380 6502 50410 6554
rect 50410 6502 50422 6554
rect 50422 6502 50436 6554
rect 50460 6502 50474 6554
rect 50474 6502 50486 6554
rect 50486 6502 50516 6554
rect 50540 6502 50550 6554
rect 50550 6502 50596 6554
rect 50300 6500 50356 6502
rect 50380 6500 50436 6502
rect 50460 6500 50516 6502
rect 50540 6500 50596 6502
rect 50300 5466 50356 5468
rect 50380 5466 50436 5468
rect 50460 5466 50516 5468
rect 50540 5466 50596 5468
rect 50300 5414 50346 5466
rect 50346 5414 50356 5466
rect 50380 5414 50410 5466
rect 50410 5414 50422 5466
rect 50422 5414 50436 5466
rect 50460 5414 50474 5466
rect 50474 5414 50486 5466
rect 50486 5414 50516 5466
rect 50540 5414 50550 5466
rect 50550 5414 50596 5466
rect 50300 5412 50356 5414
rect 50380 5412 50436 5414
rect 50460 5412 50516 5414
rect 50540 5412 50596 5414
rect 50300 4378 50356 4380
rect 50380 4378 50436 4380
rect 50460 4378 50516 4380
rect 50540 4378 50596 4380
rect 50300 4326 50346 4378
rect 50346 4326 50356 4378
rect 50380 4326 50410 4378
rect 50410 4326 50422 4378
rect 50422 4326 50436 4378
rect 50460 4326 50474 4378
rect 50474 4326 50486 4378
rect 50486 4326 50516 4378
rect 50540 4326 50550 4378
rect 50550 4326 50596 4378
rect 50300 4324 50356 4326
rect 50380 4324 50436 4326
rect 50460 4324 50516 4326
rect 50540 4324 50596 4326
rect 50300 3290 50356 3292
rect 50380 3290 50436 3292
rect 50460 3290 50516 3292
rect 50540 3290 50596 3292
rect 50300 3238 50346 3290
rect 50346 3238 50356 3290
rect 50380 3238 50410 3290
rect 50410 3238 50422 3290
rect 50422 3238 50436 3290
rect 50460 3238 50474 3290
rect 50474 3238 50486 3290
rect 50486 3238 50516 3290
rect 50540 3238 50550 3290
rect 50550 3238 50596 3290
rect 50300 3236 50356 3238
rect 50380 3236 50436 3238
rect 50460 3236 50516 3238
rect 50540 3236 50596 3238
rect 51722 10668 51778 10704
rect 51722 10648 51724 10668
rect 51724 10648 51776 10668
rect 51776 10648 51778 10668
rect 53562 15564 53618 15600
rect 53562 15544 53564 15564
rect 53564 15544 53616 15564
rect 53616 15544 53618 15564
rect 52734 11600 52790 11656
rect 56782 24132 56838 24168
rect 56782 24112 56784 24132
rect 56784 24112 56836 24132
rect 56836 24112 56838 24132
rect 50300 2202 50356 2204
rect 50380 2202 50436 2204
rect 50460 2202 50516 2204
rect 50540 2202 50596 2204
rect 50300 2150 50346 2202
rect 50346 2150 50356 2202
rect 50380 2150 50410 2202
rect 50410 2150 50422 2202
rect 50422 2150 50436 2202
rect 50460 2150 50474 2202
rect 50474 2150 50486 2202
rect 50486 2150 50516 2202
rect 50540 2150 50550 2202
rect 50550 2150 50596 2202
rect 50300 2148 50356 2150
rect 50380 2148 50436 2150
rect 50460 2148 50516 2150
rect 50540 2148 50596 2150
rect 56046 11756 56102 11792
rect 56046 11736 56048 11756
rect 56048 11736 56100 11756
rect 56100 11736 56102 11756
rect 57886 35672 57942 35728
rect 58162 35400 58218 35456
rect 58162 33360 58218 33416
rect 57886 31320 57942 31376
rect 58162 29280 58218 29336
rect 58162 27240 58218 27296
rect 58070 25200 58126 25256
rect 57886 23160 57942 23216
rect 57518 7812 57574 7848
rect 57518 7792 57520 7812
rect 57520 7792 57572 7812
rect 57572 7792 57574 7812
rect 56782 6740 56784 6760
rect 56784 6740 56836 6760
rect 56836 6740 56838 6760
rect 56782 6704 56838 6740
rect 58162 20476 58164 20496
rect 58164 20476 58216 20496
rect 58216 20476 58218 20496
rect 58162 20440 58218 20476
rect 58070 18400 58126 18456
rect 58162 16360 58218 16416
rect 58070 14320 58126 14376
rect 58162 12280 58218 12336
rect 58070 10240 58126 10296
rect 58070 8200 58126 8256
rect 58070 6180 58126 6216
rect 58070 6160 58072 6180
rect 58072 6160 58124 6180
rect 58124 6160 58126 6180
rect 58070 3476 58072 3496
rect 58072 3476 58124 3496
rect 58124 3476 58126 3496
rect 58070 3440 58126 3476
rect 57242 1400 57298 1456
<< metal3 >>
rect 0 38178 800 38208
rect 1485 38178 1551 38181
rect 0 38176 1551 38178
rect 0 38120 1490 38176
rect 1546 38120 1551 38176
rect 0 38118 1551 38120
rect 0 38088 800 38118
rect 1485 38115 1551 38118
rect 4208 37568 4528 37569
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 37503 4528 37504
rect 34928 37568 35248 37569
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 37503 35248 37504
rect 57881 37498 57947 37501
rect 59200 37498 60000 37528
rect 57881 37496 60000 37498
rect 57881 37440 57886 37496
rect 57942 37440 60000 37496
rect 57881 37438 60000 37440
rect 57881 37435 57947 37438
rect 59200 37408 60000 37438
rect 19568 37024 19888 37025
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 36959 19888 36960
rect 50288 37024 50608 37025
rect 50288 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50608 37024
rect 50288 36959 50608 36960
rect 28073 36818 28139 36821
rect 42517 36818 42583 36821
rect 42701 36818 42767 36821
rect 28073 36816 42767 36818
rect 28073 36760 28078 36816
rect 28134 36760 42522 36816
rect 42578 36760 42706 36816
rect 42762 36760 42767 36816
rect 28073 36758 42767 36760
rect 28073 36755 28139 36758
rect 42517 36755 42583 36758
rect 42701 36755 42767 36758
rect 4208 36480 4528 36481
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 36415 4528 36416
rect 34928 36480 35248 36481
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 36415 35248 36416
rect 0 36138 800 36168
rect 1485 36138 1551 36141
rect 0 36136 1551 36138
rect 0 36080 1490 36136
rect 1546 36080 1551 36136
rect 0 36078 1551 36080
rect 0 36048 800 36078
rect 1485 36075 1551 36078
rect 19568 35936 19888 35937
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 35871 19888 35872
rect 50288 35936 50608 35937
rect 50288 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50608 35936
rect 50288 35871 50608 35872
rect 9581 35730 9647 35733
rect 57881 35730 57947 35733
rect 9581 35728 57947 35730
rect 9581 35672 9586 35728
rect 9642 35672 57886 35728
rect 57942 35672 57947 35728
rect 9581 35670 57947 35672
rect 9581 35667 9647 35670
rect 57881 35667 57947 35670
rect 58157 35458 58223 35461
rect 59200 35458 60000 35488
rect 58157 35456 60000 35458
rect 58157 35400 58162 35456
rect 58218 35400 60000 35456
rect 58157 35398 60000 35400
rect 58157 35395 58223 35398
rect 4208 35392 4528 35393
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 35327 4528 35328
rect 34928 35392 35248 35393
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 59200 35368 60000 35398
rect 34928 35327 35248 35328
rect 19568 34848 19888 34849
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 34783 19888 34784
rect 50288 34848 50608 34849
rect 50288 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50608 34848
rect 50288 34783 50608 34784
rect 4208 34304 4528 34305
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 34239 4528 34240
rect 34928 34304 35248 34305
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 34239 35248 34240
rect 19568 33760 19888 33761
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 33695 19888 33696
rect 50288 33760 50608 33761
rect 50288 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50608 33760
rect 50288 33695 50608 33696
rect 0 33418 800 33448
rect 1577 33418 1643 33421
rect 0 33416 1643 33418
rect 0 33360 1582 33416
rect 1638 33360 1643 33416
rect 0 33358 1643 33360
rect 0 33328 800 33358
rect 1577 33355 1643 33358
rect 58157 33418 58223 33421
rect 59200 33418 60000 33448
rect 58157 33416 60000 33418
rect 58157 33360 58162 33416
rect 58218 33360 60000 33416
rect 58157 33358 60000 33360
rect 58157 33355 58223 33358
rect 59200 33328 60000 33358
rect 4208 33216 4528 33217
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 33151 4528 33152
rect 34928 33216 35248 33217
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 33151 35248 33152
rect 19568 32672 19888 32673
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 32607 19888 32608
rect 50288 32672 50608 32673
rect 50288 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50608 32672
rect 50288 32607 50608 32608
rect 4208 32128 4528 32129
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 32063 4528 32064
rect 34928 32128 35248 32129
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 32063 35248 32064
rect 19568 31584 19888 31585
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 31519 19888 31520
rect 50288 31584 50608 31585
rect 50288 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50608 31584
rect 50288 31519 50608 31520
rect 0 31378 800 31408
rect 1577 31378 1643 31381
rect 0 31376 1643 31378
rect 0 31320 1582 31376
rect 1638 31320 1643 31376
rect 0 31318 1643 31320
rect 0 31288 800 31318
rect 1577 31315 1643 31318
rect 3233 31378 3299 31381
rect 54937 31378 55003 31381
rect 3233 31376 55003 31378
rect 3233 31320 3238 31376
rect 3294 31320 54942 31376
rect 54998 31320 55003 31376
rect 3233 31318 55003 31320
rect 3233 31315 3299 31318
rect 54937 31315 55003 31318
rect 57881 31378 57947 31381
rect 59200 31378 60000 31408
rect 57881 31376 60000 31378
rect 57881 31320 57886 31376
rect 57942 31320 60000 31376
rect 57881 31318 60000 31320
rect 57881 31315 57947 31318
rect 59200 31288 60000 31318
rect 4208 31040 4528 31041
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 30975 4528 30976
rect 34928 31040 35248 31041
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 30975 35248 30976
rect 19568 30496 19888 30497
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 30431 19888 30432
rect 50288 30496 50608 30497
rect 50288 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50608 30496
rect 50288 30431 50608 30432
rect 11053 30018 11119 30021
rect 18045 30018 18111 30021
rect 11053 30016 18111 30018
rect 11053 29960 11058 30016
rect 11114 29960 18050 30016
rect 18106 29960 18111 30016
rect 11053 29958 18111 29960
rect 11053 29955 11119 29958
rect 18045 29955 18111 29958
rect 4208 29952 4528 29953
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 29887 4528 29888
rect 34928 29952 35248 29953
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 29887 35248 29888
rect 19568 29408 19888 29409
rect 0 29338 800 29368
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 29343 19888 29344
rect 50288 29408 50608 29409
rect 50288 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50608 29408
rect 50288 29343 50608 29344
rect 1485 29338 1551 29341
rect 0 29336 1551 29338
rect 0 29280 1490 29336
rect 1546 29280 1551 29336
rect 0 29278 1551 29280
rect 0 29248 800 29278
rect 1485 29275 1551 29278
rect 13077 29338 13143 29341
rect 13905 29338 13971 29341
rect 16021 29338 16087 29341
rect 13077 29336 16087 29338
rect 13077 29280 13082 29336
rect 13138 29280 13910 29336
rect 13966 29280 16026 29336
rect 16082 29280 16087 29336
rect 13077 29278 16087 29280
rect 13077 29275 13143 29278
rect 13905 29275 13971 29278
rect 16021 29275 16087 29278
rect 58157 29338 58223 29341
rect 59200 29338 60000 29368
rect 58157 29336 60000 29338
rect 58157 29280 58162 29336
rect 58218 29280 60000 29336
rect 58157 29278 60000 29280
rect 58157 29275 58223 29278
rect 59200 29248 60000 29278
rect 13629 29202 13695 29205
rect 14917 29202 14983 29205
rect 13629 29200 14983 29202
rect 13629 29144 13634 29200
rect 13690 29144 14922 29200
rect 14978 29144 14983 29200
rect 13629 29142 14983 29144
rect 13629 29139 13695 29142
rect 14917 29139 14983 29142
rect 10777 29066 10843 29069
rect 13997 29066 14063 29069
rect 14641 29066 14707 29069
rect 10777 29064 14707 29066
rect 10777 29008 10782 29064
rect 10838 29008 14002 29064
rect 14058 29008 14646 29064
rect 14702 29008 14707 29064
rect 10777 29006 14707 29008
rect 10777 29003 10843 29006
rect 13997 29003 14063 29006
rect 14641 29003 14707 29006
rect 16205 29066 16271 29069
rect 19333 29066 19399 29069
rect 23289 29066 23355 29069
rect 16205 29064 23355 29066
rect 16205 29008 16210 29064
rect 16266 29008 19338 29064
rect 19394 29008 23294 29064
rect 23350 29008 23355 29064
rect 16205 29006 23355 29008
rect 16205 29003 16271 29006
rect 19333 29003 19399 29006
rect 23289 29003 23355 29006
rect 4208 28864 4528 28865
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 28799 4528 28800
rect 34928 28864 35248 28865
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 28799 35248 28800
rect 19568 28320 19888 28321
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 28255 19888 28256
rect 50288 28320 50608 28321
rect 50288 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50608 28320
rect 50288 28255 50608 28256
rect 22001 27978 22067 27981
rect 37273 27978 37339 27981
rect 22001 27976 37339 27978
rect 22001 27920 22006 27976
rect 22062 27920 37278 27976
rect 37334 27920 37339 27976
rect 22001 27918 37339 27920
rect 22001 27915 22067 27918
rect 37273 27915 37339 27918
rect 4208 27776 4528 27777
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 27711 4528 27712
rect 34928 27776 35248 27777
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 27711 35248 27712
rect 15653 27434 15719 27437
rect 19333 27434 19399 27437
rect 15653 27432 19399 27434
rect 15653 27376 15658 27432
rect 15714 27376 19338 27432
rect 19394 27376 19399 27432
rect 15653 27374 19399 27376
rect 15653 27371 15719 27374
rect 19333 27371 19399 27374
rect 0 27298 800 27328
rect 1853 27298 1919 27301
rect 0 27296 1919 27298
rect 0 27240 1858 27296
rect 1914 27240 1919 27296
rect 0 27238 1919 27240
rect 0 27208 800 27238
rect 1853 27235 1919 27238
rect 58157 27298 58223 27301
rect 59200 27298 60000 27328
rect 58157 27296 60000 27298
rect 58157 27240 58162 27296
rect 58218 27240 60000 27296
rect 58157 27238 60000 27240
rect 58157 27235 58223 27238
rect 19568 27232 19888 27233
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 27167 19888 27168
rect 50288 27232 50608 27233
rect 50288 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50608 27232
rect 59200 27208 60000 27238
rect 50288 27167 50608 27168
rect 4208 26688 4528 26689
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 26623 4528 26624
rect 34928 26688 35248 26689
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 34928 26623 35248 26624
rect 20805 26618 20871 26621
rect 21214 26618 21220 26620
rect 20805 26616 21220 26618
rect 20805 26560 20810 26616
rect 20866 26560 21220 26616
rect 20805 26558 21220 26560
rect 20805 26555 20871 26558
rect 21214 26556 21220 26558
rect 21284 26556 21290 26620
rect 18689 26346 18755 26349
rect 19701 26346 19767 26349
rect 18689 26344 19767 26346
rect 18689 26288 18694 26344
rect 18750 26288 19706 26344
rect 19762 26288 19767 26344
rect 18689 26286 19767 26288
rect 18689 26283 18755 26286
rect 19701 26283 19767 26286
rect 19568 26144 19888 26145
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 26079 19888 26080
rect 50288 26144 50608 26145
rect 50288 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50608 26144
rect 50288 26079 50608 26080
rect 23606 25876 23612 25940
rect 23676 25938 23682 25940
rect 52453 25938 52519 25941
rect 23676 25936 52519 25938
rect 23676 25880 52458 25936
rect 52514 25880 52519 25936
rect 23676 25878 52519 25880
rect 23676 25876 23682 25878
rect 52453 25875 52519 25878
rect 4208 25600 4528 25601
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 25535 4528 25536
rect 34928 25600 35248 25601
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 25535 35248 25536
rect 7465 25530 7531 25533
rect 30373 25530 30439 25533
rect 7465 25528 30439 25530
rect 7465 25472 7470 25528
rect 7526 25472 30378 25528
rect 30434 25472 30439 25528
rect 7465 25470 30439 25472
rect 7465 25467 7531 25470
rect 30373 25467 30439 25470
rect 0 25258 800 25288
rect 1853 25258 1919 25261
rect 0 25256 1919 25258
rect 0 25200 1858 25256
rect 1914 25200 1919 25256
rect 0 25198 1919 25200
rect 0 25168 800 25198
rect 1853 25195 1919 25198
rect 14733 25258 14799 25261
rect 31293 25258 31359 25261
rect 14733 25256 31359 25258
rect 14733 25200 14738 25256
rect 14794 25200 31298 25256
rect 31354 25200 31359 25256
rect 14733 25198 31359 25200
rect 14733 25195 14799 25198
rect 31293 25195 31359 25198
rect 58065 25258 58131 25261
rect 59200 25258 60000 25288
rect 58065 25256 60000 25258
rect 58065 25200 58070 25256
rect 58126 25200 60000 25256
rect 58065 25198 60000 25200
rect 58065 25195 58131 25198
rect 59200 25168 60000 25198
rect 19568 25056 19888 25057
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 24991 19888 24992
rect 50288 25056 50608 25057
rect 50288 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50608 25056
rect 50288 24991 50608 24992
rect 15193 24850 15259 24853
rect 19977 24850 20043 24853
rect 20345 24850 20411 24853
rect 15193 24848 20411 24850
rect 15193 24792 15198 24848
rect 15254 24792 19982 24848
rect 20038 24792 20350 24848
rect 20406 24792 20411 24848
rect 15193 24790 20411 24792
rect 15193 24787 15259 24790
rect 19977 24787 20043 24790
rect 20345 24787 20411 24790
rect 4208 24512 4528 24513
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 24447 4528 24448
rect 34928 24512 35248 24513
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 24447 35248 24448
rect 14733 24306 14799 24309
rect 33225 24306 33291 24309
rect 14733 24304 33291 24306
rect 14733 24248 14738 24304
rect 14794 24248 33230 24304
rect 33286 24248 33291 24304
rect 14733 24246 33291 24248
rect 14733 24243 14799 24246
rect 33225 24243 33291 24246
rect 8385 24170 8451 24173
rect 8937 24170 9003 24173
rect 56777 24170 56843 24173
rect 8385 24168 56843 24170
rect 8385 24112 8390 24168
rect 8446 24112 8942 24168
rect 8998 24112 56782 24168
rect 56838 24112 56843 24168
rect 8385 24110 56843 24112
rect 8385 24107 8451 24110
rect 8937 24107 9003 24110
rect 56777 24107 56843 24110
rect 20161 24034 20227 24037
rect 24853 24034 24919 24037
rect 20161 24032 24919 24034
rect 20161 23976 20166 24032
rect 20222 23976 24858 24032
rect 24914 23976 24919 24032
rect 20161 23974 24919 23976
rect 20161 23971 20227 23974
rect 24853 23971 24919 23974
rect 19568 23968 19888 23969
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 23903 19888 23904
rect 50288 23968 50608 23969
rect 50288 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50608 23968
rect 50288 23903 50608 23904
rect 10777 23490 10843 23493
rect 15101 23490 15167 23493
rect 10777 23488 15167 23490
rect 10777 23432 10782 23488
rect 10838 23432 15106 23488
rect 15162 23432 15167 23488
rect 10777 23430 15167 23432
rect 10777 23427 10843 23430
rect 15101 23427 15167 23430
rect 23422 23428 23428 23492
rect 23492 23490 23498 23492
rect 29637 23490 29703 23493
rect 23492 23488 29703 23490
rect 23492 23432 29642 23488
rect 29698 23432 29703 23488
rect 23492 23430 29703 23432
rect 23492 23428 23498 23430
rect 29637 23427 29703 23430
rect 4208 23424 4528 23425
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 23359 4528 23360
rect 34928 23424 35248 23425
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 23359 35248 23360
rect 0 23218 800 23248
rect 1853 23218 1919 23221
rect 0 23216 1919 23218
rect 0 23160 1858 23216
rect 1914 23160 1919 23216
rect 0 23158 1919 23160
rect 0 23128 800 23158
rect 1853 23155 1919 23158
rect 57881 23218 57947 23221
rect 59200 23218 60000 23248
rect 57881 23216 60000 23218
rect 57881 23160 57886 23216
rect 57942 23160 60000 23216
rect 57881 23158 60000 23160
rect 57881 23155 57947 23158
rect 59200 23128 60000 23158
rect 2037 23082 2103 23085
rect 23381 23082 23447 23085
rect 2037 23080 23447 23082
rect 2037 23024 2042 23080
rect 2098 23024 23386 23080
rect 23442 23024 23447 23080
rect 2037 23022 23447 23024
rect 2037 23019 2103 23022
rect 23381 23019 23447 23022
rect 19568 22880 19888 22881
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 22815 19888 22816
rect 50288 22880 50608 22881
rect 50288 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50608 22880
rect 50288 22815 50608 22816
rect 15193 22674 15259 22677
rect 33501 22674 33567 22677
rect 15193 22672 33567 22674
rect 15193 22616 15198 22672
rect 15254 22616 33506 22672
rect 33562 22616 33567 22672
rect 15193 22614 33567 22616
rect 15193 22611 15259 22614
rect 33501 22611 33567 22614
rect 14457 22538 14523 22541
rect 36629 22538 36695 22541
rect 14457 22536 36695 22538
rect 14457 22480 14462 22536
rect 14518 22480 36634 22536
rect 36690 22480 36695 22536
rect 14457 22478 36695 22480
rect 14457 22475 14523 22478
rect 36629 22475 36695 22478
rect 14181 22402 14247 22405
rect 17033 22402 17099 22405
rect 14181 22400 17099 22402
rect 14181 22344 14186 22400
rect 14242 22344 17038 22400
rect 17094 22344 17099 22400
rect 14181 22342 17099 22344
rect 14181 22339 14247 22342
rect 17033 22339 17099 22342
rect 4208 22336 4528 22337
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 22271 4528 22272
rect 34928 22336 35248 22337
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 22271 35248 22272
rect 15469 22130 15535 22133
rect 23105 22130 23171 22133
rect 15469 22128 23171 22130
rect 15469 22072 15474 22128
rect 15530 22072 23110 22128
rect 23166 22072 23171 22128
rect 15469 22070 23171 22072
rect 15469 22067 15535 22070
rect 23105 22067 23171 22070
rect 19977 21858 20043 21861
rect 22093 21858 22159 21861
rect 19977 21856 22159 21858
rect 19977 21800 19982 21856
rect 20038 21800 22098 21856
rect 22154 21800 22159 21856
rect 19977 21798 22159 21800
rect 19977 21795 20043 21798
rect 22093 21795 22159 21798
rect 19568 21792 19888 21793
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 21727 19888 21728
rect 50288 21792 50608 21793
rect 50288 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50608 21792
rect 50288 21727 50608 21728
rect 9765 21586 9831 21589
rect 27613 21586 27679 21589
rect 9765 21584 27679 21586
rect 9765 21528 9770 21584
rect 9826 21528 27618 21584
rect 27674 21528 27679 21584
rect 9765 21526 27679 21528
rect 9765 21523 9831 21526
rect 27613 21523 27679 21526
rect 10501 21450 10567 21453
rect 33317 21450 33383 21453
rect 10501 21448 33383 21450
rect 10501 21392 10506 21448
rect 10562 21392 33322 21448
rect 33378 21392 33383 21448
rect 10501 21390 33383 21392
rect 10501 21387 10567 21390
rect 33317 21387 33383 21390
rect 11053 21314 11119 21317
rect 14089 21314 14155 21317
rect 11053 21312 14155 21314
rect 11053 21256 11058 21312
rect 11114 21256 14094 21312
rect 14150 21256 14155 21312
rect 11053 21254 14155 21256
rect 11053 21251 11119 21254
rect 14089 21251 14155 21254
rect 16113 21314 16179 21317
rect 19333 21314 19399 21317
rect 20345 21314 20411 21317
rect 16113 21312 20411 21314
rect 16113 21256 16118 21312
rect 16174 21256 19338 21312
rect 19394 21256 20350 21312
rect 20406 21256 20411 21312
rect 16113 21254 20411 21256
rect 16113 21251 16179 21254
rect 19333 21251 19399 21254
rect 20345 21251 20411 21254
rect 21817 21314 21883 21317
rect 22185 21314 22251 21317
rect 21817 21312 22251 21314
rect 21817 21256 21822 21312
rect 21878 21256 22190 21312
rect 22246 21256 22251 21312
rect 21817 21254 22251 21256
rect 21817 21251 21883 21254
rect 22185 21251 22251 21254
rect 4208 21248 4528 21249
rect 0 21178 800 21208
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 21183 4528 21184
rect 34928 21248 35248 21249
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 21183 35248 21184
rect 1393 21178 1459 21181
rect 0 21176 1459 21178
rect 0 21120 1398 21176
rect 1454 21120 1459 21176
rect 0 21118 1459 21120
rect 0 21088 800 21118
rect 1393 21115 1459 21118
rect 20253 21178 20319 21181
rect 30557 21178 30623 21181
rect 20253 21176 30623 21178
rect 20253 21120 20258 21176
rect 20314 21120 30562 21176
rect 30618 21120 30623 21176
rect 20253 21118 30623 21120
rect 20253 21115 20319 21118
rect 30557 21115 30623 21118
rect 15009 21042 15075 21045
rect 27337 21042 27403 21045
rect 15009 21040 27403 21042
rect 15009 20984 15014 21040
rect 15070 20984 27342 21040
rect 27398 20984 27403 21040
rect 15009 20982 27403 20984
rect 15009 20979 15075 20982
rect 27337 20979 27403 20982
rect 16481 20906 16547 20909
rect 38193 20906 38259 20909
rect 16481 20904 38259 20906
rect 16481 20848 16486 20904
rect 16542 20848 38198 20904
rect 38254 20848 38259 20904
rect 16481 20846 38259 20848
rect 16481 20843 16547 20846
rect 38193 20843 38259 20846
rect 19568 20704 19888 20705
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 20639 19888 20640
rect 50288 20704 50608 20705
rect 50288 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50608 20704
rect 50288 20639 50608 20640
rect 10409 20498 10475 20501
rect 34605 20498 34671 20501
rect 10409 20496 34671 20498
rect 10409 20440 10414 20496
rect 10470 20440 34610 20496
rect 34666 20440 34671 20496
rect 10409 20438 34671 20440
rect 10409 20435 10475 20438
rect 34605 20435 34671 20438
rect 58157 20498 58223 20501
rect 59200 20498 60000 20528
rect 58157 20496 60000 20498
rect 58157 20440 58162 20496
rect 58218 20440 60000 20496
rect 58157 20438 60000 20440
rect 58157 20435 58223 20438
rect 59200 20408 60000 20438
rect 13077 20362 13143 20365
rect 30373 20362 30439 20365
rect 13077 20360 30439 20362
rect 13077 20304 13082 20360
rect 13138 20304 30378 20360
rect 30434 20304 30439 20360
rect 13077 20302 30439 20304
rect 13077 20299 13143 20302
rect 30373 20299 30439 20302
rect 15745 20226 15811 20229
rect 16297 20226 16363 20229
rect 26509 20226 26575 20229
rect 15745 20224 26575 20226
rect 15745 20168 15750 20224
rect 15806 20168 16302 20224
rect 16358 20168 26514 20224
rect 26570 20168 26575 20224
rect 15745 20166 26575 20168
rect 15745 20163 15811 20166
rect 16297 20163 16363 20166
rect 26509 20163 26575 20166
rect 4208 20160 4528 20161
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 20095 4528 20096
rect 34928 20160 35248 20161
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 20095 35248 20096
rect 19568 19616 19888 19617
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 19551 19888 19552
rect 50288 19616 50608 19617
rect 50288 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50608 19616
rect 50288 19551 50608 19552
rect 15929 19410 15995 19413
rect 43345 19410 43411 19413
rect 15929 19408 43411 19410
rect 15929 19352 15934 19408
rect 15990 19352 43350 19408
rect 43406 19352 43411 19408
rect 15929 19350 43411 19352
rect 15929 19347 15995 19350
rect 43345 19347 43411 19350
rect 23381 19274 23447 19277
rect 38009 19274 38075 19277
rect 23381 19272 38075 19274
rect 23381 19216 23386 19272
rect 23442 19216 38014 19272
rect 38070 19216 38075 19272
rect 23381 19214 38075 19216
rect 23381 19211 23447 19214
rect 38009 19211 38075 19214
rect 0 19138 800 19168
rect 1393 19138 1459 19141
rect 0 19136 1459 19138
rect 0 19080 1398 19136
rect 1454 19080 1459 19136
rect 0 19078 1459 19080
rect 0 19048 800 19078
rect 1393 19075 1459 19078
rect 4208 19072 4528 19073
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 19007 4528 19008
rect 34928 19072 35248 19073
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 34928 19007 35248 19008
rect 2681 18866 2747 18869
rect 23606 18866 23612 18868
rect 2681 18864 23612 18866
rect 2681 18808 2686 18864
rect 2742 18808 23612 18864
rect 2681 18806 23612 18808
rect 2681 18803 2747 18806
rect 23606 18804 23612 18806
rect 23676 18804 23682 18868
rect 14917 18730 14983 18733
rect 41781 18730 41847 18733
rect 14917 18728 41847 18730
rect 14917 18672 14922 18728
rect 14978 18672 41786 18728
rect 41842 18672 41847 18728
rect 14917 18670 41847 18672
rect 14917 18667 14983 18670
rect 41781 18667 41847 18670
rect 19568 18528 19888 18529
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 18463 19888 18464
rect 50288 18528 50608 18529
rect 50288 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50608 18528
rect 50288 18463 50608 18464
rect 58065 18458 58131 18461
rect 59200 18458 60000 18488
rect 58065 18456 60000 18458
rect 58065 18400 58070 18456
rect 58126 18400 60000 18456
rect 58065 18398 60000 18400
rect 58065 18395 58131 18398
rect 59200 18368 60000 18398
rect 24117 18322 24183 18325
rect 25037 18322 25103 18325
rect 24117 18320 25103 18322
rect 24117 18264 24122 18320
rect 24178 18264 25042 18320
rect 25098 18264 25103 18320
rect 24117 18262 25103 18264
rect 24117 18259 24183 18262
rect 25037 18259 25103 18262
rect 4208 17984 4528 17985
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 17919 4528 17920
rect 34928 17984 35248 17985
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 17919 35248 17920
rect 15561 17642 15627 17645
rect 50153 17642 50219 17645
rect 15561 17640 50219 17642
rect 15561 17584 15566 17640
rect 15622 17584 50158 17640
rect 50214 17584 50219 17640
rect 15561 17582 50219 17584
rect 15561 17579 15627 17582
rect 50153 17579 50219 17582
rect 20805 17506 20871 17509
rect 40217 17506 40283 17509
rect 20805 17504 40283 17506
rect 20805 17448 20810 17504
rect 20866 17448 40222 17504
rect 40278 17448 40283 17504
rect 20805 17446 40283 17448
rect 20805 17443 20871 17446
rect 40217 17443 40283 17446
rect 19568 17440 19888 17441
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 17375 19888 17376
rect 50288 17440 50608 17441
rect 50288 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50608 17440
rect 50288 17375 50608 17376
rect 26233 17098 26299 17101
rect 38745 17098 38811 17101
rect 26233 17096 38811 17098
rect 26233 17040 26238 17096
rect 26294 17040 38750 17096
rect 38806 17040 38811 17096
rect 26233 17038 38811 17040
rect 26233 17035 26299 17038
rect 38745 17035 38811 17038
rect 4208 16896 4528 16897
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 16831 4528 16832
rect 34928 16896 35248 16897
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 34928 16831 35248 16832
rect 13537 16826 13603 16829
rect 23422 16826 23428 16828
rect 13537 16824 23428 16826
rect 13537 16768 13542 16824
rect 13598 16768 23428 16824
rect 13537 16766 23428 16768
rect 13537 16763 13603 16766
rect 23422 16764 23428 16766
rect 23492 16764 23498 16828
rect 19701 16690 19767 16693
rect 40033 16690 40099 16693
rect 19701 16688 40099 16690
rect 19701 16632 19706 16688
rect 19762 16632 40038 16688
rect 40094 16632 40099 16688
rect 19701 16630 40099 16632
rect 19701 16627 19767 16630
rect 40033 16627 40099 16630
rect 0 16418 800 16448
rect 1853 16418 1919 16421
rect 0 16416 1919 16418
rect 0 16360 1858 16416
rect 1914 16360 1919 16416
rect 0 16358 1919 16360
rect 0 16328 800 16358
rect 1853 16355 1919 16358
rect 58157 16418 58223 16421
rect 59200 16418 60000 16448
rect 58157 16416 60000 16418
rect 58157 16360 58162 16416
rect 58218 16360 60000 16416
rect 58157 16358 60000 16360
rect 58157 16355 58223 16358
rect 19568 16352 19888 16353
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 16287 19888 16288
rect 50288 16352 50608 16353
rect 50288 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50608 16352
rect 59200 16328 60000 16358
rect 50288 16287 50608 16288
rect 7557 16146 7623 16149
rect 11881 16146 11947 16149
rect 7557 16144 11947 16146
rect 7557 16088 7562 16144
rect 7618 16088 11886 16144
rect 11942 16088 11947 16144
rect 7557 16086 11947 16088
rect 7557 16083 7623 16086
rect 11881 16083 11947 16086
rect 20621 16010 20687 16013
rect 39849 16010 39915 16013
rect 20621 16008 39915 16010
rect 20621 15952 20626 16008
rect 20682 15952 39854 16008
rect 39910 15952 39915 16008
rect 20621 15950 39915 15952
rect 20621 15947 20687 15950
rect 39849 15947 39915 15950
rect 13721 15874 13787 15877
rect 31017 15874 31083 15877
rect 13721 15872 31083 15874
rect 13721 15816 13726 15872
rect 13782 15816 31022 15872
rect 31078 15816 31083 15872
rect 13721 15814 31083 15816
rect 13721 15811 13787 15814
rect 31017 15811 31083 15814
rect 4208 15808 4528 15809
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 15743 4528 15744
rect 34928 15808 35248 15809
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 34928 15743 35248 15744
rect 21081 15738 21147 15741
rect 24761 15738 24827 15741
rect 21081 15736 24827 15738
rect 21081 15680 21086 15736
rect 21142 15680 24766 15736
rect 24822 15680 24827 15736
rect 21081 15678 24827 15680
rect 21081 15675 21147 15678
rect 24761 15675 24827 15678
rect 33041 15602 33107 15605
rect 53557 15602 53623 15605
rect 33041 15600 53623 15602
rect 33041 15544 33046 15600
rect 33102 15544 53562 15600
rect 53618 15544 53623 15600
rect 33041 15542 53623 15544
rect 33041 15539 33107 15542
rect 53557 15539 53623 15542
rect 15193 15466 15259 15469
rect 41965 15466 42031 15469
rect 15193 15464 42031 15466
rect 15193 15408 15198 15464
rect 15254 15408 41970 15464
rect 42026 15408 42031 15464
rect 15193 15406 42031 15408
rect 15193 15403 15259 15406
rect 41965 15403 42031 15406
rect 21214 15268 21220 15332
rect 21284 15330 21290 15332
rect 23381 15330 23447 15333
rect 21284 15328 23447 15330
rect 21284 15272 23386 15328
rect 23442 15272 23447 15328
rect 21284 15270 23447 15272
rect 21284 15268 21290 15270
rect 23381 15267 23447 15270
rect 19568 15264 19888 15265
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 15199 19888 15200
rect 50288 15264 50608 15265
rect 50288 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50608 15264
rect 50288 15199 50608 15200
rect 20713 15194 20779 15197
rect 40033 15194 40099 15197
rect 20713 15192 40099 15194
rect 20713 15136 20718 15192
rect 20774 15136 40038 15192
rect 40094 15136 40099 15192
rect 20713 15134 40099 15136
rect 20713 15131 20779 15134
rect 40033 15131 40099 15134
rect 15837 15058 15903 15061
rect 19517 15058 19583 15061
rect 15837 15056 19583 15058
rect 15837 15000 15842 15056
rect 15898 15000 19522 15056
rect 19578 15000 19583 15056
rect 15837 14998 19583 15000
rect 15837 14995 15903 14998
rect 19517 14995 19583 14998
rect 15561 14922 15627 14925
rect 16849 14922 16915 14925
rect 15561 14920 16915 14922
rect 15561 14864 15566 14920
rect 15622 14864 16854 14920
rect 16910 14864 16915 14920
rect 15561 14862 16915 14864
rect 15561 14859 15627 14862
rect 16849 14859 16915 14862
rect 17677 14922 17743 14925
rect 49785 14922 49851 14925
rect 17677 14920 49851 14922
rect 17677 14864 17682 14920
rect 17738 14864 49790 14920
rect 49846 14864 49851 14920
rect 17677 14862 49851 14864
rect 17677 14859 17743 14862
rect 49785 14859 49851 14862
rect 12065 14786 12131 14789
rect 12617 14786 12683 14789
rect 20713 14786 20779 14789
rect 12065 14784 20779 14786
rect 12065 14728 12070 14784
rect 12126 14728 12622 14784
rect 12678 14728 20718 14784
rect 20774 14728 20779 14784
rect 12065 14726 20779 14728
rect 12065 14723 12131 14726
rect 12617 14723 12683 14726
rect 20713 14723 20779 14726
rect 4208 14720 4528 14721
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 14655 4528 14656
rect 34928 14720 35248 14721
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 14655 35248 14656
rect 0 14378 800 14408
rect 1393 14378 1459 14381
rect 0 14376 1459 14378
rect 0 14320 1398 14376
rect 1454 14320 1459 14376
rect 0 14318 1459 14320
rect 0 14288 800 14318
rect 1393 14315 1459 14318
rect 19333 14378 19399 14381
rect 31385 14378 31451 14381
rect 19333 14376 31451 14378
rect 19333 14320 19338 14376
rect 19394 14320 31390 14376
rect 31446 14320 31451 14376
rect 19333 14318 31451 14320
rect 19333 14315 19399 14318
rect 31385 14315 31451 14318
rect 32949 14378 33015 14381
rect 44357 14378 44423 14381
rect 32949 14376 44423 14378
rect 32949 14320 32954 14376
rect 33010 14320 44362 14376
rect 44418 14320 44423 14376
rect 32949 14318 44423 14320
rect 32949 14315 33015 14318
rect 44357 14315 44423 14318
rect 58065 14378 58131 14381
rect 59200 14378 60000 14408
rect 58065 14376 60000 14378
rect 58065 14320 58070 14376
rect 58126 14320 60000 14376
rect 58065 14318 60000 14320
rect 58065 14315 58131 14318
rect 59200 14288 60000 14318
rect 19568 14176 19888 14177
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 14111 19888 14112
rect 50288 14176 50608 14177
rect 50288 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50608 14176
rect 50288 14111 50608 14112
rect 15837 13970 15903 13973
rect 16297 13970 16363 13973
rect 15837 13968 16363 13970
rect 15837 13912 15842 13968
rect 15898 13912 16302 13968
rect 16358 13912 16363 13968
rect 15837 13910 16363 13912
rect 15837 13907 15903 13910
rect 16297 13907 16363 13910
rect 20897 13834 20963 13837
rect 21817 13834 21883 13837
rect 20897 13832 21883 13834
rect 20897 13776 20902 13832
rect 20958 13776 21822 13832
rect 21878 13776 21883 13832
rect 20897 13774 21883 13776
rect 20897 13771 20963 13774
rect 21817 13771 21883 13774
rect 4208 13632 4528 13633
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 13567 4528 13568
rect 34928 13632 35248 13633
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 13567 35248 13568
rect 19977 13290 20043 13293
rect 46657 13290 46723 13293
rect 19977 13288 46723 13290
rect 19977 13232 19982 13288
rect 20038 13232 46662 13288
rect 46718 13232 46723 13288
rect 19977 13230 46723 13232
rect 19977 13227 20043 13230
rect 46657 13227 46723 13230
rect 22461 13154 22527 13157
rect 30281 13154 30347 13157
rect 22461 13152 30347 13154
rect 22461 13096 22466 13152
rect 22522 13096 30286 13152
rect 30342 13096 30347 13152
rect 22461 13094 30347 13096
rect 22461 13091 22527 13094
rect 30281 13091 30347 13094
rect 19568 13088 19888 13089
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 13023 19888 13024
rect 50288 13088 50608 13089
rect 50288 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50608 13088
rect 50288 13023 50608 13024
rect 16481 12746 16547 12749
rect 37549 12746 37615 12749
rect 16481 12744 37615 12746
rect 16481 12688 16486 12744
rect 16542 12688 37554 12744
rect 37610 12688 37615 12744
rect 16481 12686 37615 12688
rect 16481 12683 16547 12686
rect 37549 12683 37615 12686
rect 10961 12610 11027 12613
rect 23473 12610 23539 12613
rect 10961 12608 23539 12610
rect 10961 12552 10966 12608
rect 11022 12552 23478 12608
rect 23534 12552 23539 12608
rect 10961 12550 23539 12552
rect 10961 12547 11027 12550
rect 23473 12547 23539 12550
rect 4208 12544 4528 12545
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 12479 4528 12480
rect 34928 12544 35248 12545
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 12479 35248 12480
rect 13537 12474 13603 12477
rect 23013 12474 23079 12477
rect 31569 12474 31635 12477
rect 13537 12472 31635 12474
rect 13537 12416 13542 12472
rect 13598 12416 23018 12472
rect 23074 12416 31574 12472
rect 31630 12416 31635 12472
rect 13537 12414 31635 12416
rect 13537 12411 13603 12414
rect 0 12338 800 12368
rect 17174 12341 17234 12414
rect 23013 12411 23079 12414
rect 31569 12411 31635 12414
rect 1393 12338 1459 12341
rect 0 12336 1459 12338
rect 0 12280 1398 12336
rect 1454 12280 1459 12336
rect 0 12278 1459 12280
rect 17174 12336 17283 12341
rect 17174 12280 17222 12336
rect 17278 12280 17283 12336
rect 17174 12278 17283 12280
rect 0 12248 800 12278
rect 1393 12275 1459 12278
rect 17217 12275 17283 12278
rect 21449 12338 21515 12341
rect 25221 12338 25287 12341
rect 21449 12336 25287 12338
rect 21449 12280 21454 12336
rect 21510 12280 25226 12336
rect 25282 12280 25287 12336
rect 21449 12278 25287 12280
rect 21449 12275 21515 12278
rect 25221 12275 25287 12278
rect 58157 12338 58223 12341
rect 59200 12338 60000 12368
rect 58157 12336 60000 12338
rect 58157 12280 58162 12336
rect 58218 12280 60000 12336
rect 58157 12278 60000 12280
rect 58157 12275 58223 12278
rect 59200 12248 60000 12278
rect 20621 12202 20687 12205
rect 40309 12202 40375 12205
rect 20621 12200 40375 12202
rect 20621 12144 20626 12200
rect 20682 12144 40314 12200
rect 40370 12144 40375 12200
rect 20621 12142 40375 12144
rect 20621 12139 20687 12142
rect 40309 12139 40375 12142
rect 19568 12000 19888 12001
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 11935 19888 11936
rect 50288 12000 50608 12001
rect 50288 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50608 12000
rect 50288 11935 50608 11936
rect 23473 11794 23539 11797
rect 56041 11794 56107 11797
rect 23473 11792 56107 11794
rect 23473 11736 23478 11792
rect 23534 11736 56046 11792
rect 56102 11736 56107 11792
rect 23473 11734 56107 11736
rect 23473 11731 23539 11734
rect 56041 11731 56107 11734
rect 7097 11658 7163 11661
rect 52729 11658 52795 11661
rect 7097 11656 52795 11658
rect 7097 11600 7102 11656
rect 7158 11600 52734 11656
rect 52790 11600 52795 11656
rect 7097 11598 52795 11600
rect 7097 11595 7163 11598
rect 52729 11595 52795 11598
rect 4208 11456 4528 11457
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 11391 4528 11392
rect 34928 11456 35248 11457
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 11391 35248 11392
rect 23013 11250 23079 11253
rect 37365 11250 37431 11253
rect 23013 11248 37431 11250
rect 23013 11192 23018 11248
rect 23074 11192 37370 11248
rect 37426 11192 37431 11248
rect 23013 11190 37431 11192
rect 23013 11187 23079 11190
rect 37365 11187 37431 11190
rect 21909 10978 21975 10981
rect 24393 10978 24459 10981
rect 21909 10976 24459 10978
rect 21909 10920 21914 10976
rect 21970 10920 24398 10976
rect 24454 10920 24459 10976
rect 21909 10918 24459 10920
rect 21909 10915 21975 10918
rect 24393 10915 24459 10918
rect 19568 10912 19888 10913
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 10847 19888 10848
rect 50288 10912 50608 10913
rect 50288 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50608 10912
rect 50288 10847 50608 10848
rect 10869 10706 10935 10709
rect 51717 10706 51783 10709
rect 10869 10704 51783 10706
rect 10869 10648 10874 10704
rect 10930 10648 51722 10704
rect 51778 10648 51783 10704
rect 10869 10646 51783 10648
rect 10869 10643 10935 10646
rect 51717 10643 51783 10646
rect 10685 10570 10751 10573
rect 26877 10570 26943 10573
rect 10685 10568 26943 10570
rect 10685 10512 10690 10568
rect 10746 10512 26882 10568
rect 26938 10512 26943 10568
rect 10685 10510 26943 10512
rect 10685 10507 10751 10510
rect 26877 10507 26943 10510
rect 4208 10368 4528 10369
rect 0 10298 800 10328
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 10303 4528 10304
rect 34928 10368 35248 10369
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 10303 35248 10304
rect 1393 10298 1459 10301
rect 0 10296 1459 10298
rect 0 10240 1398 10296
rect 1454 10240 1459 10296
rect 0 10238 1459 10240
rect 0 10208 800 10238
rect 1393 10235 1459 10238
rect 58065 10298 58131 10301
rect 59200 10298 60000 10328
rect 58065 10296 60000 10298
rect 58065 10240 58070 10296
rect 58126 10240 60000 10296
rect 58065 10238 60000 10240
rect 58065 10235 58131 10238
rect 59200 10208 60000 10238
rect 10225 10162 10291 10165
rect 47761 10162 47827 10165
rect 10225 10160 47827 10162
rect 10225 10104 10230 10160
rect 10286 10104 47766 10160
rect 47822 10104 47827 10160
rect 10225 10102 47827 10104
rect 10225 10099 10291 10102
rect 47761 10099 47827 10102
rect 9857 10026 9923 10029
rect 51165 10026 51231 10029
rect 9857 10024 51231 10026
rect 9857 9968 9862 10024
rect 9918 9968 51170 10024
rect 51226 9968 51231 10024
rect 9857 9966 51231 9968
rect 9857 9963 9923 9966
rect 51165 9963 51231 9966
rect 24025 9890 24091 9893
rect 35341 9890 35407 9893
rect 24025 9888 35407 9890
rect 24025 9832 24030 9888
rect 24086 9832 35346 9888
rect 35402 9832 35407 9888
rect 24025 9830 35407 9832
rect 24025 9827 24091 9830
rect 35341 9827 35407 9830
rect 19568 9824 19888 9825
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 9759 19888 9760
rect 50288 9824 50608 9825
rect 50288 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50608 9824
rect 50288 9759 50608 9760
rect 19333 9618 19399 9621
rect 22645 9618 22711 9621
rect 26325 9618 26391 9621
rect 19333 9616 26391 9618
rect 19333 9560 19338 9616
rect 19394 9560 22650 9616
rect 22706 9560 26330 9616
rect 26386 9560 26391 9616
rect 19333 9558 26391 9560
rect 19333 9555 19399 9558
rect 22645 9555 22711 9558
rect 26325 9555 26391 9558
rect 29821 9618 29887 9621
rect 30741 9618 30807 9621
rect 29821 9616 30807 9618
rect 29821 9560 29826 9616
rect 29882 9560 30746 9616
rect 30802 9560 30807 9616
rect 29821 9558 30807 9560
rect 29821 9555 29887 9558
rect 30741 9555 30807 9558
rect 9581 9482 9647 9485
rect 35893 9482 35959 9485
rect 9581 9480 35959 9482
rect 9581 9424 9586 9480
rect 9642 9424 35898 9480
rect 35954 9424 35959 9480
rect 9581 9422 35959 9424
rect 9581 9419 9647 9422
rect 35893 9419 35959 9422
rect 20713 9346 20779 9349
rect 24025 9346 24091 9349
rect 20713 9344 24091 9346
rect 20713 9288 20718 9344
rect 20774 9288 24030 9344
rect 24086 9288 24091 9344
rect 20713 9286 24091 9288
rect 20713 9283 20779 9286
rect 24025 9283 24091 9286
rect 28349 9346 28415 9349
rect 28901 9346 28967 9349
rect 28349 9344 28967 9346
rect 28349 9288 28354 9344
rect 28410 9288 28906 9344
rect 28962 9288 28967 9344
rect 28349 9286 28967 9288
rect 28349 9283 28415 9286
rect 28901 9283 28967 9286
rect 4208 9280 4528 9281
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 9215 4528 9216
rect 34928 9280 35248 9281
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 9215 35248 9216
rect 17769 9210 17835 9213
rect 31017 9210 31083 9213
rect 17769 9208 31083 9210
rect 17769 9152 17774 9208
rect 17830 9152 31022 9208
rect 31078 9152 31083 9208
rect 17769 9150 31083 9152
rect 17769 9147 17835 9150
rect 31017 9147 31083 9150
rect 17493 9074 17559 9077
rect 27797 9074 27863 9077
rect 17493 9072 27863 9074
rect 17493 9016 17498 9072
rect 17554 9016 27802 9072
rect 27858 9016 27863 9072
rect 17493 9014 27863 9016
rect 17493 9011 17559 9014
rect 27797 9011 27863 9014
rect 10041 8938 10107 8941
rect 39113 8938 39179 8941
rect 10041 8936 39179 8938
rect 10041 8880 10046 8936
rect 10102 8880 39118 8936
rect 39174 8880 39179 8936
rect 10041 8878 39179 8880
rect 10041 8875 10107 8878
rect 39113 8875 39179 8878
rect 19568 8736 19888 8737
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 8671 19888 8672
rect 50288 8736 50608 8737
rect 50288 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50608 8736
rect 50288 8671 50608 8672
rect 0 8258 800 8288
rect 1485 8258 1551 8261
rect 0 8256 1551 8258
rect 0 8200 1490 8256
rect 1546 8200 1551 8256
rect 0 8198 1551 8200
rect 0 8168 800 8198
rect 1485 8195 1551 8198
rect 58065 8258 58131 8261
rect 59200 8258 60000 8288
rect 58065 8256 60000 8258
rect 58065 8200 58070 8256
rect 58126 8200 60000 8256
rect 58065 8198 60000 8200
rect 58065 8195 58131 8198
rect 4208 8192 4528 8193
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 8127 4528 8128
rect 34928 8192 35248 8193
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 59200 8168 60000 8198
rect 34928 8127 35248 8128
rect 5349 7850 5415 7853
rect 57513 7850 57579 7853
rect 5349 7848 57579 7850
rect 5349 7792 5354 7848
rect 5410 7792 57518 7848
rect 57574 7792 57579 7848
rect 5349 7790 57579 7792
rect 5349 7787 5415 7790
rect 57513 7787 57579 7790
rect 19568 7648 19888 7649
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 7583 19888 7584
rect 50288 7648 50608 7649
rect 50288 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50608 7648
rect 50288 7583 50608 7584
rect 13721 7306 13787 7309
rect 39665 7306 39731 7309
rect 13721 7304 39731 7306
rect 13721 7248 13726 7304
rect 13782 7248 39670 7304
rect 39726 7248 39731 7304
rect 13721 7246 39731 7248
rect 13721 7243 13787 7246
rect 39665 7243 39731 7246
rect 4208 7104 4528 7105
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 7039 4528 7040
rect 34928 7104 35248 7105
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 7039 35248 7040
rect 8661 6762 8727 6765
rect 56777 6762 56843 6765
rect 8661 6760 56843 6762
rect 8661 6704 8666 6760
rect 8722 6704 56782 6760
rect 56838 6704 56843 6760
rect 8661 6702 56843 6704
rect 8661 6699 8727 6702
rect 56777 6699 56843 6702
rect 19568 6560 19888 6561
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 6495 19888 6496
rect 50288 6560 50608 6561
rect 50288 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50608 6560
rect 50288 6495 50608 6496
rect 0 6218 800 6248
rect 1577 6218 1643 6221
rect 0 6216 1643 6218
rect 0 6160 1582 6216
rect 1638 6160 1643 6216
rect 0 6158 1643 6160
rect 0 6128 800 6158
rect 1577 6155 1643 6158
rect 58065 6218 58131 6221
rect 59200 6218 60000 6248
rect 58065 6216 60000 6218
rect 58065 6160 58070 6216
rect 58126 6160 60000 6216
rect 58065 6158 60000 6160
rect 58065 6155 58131 6158
rect 59200 6128 60000 6158
rect 4208 6016 4528 6017
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 5951 4528 5952
rect 34928 6016 35248 6017
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 5951 35248 5952
rect 19568 5472 19888 5473
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 5407 19888 5408
rect 50288 5472 50608 5473
rect 50288 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50608 5472
rect 50288 5407 50608 5408
rect 4208 4928 4528 4929
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 4863 4528 4864
rect 34928 4928 35248 4929
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 4863 35248 4864
rect 19568 4384 19888 4385
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 4319 19888 4320
rect 50288 4384 50608 4385
rect 50288 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50608 4384
rect 50288 4319 50608 4320
rect 0 4178 800 4208
rect 1485 4178 1551 4181
rect 0 4176 1551 4178
rect 0 4120 1490 4176
rect 1546 4120 1551 4176
rect 0 4118 1551 4120
rect 0 4088 800 4118
rect 1485 4115 1551 4118
rect 4208 3840 4528 3841
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 3775 4528 3776
rect 34928 3840 35248 3841
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 3775 35248 3776
rect 58065 3498 58131 3501
rect 59200 3498 60000 3528
rect 58065 3496 60000 3498
rect 58065 3440 58070 3496
rect 58126 3440 60000 3496
rect 58065 3438 60000 3440
rect 58065 3435 58131 3438
rect 59200 3408 60000 3438
rect 19568 3296 19888 3297
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 3231 19888 3232
rect 50288 3296 50608 3297
rect 50288 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50608 3296
rect 50288 3231 50608 3232
rect 18045 3090 18111 3093
rect 23933 3090 23999 3093
rect 18045 3088 23999 3090
rect 18045 3032 18050 3088
rect 18106 3032 23938 3088
rect 23994 3032 23999 3088
rect 18045 3030 23999 3032
rect 18045 3027 18111 3030
rect 23933 3027 23999 3030
rect 24301 3090 24367 3093
rect 26877 3090 26943 3093
rect 24301 3088 26943 3090
rect 24301 3032 24306 3088
rect 24362 3032 26882 3088
rect 26938 3032 26943 3088
rect 24301 3030 26943 3032
rect 24301 3027 24367 3030
rect 26877 3027 26943 3030
rect 4208 2752 4528 2753
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2687 4528 2688
rect 34928 2752 35248 2753
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2687 35248 2688
rect 19568 2208 19888 2209
rect 0 2138 800 2168
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2143 19888 2144
rect 50288 2208 50608 2209
rect 50288 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50608 2208
rect 50288 2143 50608 2144
rect 1393 2138 1459 2141
rect 0 2136 1459 2138
rect 0 2080 1398 2136
rect 1454 2080 1459 2136
rect 0 2078 1459 2080
rect 0 2048 800 2078
rect 1393 2075 1459 2078
rect 57237 1458 57303 1461
rect 59200 1458 60000 1488
rect 57237 1456 60000 1458
rect 57237 1400 57242 1456
rect 57298 1400 60000 1456
rect 57237 1398 60000 1400
rect 57237 1395 57303 1398
rect 59200 1368 60000 1398
<< via3 >>
rect 4216 37564 4280 37568
rect 4216 37508 4220 37564
rect 4220 37508 4276 37564
rect 4276 37508 4280 37564
rect 4216 37504 4280 37508
rect 4296 37564 4360 37568
rect 4296 37508 4300 37564
rect 4300 37508 4356 37564
rect 4356 37508 4360 37564
rect 4296 37504 4360 37508
rect 4376 37564 4440 37568
rect 4376 37508 4380 37564
rect 4380 37508 4436 37564
rect 4436 37508 4440 37564
rect 4376 37504 4440 37508
rect 4456 37564 4520 37568
rect 4456 37508 4460 37564
rect 4460 37508 4516 37564
rect 4516 37508 4520 37564
rect 4456 37504 4520 37508
rect 34936 37564 35000 37568
rect 34936 37508 34940 37564
rect 34940 37508 34996 37564
rect 34996 37508 35000 37564
rect 34936 37504 35000 37508
rect 35016 37564 35080 37568
rect 35016 37508 35020 37564
rect 35020 37508 35076 37564
rect 35076 37508 35080 37564
rect 35016 37504 35080 37508
rect 35096 37564 35160 37568
rect 35096 37508 35100 37564
rect 35100 37508 35156 37564
rect 35156 37508 35160 37564
rect 35096 37504 35160 37508
rect 35176 37564 35240 37568
rect 35176 37508 35180 37564
rect 35180 37508 35236 37564
rect 35236 37508 35240 37564
rect 35176 37504 35240 37508
rect 19576 37020 19640 37024
rect 19576 36964 19580 37020
rect 19580 36964 19636 37020
rect 19636 36964 19640 37020
rect 19576 36960 19640 36964
rect 19656 37020 19720 37024
rect 19656 36964 19660 37020
rect 19660 36964 19716 37020
rect 19716 36964 19720 37020
rect 19656 36960 19720 36964
rect 19736 37020 19800 37024
rect 19736 36964 19740 37020
rect 19740 36964 19796 37020
rect 19796 36964 19800 37020
rect 19736 36960 19800 36964
rect 19816 37020 19880 37024
rect 19816 36964 19820 37020
rect 19820 36964 19876 37020
rect 19876 36964 19880 37020
rect 19816 36960 19880 36964
rect 50296 37020 50360 37024
rect 50296 36964 50300 37020
rect 50300 36964 50356 37020
rect 50356 36964 50360 37020
rect 50296 36960 50360 36964
rect 50376 37020 50440 37024
rect 50376 36964 50380 37020
rect 50380 36964 50436 37020
rect 50436 36964 50440 37020
rect 50376 36960 50440 36964
rect 50456 37020 50520 37024
rect 50456 36964 50460 37020
rect 50460 36964 50516 37020
rect 50516 36964 50520 37020
rect 50456 36960 50520 36964
rect 50536 37020 50600 37024
rect 50536 36964 50540 37020
rect 50540 36964 50596 37020
rect 50596 36964 50600 37020
rect 50536 36960 50600 36964
rect 4216 36476 4280 36480
rect 4216 36420 4220 36476
rect 4220 36420 4276 36476
rect 4276 36420 4280 36476
rect 4216 36416 4280 36420
rect 4296 36476 4360 36480
rect 4296 36420 4300 36476
rect 4300 36420 4356 36476
rect 4356 36420 4360 36476
rect 4296 36416 4360 36420
rect 4376 36476 4440 36480
rect 4376 36420 4380 36476
rect 4380 36420 4436 36476
rect 4436 36420 4440 36476
rect 4376 36416 4440 36420
rect 4456 36476 4520 36480
rect 4456 36420 4460 36476
rect 4460 36420 4516 36476
rect 4516 36420 4520 36476
rect 4456 36416 4520 36420
rect 34936 36476 35000 36480
rect 34936 36420 34940 36476
rect 34940 36420 34996 36476
rect 34996 36420 35000 36476
rect 34936 36416 35000 36420
rect 35016 36476 35080 36480
rect 35016 36420 35020 36476
rect 35020 36420 35076 36476
rect 35076 36420 35080 36476
rect 35016 36416 35080 36420
rect 35096 36476 35160 36480
rect 35096 36420 35100 36476
rect 35100 36420 35156 36476
rect 35156 36420 35160 36476
rect 35096 36416 35160 36420
rect 35176 36476 35240 36480
rect 35176 36420 35180 36476
rect 35180 36420 35236 36476
rect 35236 36420 35240 36476
rect 35176 36416 35240 36420
rect 19576 35932 19640 35936
rect 19576 35876 19580 35932
rect 19580 35876 19636 35932
rect 19636 35876 19640 35932
rect 19576 35872 19640 35876
rect 19656 35932 19720 35936
rect 19656 35876 19660 35932
rect 19660 35876 19716 35932
rect 19716 35876 19720 35932
rect 19656 35872 19720 35876
rect 19736 35932 19800 35936
rect 19736 35876 19740 35932
rect 19740 35876 19796 35932
rect 19796 35876 19800 35932
rect 19736 35872 19800 35876
rect 19816 35932 19880 35936
rect 19816 35876 19820 35932
rect 19820 35876 19876 35932
rect 19876 35876 19880 35932
rect 19816 35872 19880 35876
rect 50296 35932 50360 35936
rect 50296 35876 50300 35932
rect 50300 35876 50356 35932
rect 50356 35876 50360 35932
rect 50296 35872 50360 35876
rect 50376 35932 50440 35936
rect 50376 35876 50380 35932
rect 50380 35876 50436 35932
rect 50436 35876 50440 35932
rect 50376 35872 50440 35876
rect 50456 35932 50520 35936
rect 50456 35876 50460 35932
rect 50460 35876 50516 35932
rect 50516 35876 50520 35932
rect 50456 35872 50520 35876
rect 50536 35932 50600 35936
rect 50536 35876 50540 35932
rect 50540 35876 50596 35932
rect 50596 35876 50600 35932
rect 50536 35872 50600 35876
rect 4216 35388 4280 35392
rect 4216 35332 4220 35388
rect 4220 35332 4276 35388
rect 4276 35332 4280 35388
rect 4216 35328 4280 35332
rect 4296 35388 4360 35392
rect 4296 35332 4300 35388
rect 4300 35332 4356 35388
rect 4356 35332 4360 35388
rect 4296 35328 4360 35332
rect 4376 35388 4440 35392
rect 4376 35332 4380 35388
rect 4380 35332 4436 35388
rect 4436 35332 4440 35388
rect 4376 35328 4440 35332
rect 4456 35388 4520 35392
rect 4456 35332 4460 35388
rect 4460 35332 4516 35388
rect 4516 35332 4520 35388
rect 4456 35328 4520 35332
rect 34936 35388 35000 35392
rect 34936 35332 34940 35388
rect 34940 35332 34996 35388
rect 34996 35332 35000 35388
rect 34936 35328 35000 35332
rect 35016 35388 35080 35392
rect 35016 35332 35020 35388
rect 35020 35332 35076 35388
rect 35076 35332 35080 35388
rect 35016 35328 35080 35332
rect 35096 35388 35160 35392
rect 35096 35332 35100 35388
rect 35100 35332 35156 35388
rect 35156 35332 35160 35388
rect 35096 35328 35160 35332
rect 35176 35388 35240 35392
rect 35176 35332 35180 35388
rect 35180 35332 35236 35388
rect 35236 35332 35240 35388
rect 35176 35328 35240 35332
rect 19576 34844 19640 34848
rect 19576 34788 19580 34844
rect 19580 34788 19636 34844
rect 19636 34788 19640 34844
rect 19576 34784 19640 34788
rect 19656 34844 19720 34848
rect 19656 34788 19660 34844
rect 19660 34788 19716 34844
rect 19716 34788 19720 34844
rect 19656 34784 19720 34788
rect 19736 34844 19800 34848
rect 19736 34788 19740 34844
rect 19740 34788 19796 34844
rect 19796 34788 19800 34844
rect 19736 34784 19800 34788
rect 19816 34844 19880 34848
rect 19816 34788 19820 34844
rect 19820 34788 19876 34844
rect 19876 34788 19880 34844
rect 19816 34784 19880 34788
rect 50296 34844 50360 34848
rect 50296 34788 50300 34844
rect 50300 34788 50356 34844
rect 50356 34788 50360 34844
rect 50296 34784 50360 34788
rect 50376 34844 50440 34848
rect 50376 34788 50380 34844
rect 50380 34788 50436 34844
rect 50436 34788 50440 34844
rect 50376 34784 50440 34788
rect 50456 34844 50520 34848
rect 50456 34788 50460 34844
rect 50460 34788 50516 34844
rect 50516 34788 50520 34844
rect 50456 34784 50520 34788
rect 50536 34844 50600 34848
rect 50536 34788 50540 34844
rect 50540 34788 50596 34844
rect 50596 34788 50600 34844
rect 50536 34784 50600 34788
rect 4216 34300 4280 34304
rect 4216 34244 4220 34300
rect 4220 34244 4276 34300
rect 4276 34244 4280 34300
rect 4216 34240 4280 34244
rect 4296 34300 4360 34304
rect 4296 34244 4300 34300
rect 4300 34244 4356 34300
rect 4356 34244 4360 34300
rect 4296 34240 4360 34244
rect 4376 34300 4440 34304
rect 4376 34244 4380 34300
rect 4380 34244 4436 34300
rect 4436 34244 4440 34300
rect 4376 34240 4440 34244
rect 4456 34300 4520 34304
rect 4456 34244 4460 34300
rect 4460 34244 4516 34300
rect 4516 34244 4520 34300
rect 4456 34240 4520 34244
rect 34936 34300 35000 34304
rect 34936 34244 34940 34300
rect 34940 34244 34996 34300
rect 34996 34244 35000 34300
rect 34936 34240 35000 34244
rect 35016 34300 35080 34304
rect 35016 34244 35020 34300
rect 35020 34244 35076 34300
rect 35076 34244 35080 34300
rect 35016 34240 35080 34244
rect 35096 34300 35160 34304
rect 35096 34244 35100 34300
rect 35100 34244 35156 34300
rect 35156 34244 35160 34300
rect 35096 34240 35160 34244
rect 35176 34300 35240 34304
rect 35176 34244 35180 34300
rect 35180 34244 35236 34300
rect 35236 34244 35240 34300
rect 35176 34240 35240 34244
rect 19576 33756 19640 33760
rect 19576 33700 19580 33756
rect 19580 33700 19636 33756
rect 19636 33700 19640 33756
rect 19576 33696 19640 33700
rect 19656 33756 19720 33760
rect 19656 33700 19660 33756
rect 19660 33700 19716 33756
rect 19716 33700 19720 33756
rect 19656 33696 19720 33700
rect 19736 33756 19800 33760
rect 19736 33700 19740 33756
rect 19740 33700 19796 33756
rect 19796 33700 19800 33756
rect 19736 33696 19800 33700
rect 19816 33756 19880 33760
rect 19816 33700 19820 33756
rect 19820 33700 19876 33756
rect 19876 33700 19880 33756
rect 19816 33696 19880 33700
rect 50296 33756 50360 33760
rect 50296 33700 50300 33756
rect 50300 33700 50356 33756
rect 50356 33700 50360 33756
rect 50296 33696 50360 33700
rect 50376 33756 50440 33760
rect 50376 33700 50380 33756
rect 50380 33700 50436 33756
rect 50436 33700 50440 33756
rect 50376 33696 50440 33700
rect 50456 33756 50520 33760
rect 50456 33700 50460 33756
rect 50460 33700 50516 33756
rect 50516 33700 50520 33756
rect 50456 33696 50520 33700
rect 50536 33756 50600 33760
rect 50536 33700 50540 33756
rect 50540 33700 50596 33756
rect 50596 33700 50600 33756
rect 50536 33696 50600 33700
rect 4216 33212 4280 33216
rect 4216 33156 4220 33212
rect 4220 33156 4276 33212
rect 4276 33156 4280 33212
rect 4216 33152 4280 33156
rect 4296 33212 4360 33216
rect 4296 33156 4300 33212
rect 4300 33156 4356 33212
rect 4356 33156 4360 33212
rect 4296 33152 4360 33156
rect 4376 33212 4440 33216
rect 4376 33156 4380 33212
rect 4380 33156 4436 33212
rect 4436 33156 4440 33212
rect 4376 33152 4440 33156
rect 4456 33212 4520 33216
rect 4456 33156 4460 33212
rect 4460 33156 4516 33212
rect 4516 33156 4520 33212
rect 4456 33152 4520 33156
rect 34936 33212 35000 33216
rect 34936 33156 34940 33212
rect 34940 33156 34996 33212
rect 34996 33156 35000 33212
rect 34936 33152 35000 33156
rect 35016 33212 35080 33216
rect 35016 33156 35020 33212
rect 35020 33156 35076 33212
rect 35076 33156 35080 33212
rect 35016 33152 35080 33156
rect 35096 33212 35160 33216
rect 35096 33156 35100 33212
rect 35100 33156 35156 33212
rect 35156 33156 35160 33212
rect 35096 33152 35160 33156
rect 35176 33212 35240 33216
rect 35176 33156 35180 33212
rect 35180 33156 35236 33212
rect 35236 33156 35240 33212
rect 35176 33152 35240 33156
rect 19576 32668 19640 32672
rect 19576 32612 19580 32668
rect 19580 32612 19636 32668
rect 19636 32612 19640 32668
rect 19576 32608 19640 32612
rect 19656 32668 19720 32672
rect 19656 32612 19660 32668
rect 19660 32612 19716 32668
rect 19716 32612 19720 32668
rect 19656 32608 19720 32612
rect 19736 32668 19800 32672
rect 19736 32612 19740 32668
rect 19740 32612 19796 32668
rect 19796 32612 19800 32668
rect 19736 32608 19800 32612
rect 19816 32668 19880 32672
rect 19816 32612 19820 32668
rect 19820 32612 19876 32668
rect 19876 32612 19880 32668
rect 19816 32608 19880 32612
rect 50296 32668 50360 32672
rect 50296 32612 50300 32668
rect 50300 32612 50356 32668
rect 50356 32612 50360 32668
rect 50296 32608 50360 32612
rect 50376 32668 50440 32672
rect 50376 32612 50380 32668
rect 50380 32612 50436 32668
rect 50436 32612 50440 32668
rect 50376 32608 50440 32612
rect 50456 32668 50520 32672
rect 50456 32612 50460 32668
rect 50460 32612 50516 32668
rect 50516 32612 50520 32668
rect 50456 32608 50520 32612
rect 50536 32668 50600 32672
rect 50536 32612 50540 32668
rect 50540 32612 50596 32668
rect 50596 32612 50600 32668
rect 50536 32608 50600 32612
rect 4216 32124 4280 32128
rect 4216 32068 4220 32124
rect 4220 32068 4276 32124
rect 4276 32068 4280 32124
rect 4216 32064 4280 32068
rect 4296 32124 4360 32128
rect 4296 32068 4300 32124
rect 4300 32068 4356 32124
rect 4356 32068 4360 32124
rect 4296 32064 4360 32068
rect 4376 32124 4440 32128
rect 4376 32068 4380 32124
rect 4380 32068 4436 32124
rect 4436 32068 4440 32124
rect 4376 32064 4440 32068
rect 4456 32124 4520 32128
rect 4456 32068 4460 32124
rect 4460 32068 4516 32124
rect 4516 32068 4520 32124
rect 4456 32064 4520 32068
rect 34936 32124 35000 32128
rect 34936 32068 34940 32124
rect 34940 32068 34996 32124
rect 34996 32068 35000 32124
rect 34936 32064 35000 32068
rect 35016 32124 35080 32128
rect 35016 32068 35020 32124
rect 35020 32068 35076 32124
rect 35076 32068 35080 32124
rect 35016 32064 35080 32068
rect 35096 32124 35160 32128
rect 35096 32068 35100 32124
rect 35100 32068 35156 32124
rect 35156 32068 35160 32124
rect 35096 32064 35160 32068
rect 35176 32124 35240 32128
rect 35176 32068 35180 32124
rect 35180 32068 35236 32124
rect 35236 32068 35240 32124
rect 35176 32064 35240 32068
rect 19576 31580 19640 31584
rect 19576 31524 19580 31580
rect 19580 31524 19636 31580
rect 19636 31524 19640 31580
rect 19576 31520 19640 31524
rect 19656 31580 19720 31584
rect 19656 31524 19660 31580
rect 19660 31524 19716 31580
rect 19716 31524 19720 31580
rect 19656 31520 19720 31524
rect 19736 31580 19800 31584
rect 19736 31524 19740 31580
rect 19740 31524 19796 31580
rect 19796 31524 19800 31580
rect 19736 31520 19800 31524
rect 19816 31580 19880 31584
rect 19816 31524 19820 31580
rect 19820 31524 19876 31580
rect 19876 31524 19880 31580
rect 19816 31520 19880 31524
rect 50296 31580 50360 31584
rect 50296 31524 50300 31580
rect 50300 31524 50356 31580
rect 50356 31524 50360 31580
rect 50296 31520 50360 31524
rect 50376 31580 50440 31584
rect 50376 31524 50380 31580
rect 50380 31524 50436 31580
rect 50436 31524 50440 31580
rect 50376 31520 50440 31524
rect 50456 31580 50520 31584
rect 50456 31524 50460 31580
rect 50460 31524 50516 31580
rect 50516 31524 50520 31580
rect 50456 31520 50520 31524
rect 50536 31580 50600 31584
rect 50536 31524 50540 31580
rect 50540 31524 50596 31580
rect 50596 31524 50600 31580
rect 50536 31520 50600 31524
rect 4216 31036 4280 31040
rect 4216 30980 4220 31036
rect 4220 30980 4276 31036
rect 4276 30980 4280 31036
rect 4216 30976 4280 30980
rect 4296 31036 4360 31040
rect 4296 30980 4300 31036
rect 4300 30980 4356 31036
rect 4356 30980 4360 31036
rect 4296 30976 4360 30980
rect 4376 31036 4440 31040
rect 4376 30980 4380 31036
rect 4380 30980 4436 31036
rect 4436 30980 4440 31036
rect 4376 30976 4440 30980
rect 4456 31036 4520 31040
rect 4456 30980 4460 31036
rect 4460 30980 4516 31036
rect 4516 30980 4520 31036
rect 4456 30976 4520 30980
rect 34936 31036 35000 31040
rect 34936 30980 34940 31036
rect 34940 30980 34996 31036
rect 34996 30980 35000 31036
rect 34936 30976 35000 30980
rect 35016 31036 35080 31040
rect 35016 30980 35020 31036
rect 35020 30980 35076 31036
rect 35076 30980 35080 31036
rect 35016 30976 35080 30980
rect 35096 31036 35160 31040
rect 35096 30980 35100 31036
rect 35100 30980 35156 31036
rect 35156 30980 35160 31036
rect 35096 30976 35160 30980
rect 35176 31036 35240 31040
rect 35176 30980 35180 31036
rect 35180 30980 35236 31036
rect 35236 30980 35240 31036
rect 35176 30976 35240 30980
rect 19576 30492 19640 30496
rect 19576 30436 19580 30492
rect 19580 30436 19636 30492
rect 19636 30436 19640 30492
rect 19576 30432 19640 30436
rect 19656 30492 19720 30496
rect 19656 30436 19660 30492
rect 19660 30436 19716 30492
rect 19716 30436 19720 30492
rect 19656 30432 19720 30436
rect 19736 30492 19800 30496
rect 19736 30436 19740 30492
rect 19740 30436 19796 30492
rect 19796 30436 19800 30492
rect 19736 30432 19800 30436
rect 19816 30492 19880 30496
rect 19816 30436 19820 30492
rect 19820 30436 19876 30492
rect 19876 30436 19880 30492
rect 19816 30432 19880 30436
rect 50296 30492 50360 30496
rect 50296 30436 50300 30492
rect 50300 30436 50356 30492
rect 50356 30436 50360 30492
rect 50296 30432 50360 30436
rect 50376 30492 50440 30496
rect 50376 30436 50380 30492
rect 50380 30436 50436 30492
rect 50436 30436 50440 30492
rect 50376 30432 50440 30436
rect 50456 30492 50520 30496
rect 50456 30436 50460 30492
rect 50460 30436 50516 30492
rect 50516 30436 50520 30492
rect 50456 30432 50520 30436
rect 50536 30492 50600 30496
rect 50536 30436 50540 30492
rect 50540 30436 50596 30492
rect 50596 30436 50600 30492
rect 50536 30432 50600 30436
rect 4216 29948 4280 29952
rect 4216 29892 4220 29948
rect 4220 29892 4276 29948
rect 4276 29892 4280 29948
rect 4216 29888 4280 29892
rect 4296 29948 4360 29952
rect 4296 29892 4300 29948
rect 4300 29892 4356 29948
rect 4356 29892 4360 29948
rect 4296 29888 4360 29892
rect 4376 29948 4440 29952
rect 4376 29892 4380 29948
rect 4380 29892 4436 29948
rect 4436 29892 4440 29948
rect 4376 29888 4440 29892
rect 4456 29948 4520 29952
rect 4456 29892 4460 29948
rect 4460 29892 4516 29948
rect 4516 29892 4520 29948
rect 4456 29888 4520 29892
rect 34936 29948 35000 29952
rect 34936 29892 34940 29948
rect 34940 29892 34996 29948
rect 34996 29892 35000 29948
rect 34936 29888 35000 29892
rect 35016 29948 35080 29952
rect 35016 29892 35020 29948
rect 35020 29892 35076 29948
rect 35076 29892 35080 29948
rect 35016 29888 35080 29892
rect 35096 29948 35160 29952
rect 35096 29892 35100 29948
rect 35100 29892 35156 29948
rect 35156 29892 35160 29948
rect 35096 29888 35160 29892
rect 35176 29948 35240 29952
rect 35176 29892 35180 29948
rect 35180 29892 35236 29948
rect 35236 29892 35240 29948
rect 35176 29888 35240 29892
rect 19576 29404 19640 29408
rect 19576 29348 19580 29404
rect 19580 29348 19636 29404
rect 19636 29348 19640 29404
rect 19576 29344 19640 29348
rect 19656 29404 19720 29408
rect 19656 29348 19660 29404
rect 19660 29348 19716 29404
rect 19716 29348 19720 29404
rect 19656 29344 19720 29348
rect 19736 29404 19800 29408
rect 19736 29348 19740 29404
rect 19740 29348 19796 29404
rect 19796 29348 19800 29404
rect 19736 29344 19800 29348
rect 19816 29404 19880 29408
rect 19816 29348 19820 29404
rect 19820 29348 19876 29404
rect 19876 29348 19880 29404
rect 19816 29344 19880 29348
rect 50296 29404 50360 29408
rect 50296 29348 50300 29404
rect 50300 29348 50356 29404
rect 50356 29348 50360 29404
rect 50296 29344 50360 29348
rect 50376 29404 50440 29408
rect 50376 29348 50380 29404
rect 50380 29348 50436 29404
rect 50436 29348 50440 29404
rect 50376 29344 50440 29348
rect 50456 29404 50520 29408
rect 50456 29348 50460 29404
rect 50460 29348 50516 29404
rect 50516 29348 50520 29404
rect 50456 29344 50520 29348
rect 50536 29404 50600 29408
rect 50536 29348 50540 29404
rect 50540 29348 50596 29404
rect 50596 29348 50600 29404
rect 50536 29344 50600 29348
rect 4216 28860 4280 28864
rect 4216 28804 4220 28860
rect 4220 28804 4276 28860
rect 4276 28804 4280 28860
rect 4216 28800 4280 28804
rect 4296 28860 4360 28864
rect 4296 28804 4300 28860
rect 4300 28804 4356 28860
rect 4356 28804 4360 28860
rect 4296 28800 4360 28804
rect 4376 28860 4440 28864
rect 4376 28804 4380 28860
rect 4380 28804 4436 28860
rect 4436 28804 4440 28860
rect 4376 28800 4440 28804
rect 4456 28860 4520 28864
rect 4456 28804 4460 28860
rect 4460 28804 4516 28860
rect 4516 28804 4520 28860
rect 4456 28800 4520 28804
rect 34936 28860 35000 28864
rect 34936 28804 34940 28860
rect 34940 28804 34996 28860
rect 34996 28804 35000 28860
rect 34936 28800 35000 28804
rect 35016 28860 35080 28864
rect 35016 28804 35020 28860
rect 35020 28804 35076 28860
rect 35076 28804 35080 28860
rect 35016 28800 35080 28804
rect 35096 28860 35160 28864
rect 35096 28804 35100 28860
rect 35100 28804 35156 28860
rect 35156 28804 35160 28860
rect 35096 28800 35160 28804
rect 35176 28860 35240 28864
rect 35176 28804 35180 28860
rect 35180 28804 35236 28860
rect 35236 28804 35240 28860
rect 35176 28800 35240 28804
rect 19576 28316 19640 28320
rect 19576 28260 19580 28316
rect 19580 28260 19636 28316
rect 19636 28260 19640 28316
rect 19576 28256 19640 28260
rect 19656 28316 19720 28320
rect 19656 28260 19660 28316
rect 19660 28260 19716 28316
rect 19716 28260 19720 28316
rect 19656 28256 19720 28260
rect 19736 28316 19800 28320
rect 19736 28260 19740 28316
rect 19740 28260 19796 28316
rect 19796 28260 19800 28316
rect 19736 28256 19800 28260
rect 19816 28316 19880 28320
rect 19816 28260 19820 28316
rect 19820 28260 19876 28316
rect 19876 28260 19880 28316
rect 19816 28256 19880 28260
rect 50296 28316 50360 28320
rect 50296 28260 50300 28316
rect 50300 28260 50356 28316
rect 50356 28260 50360 28316
rect 50296 28256 50360 28260
rect 50376 28316 50440 28320
rect 50376 28260 50380 28316
rect 50380 28260 50436 28316
rect 50436 28260 50440 28316
rect 50376 28256 50440 28260
rect 50456 28316 50520 28320
rect 50456 28260 50460 28316
rect 50460 28260 50516 28316
rect 50516 28260 50520 28316
rect 50456 28256 50520 28260
rect 50536 28316 50600 28320
rect 50536 28260 50540 28316
rect 50540 28260 50596 28316
rect 50596 28260 50600 28316
rect 50536 28256 50600 28260
rect 4216 27772 4280 27776
rect 4216 27716 4220 27772
rect 4220 27716 4276 27772
rect 4276 27716 4280 27772
rect 4216 27712 4280 27716
rect 4296 27772 4360 27776
rect 4296 27716 4300 27772
rect 4300 27716 4356 27772
rect 4356 27716 4360 27772
rect 4296 27712 4360 27716
rect 4376 27772 4440 27776
rect 4376 27716 4380 27772
rect 4380 27716 4436 27772
rect 4436 27716 4440 27772
rect 4376 27712 4440 27716
rect 4456 27772 4520 27776
rect 4456 27716 4460 27772
rect 4460 27716 4516 27772
rect 4516 27716 4520 27772
rect 4456 27712 4520 27716
rect 34936 27772 35000 27776
rect 34936 27716 34940 27772
rect 34940 27716 34996 27772
rect 34996 27716 35000 27772
rect 34936 27712 35000 27716
rect 35016 27772 35080 27776
rect 35016 27716 35020 27772
rect 35020 27716 35076 27772
rect 35076 27716 35080 27772
rect 35016 27712 35080 27716
rect 35096 27772 35160 27776
rect 35096 27716 35100 27772
rect 35100 27716 35156 27772
rect 35156 27716 35160 27772
rect 35096 27712 35160 27716
rect 35176 27772 35240 27776
rect 35176 27716 35180 27772
rect 35180 27716 35236 27772
rect 35236 27716 35240 27772
rect 35176 27712 35240 27716
rect 19576 27228 19640 27232
rect 19576 27172 19580 27228
rect 19580 27172 19636 27228
rect 19636 27172 19640 27228
rect 19576 27168 19640 27172
rect 19656 27228 19720 27232
rect 19656 27172 19660 27228
rect 19660 27172 19716 27228
rect 19716 27172 19720 27228
rect 19656 27168 19720 27172
rect 19736 27228 19800 27232
rect 19736 27172 19740 27228
rect 19740 27172 19796 27228
rect 19796 27172 19800 27228
rect 19736 27168 19800 27172
rect 19816 27228 19880 27232
rect 19816 27172 19820 27228
rect 19820 27172 19876 27228
rect 19876 27172 19880 27228
rect 19816 27168 19880 27172
rect 50296 27228 50360 27232
rect 50296 27172 50300 27228
rect 50300 27172 50356 27228
rect 50356 27172 50360 27228
rect 50296 27168 50360 27172
rect 50376 27228 50440 27232
rect 50376 27172 50380 27228
rect 50380 27172 50436 27228
rect 50436 27172 50440 27228
rect 50376 27168 50440 27172
rect 50456 27228 50520 27232
rect 50456 27172 50460 27228
rect 50460 27172 50516 27228
rect 50516 27172 50520 27228
rect 50456 27168 50520 27172
rect 50536 27228 50600 27232
rect 50536 27172 50540 27228
rect 50540 27172 50596 27228
rect 50596 27172 50600 27228
rect 50536 27168 50600 27172
rect 4216 26684 4280 26688
rect 4216 26628 4220 26684
rect 4220 26628 4276 26684
rect 4276 26628 4280 26684
rect 4216 26624 4280 26628
rect 4296 26684 4360 26688
rect 4296 26628 4300 26684
rect 4300 26628 4356 26684
rect 4356 26628 4360 26684
rect 4296 26624 4360 26628
rect 4376 26684 4440 26688
rect 4376 26628 4380 26684
rect 4380 26628 4436 26684
rect 4436 26628 4440 26684
rect 4376 26624 4440 26628
rect 4456 26684 4520 26688
rect 4456 26628 4460 26684
rect 4460 26628 4516 26684
rect 4516 26628 4520 26684
rect 4456 26624 4520 26628
rect 34936 26684 35000 26688
rect 34936 26628 34940 26684
rect 34940 26628 34996 26684
rect 34996 26628 35000 26684
rect 34936 26624 35000 26628
rect 35016 26684 35080 26688
rect 35016 26628 35020 26684
rect 35020 26628 35076 26684
rect 35076 26628 35080 26684
rect 35016 26624 35080 26628
rect 35096 26684 35160 26688
rect 35096 26628 35100 26684
rect 35100 26628 35156 26684
rect 35156 26628 35160 26684
rect 35096 26624 35160 26628
rect 35176 26684 35240 26688
rect 35176 26628 35180 26684
rect 35180 26628 35236 26684
rect 35236 26628 35240 26684
rect 35176 26624 35240 26628
rect 21220 26556 21284 26620
rect 19576 26140 19640 26144
rect 19576 26084 19580 26140
rect 19580 26084 19636 26140
rect 19636 26084 19640 26140
rect 19576 26080 19640 26084
rect 19656 26140 19720 26144
rect 19656 26084 19660 26140
rect 19660 26084 19716 26140
rect 19716 26084 19720 26140
rect 19656 26080 19720 26084
rect 19736 26140 19800 26144
rect 19736 26084 19740 26140
rect 19740 26084 19796 26140
rect 19796 26084 19800 26140
rect 19736 26080 19800 26084
rect 19816 26140 19880 26144
rect 19816 26084 19820 26140
rect 19820 26084 19876 26140
rect 19876 26084 19880 26140
rect 19816 26080 19880 26084
rect 50296 26140 50360 26144
rect 50296 26084 50300 26140
rect 50300 26084 50356 26140
rect 50356 26084 50360 26140
rect 50296 26080 50360 26084
rect 50376 26140 50440 26144
rect 50376 26084 50380 26140
rect 50380 26084 50436 26140
rect 50436 26084 50440 26140
rect 50376 26080 50440 26084
rect 50456 26140 50520 26144
rect 50456 26084 50460 26140
rect 50460 26084 50516 26140
rect 50516 26084 50520 26140
rect 50456 26080 50520 26084
rect 50536 26140 50600 26144
rect 50536 26084 50540 26140
rect 50540 26084 50596 26140
rect 50596 26084 50600 26140
rect 50536 26080 50600 26084
rect 23612 25876 23676 25940
rect 4216 25596 4280 25600
rect 4216 25540 4220 25596
rect 4220 25540 4276 25596
rect 4276 25540 4280 25596
rect 4216 25536 4280 25540
rect 4296 25596 4360 25600
rect 4296 25540 4300 25596
rect 4300 25540 4356 25596
rect 4356 25540 4360 25596
rect 4296 25536 4360 25540
rect 4376 25596 4440 25600
rect 4376 25540 4380 25596
rect 4380 25540 4436 25596
rect 4436 25540 4440 25596
rect 4376 25536 4440 25540
rect 4456 25596 4520 25600
rect 4456 25540 4460 25596
rect 4460 25540 4516 25596
rect 4516 25540 4520 25596
rect 4456 25536 4520 25540
rect 34936 25596 35000 25600
rect 34936 25540 34940 25596
rect 34940 25540 34996 25596
rect 34996 25540 35000 25596
rect 34936 25536 35000 25540
rect 35016 25596 35080 25600
rect 35016 25540 35020 25596
rect 35020 25540 35076 25596
rect 35076 25540 35080 25596
rect 35016 25536 35080 25540
rect 35096 25596 35160 25600
rect 35096 25540 35100 25596
rect 35100 25540 35156 25596
rect 35156 25540 35160 25596
rect 35096 25536 35160 25540
rect 35176 25596 35240 25600
rect 35176 25540 35180 25596
rect 35180 25540 35236 25596
rect 35236 25540 35240 25596
rect 35176 25536 35240 25540
rect 19576 25052 19640 25056
rect 19576 24996 19580 25052
rect 19580 24996 19636 25052
rect 19636 24996 19640 25052
rect 19576 24992 19640 24996
rect 19656 25052 19720 25056
rect 19656 24996 19660 25052
rect 19660 24996 19716 25052
rect 19716 24996 19720 25052
rect 19656 24992 19720 24996
rect 19736 25052 19800 25056
rect 19736 24996 19740 25052
rect 19740 24996 19796 25052
rect 19796 24996 19800 25052
rect 19736 24992 19800 24996
rect 19816 25052 19880 25056
rect 19816 24996 19820 25052
rect 19820 24996 19876 25052
rect 19876 24996 19880 25052
rect 19816 24992 19880 24996
rect 50296 25052 50360 25056
rect 50296 24996 50300 25052
rect 50300 24996 50356 25052
rect 50356 24996 50360 25052
rect 50296 24992 50360 24996
rect 50376 25052 50440 25056
rect 50376 24996 50380 25052
rect 50380 24996 50436 25052
rect 50436 24996 50440 25052
rect 50376 24992 50440 24996
rect 50456 25052 50520 25056
rect 50456 24996 50460 25052
rect 50460 24996 50516 25052
rect 50516 24996 50520 25052
rect 50456 24992 50520 24996
rect 50536 25052 50600 25056
rect 50536 24996 50540 25052
rect 50540 24996 50596 25052
rect 50596 24996 50600 25052
rect 50536 24992 50600 24996
rect 4216 24508 4280 24512
rect 4216 24452 4220 24508
rect 4220 24452 4276 24508
rect 4276 24452 4280 24508
rect 4216 24448 4280 24452
rect 4296 24508 4360 24512
rect 4296 24452 4300 24508
rect 4300 24452 4356 24508
rect 4356 24452 4360 24508
rect 4296 24448 4360 24452
rect 4376 24508 4440 24512
rect 4376 24452 4380 24508
rect 4380 24452 4436 24508
rect 4436 24452 4440 24508
rect 4376 24448 4440 24452
rect 4456 24508 4520 24512
rect 4456 24452 4460 24508
rect 4460 24452 4516 24508
rect 4516 24452 4520 24508
rect 4456 24448 4520 24452
rect 34936 24508 35000 24512
rect 34936 24452 34940 24508
rect 34940 24452 34996 24508
rect 34996 24452 35000 24508
rect 34936 24448 35000 24452
rect 35016 24508 35080 24512
rect 35016 24452 35020 24508
rect 35020 24452 35076 24508
rect 35076 24452 35080 24508
rect 35016 24448 35080 24452
rect 35096 24508 35160 24512
rect 35096 24452 35100 24508
rect 35100 24452 35156 24508
rect 35156 24452 35160 24508
rect 35096 24448 35160 24452
rect 35176 24508 35240 24512
rect 35176 24452 35180 24508
rect 35180 24452 35236 24508
rect 35236 24452 35240 24508
rect 35176 24448 35240 24452
rect 19576 23964 19640 23968
rect 19576 23908 19580 23964
rect 19580 23908 19636 23964
rect 19636 23908 19640 23964
rect 19576 23904 19640 23908
rect 19656 23964 19720 23968
rect 19656 23908 19660 23964
rect 19660 23908 19716 23964
rect 19716 23908 19720 23964
rect 19656 23904 19720 23908
rect 19736 23964 19800 23968
rect 19736 23908 19740 23964
rect 19740 23908 19796 23964
rect 19796 23908 19800 23964
rect 19736 23904 19800 23908
rect 19816 23964 19880 23968
rect 19816 23908 19820 23964
rect 19820 23908 19876 23964
rect 19876 23908 19880 23964
rect 19816 23904 19880 23908
rect 50296 23964 50360 23968
rect 50296 23908 50300 23964
rect 50300 23908 50356 23964
rect 50356 23908 50360 23964
rect 50296 23904 50360 23908
rect 50376 23964 50440 23968
rect 50376 23908 50380 23964
rect 50380 23908 50436 23964
rect 50436 23908 50440 23964
rect 50376 23904 50440 23908
rect 50456 23964 50520 23968
rect 50456 23908 50460 23964
rect 50460 23908 50516 23964
rect 50516 23908 50520 23964
rect 50456 23904 50520 23908
rect 50536 23964 50600 23968
rect 50536 23908 50540 23964
rect 50540 23908 50596 23964
rect 50596 23908 50600 23964
rect 50536 23904 50600 23908
rect 23428 23428 23492 23492
rect 4216 23420 4280 23424
rect 4216 23364 4220 23420
rect 4220 23364 4276 23420
rect 4276 23364 4280 23420
rect 4216 23360 4280 23364
rect 4296 23420 4360 23424
rect 4296 23364 4300 23420
rect 4300 23364 4356 23420
rect 4356 23364 4360 23420
rect 4296 23360 4360 23364
rect 4376 23420 4440 23424
rect 4376 23364 4380 23420
rect 4380 23364 4436 23420
rect 4436 23364 4440 23420
rect 4376 23360 4440 23364
rect 4456 23420 4520 23424
rect 4456 23364 4460 23420
rect 4460 23364 4516 23420
rect 4516 23364 4520 23420
rect 4456 23360 4520 23364
rect 34936 23420 35000 23424
rect 34936 23364 34940 23420
rect 34940 23364 34996 23420
rect 34996 23364 35000 23420
rect 34936 23360 35000 23364
rect 35016 23420 35080 23424
rect 35016 23364 35020 23420
rect 35020 23364 35076 23420
rect 35076 23364 35080 23420
rect 35016 23360 35080 23364
rect 35096 23420 35160 23424
rect 35096 23364 35100 23420
rect 35100 23364 35156 23420
rect 35156 23364 35160 23420
rect 35096 23360 35160 23364
rect 35176 23420 35240 23424
rect 35176 23364 35180 23420
rect 35180 23364 35236 23420
rect 35236 23364 35240 23420
rect 35176 23360 35240 23364
rect 19576 22876 19640 22880
rect 19576 22820 19580 22876
rect 19580 22820 19636 22876
rect 19636 22820 19640 22876
rect 19576 22816 19640 22820
rect 19656 22876 19720 22880
rect 19656 22820 19660 22876
rect 19660 22820 19716 22876
rect 19716 22820 19720 22876
rect 19656 22816 19720 22820
rect 19736 22876 19800 22880
rect 19736 22820 19740 22876
rect 19740 22820 19796 22876
rect 19796 22820 19800 22876
rect 19736 22816 19800 22820
rect 19816 22876 19880 22880
rect 19816 22820 19820 22876
rect 19820 22820 19876 22876
rect 19876 22820 19880 22876
rect 19816 22816 19880 22820
rect 50296 22876 50360 22880
rect 50296 22820 50300 22876
rect 50300 22820 50356 22876
rect 50356 22820 50360 22876
rect 50296 22816 50360 22820
rect 50376 22876 50440 22880
rect 50376 22820 50380 22876
rect 50380 22820 50436 22876
rect 50436 22820 50440 22876
rect 50376 22816 50440 22820
rect 50456 22876 50520 22880
rect 50456 22820 50460 22876
rect 50460 22820 50516 22876
rect 50516 22820 50520 22876
rect 50456 22816 50520 22820
rect 50536 22876 50600 22880
rect 50536 22820 50540 22876
rect 50540 22820 50596 22876
rect 50596 22820 50600 22876
rect 50536 22816 50600 22820
rect 4216 22332 4280 22336
rect 4216 22276 4220 22332
rect 4220 22276 4276 22332
rect 4276 22276 4280 22332
rect 4216 22272 4280 22276
rect 4296 22332 4360 22336
rect 4296 22276 4300 22332
rect 4300 22276 4356 22332
rect 4356 22276 4360 22332
rect 4296 22272 4360 22276
rect 4376 22332 4440 22336
rect 4376 22276 4380 22332
rect 4380 22276 4436 22332
rect 4436 22276 4440 22332
rect 4376 22272 4440 22276
rect 4456 22332 4520 22336
rect 4456 22276 4460 22332
rect 4460 22276 4516 22332
rect 4516 22276 4520 22332
rect 4456 22272 4520 22276
rect 34936 22332 35000 22336
rect 34936 22276 34940 22332
rect 34940 22276 34996 22332
rect 34996 22276 35000 22332
rect 34936 22272 35000 22276
rect 35016 22332 35080 22336
rect 35016 22276 35020 22332
rect 35020 22276 35076 22332
rect 35076 22276 35080 22332
rect 35016 22272 35080 22276
rect 35096 22332 35160 22336
rect 35096 22276 35100 22332
rect 35100 22276 35156 22332
rect 35156 22276 35160 22332
rect 35096 22272 35160 22276
rect 35176 22332 35240 22336
rect 35176 22276 35180 22332
rect 35180 22276 35236 22332
rect 35236 22276 35240 22332
rect 35176 22272 35240 22276
rect 19576 21788 19640 21792
rect 19576 21732 19580 21788
rect 19580 21732 19636 21788
rect 19636 21732 19640 21788
rect 19576 21728 19640 21732
rect 19656 21788 19720 21792
rect 19656 21732 19660 21788
rect 19660 21732 19716 21788
rect 19716 21732 19720 21788
rect 19656 21728 19720 21732
rect 19736 21788 19800 21792
rect 19736 21732 19740 21788
rect 19740 21732 19796 21788
rect 19796 21732 19800 21788
rect 19736 21728 19800 21732
rect 19816 21788 19880 21792
rect 19816 21732 19820 21788
rect 19820 21732 19876 21788
rect 19876 21732 19880 21788
rect 19816 21728 19880 21732
rect 50296 21788 50360 21792
rect 50296 21732 50300 21788
rect 50300 21732 50356 21788
rect 50356 21732 50360 21788
rect 50296 21728 50360 21732
rect 50376 21788 50440 21792
rect 50376 21732 50380 21788
rect 50380 21732 50436 21788
rect 50436 21732 50440 21788
rect 50376 21728 50440 21732
rect 50456 21788 50520 21792
rect 50456 21732 50460 21788
rect 50460 21732 50516 21788
rect 50516 21732 50520 21788
rect 50456 21728 50520 21732
rect 50536 21788 50600 21792
rect 50536 21732 50540 21788
rect 50540 21732 50596 21788
rect 50596 21732 50600 21788
rect 50536 21728 50600 21732
rect 4216 21244 4280 21248
rect 4216 21188 4220 21244
rect 4220 21188 4276 21244
rect 4276 21188 4280 21244
rect 4216 21184 4280 21188
rect 4296 21244 4360 21248
rect 4296 21188 4300 21244
rect 4300 21188 4356 21244
rect 4356 21188 4360 21244
rect 4296 21184 4360 21188
rect 4376 21244 4440 21248
rect 4376 21188 4380 21244
rect 4380 21188 4436 21244
rect 4436 21188 4440 21244
rect 4376 21184 4440 21188
rect 4456 21244 4520 21248
rect 4456 21188 4460 21244
rect 4460 21188 4516 21244
rect 4516 21188 4520 21244
rect 4456 21184 4520 21188
rect 34936 21244 35000 21248
rect 34936 21188 34940 21244
rect 34940 21188 34996 21244
rect 34996 21188 35000 21244
rect 34936 21184 35000 21188
rect 35016 21244 35080 21248
rect 35016 21188 35020 21244
rect 35020 21188 35076 21244
rect 35076 21188 35080 21244
rect 35016 21184 35080 21188
rect 35096 21244 35160 21248
rect 35096 21188 35100 21244
rect 35100 21188 35156 21244
rect 35156 21188 35160 21244
rect 35096 21184 35160 21188
rect 35176 21244 35240 21248
rect 35176 21188 35180 21244
rect 35180 21188 35236 21244
rect 35236 21188 35240 21244
rect 35176 21184 35240 21188
rect 19576 20700 19640 20704
rect 19576 20644 19580 20700
rect 19580 20644 19636 20700
rect 19636 20644 19640 20700
rect 19576 20640 19640 20644
rect 19656 20700 19720 20704
rect 19656 20644 19660 20700
rect 19660 20644 19716 20700
rect 19716 20644 19720 20700
rect 19656 20640 19720 20644
rect 19736 20700 19800 20704
rect 19736 20644 19740 20700
rect 19740 20644 19796 20700
rect 19796 20644 19800 20700
rect 19736 20640 19800 20644
rect 19816 20700 19880 20704
rect 19816 20644 19820 20700
rect 19820 20644 19876 20700
rect 19876 20644 19880 20700
rect 19816 20640 19880 20644
rect 50296 20700 50360 20704
rect 50296 20644 50300 20700
rect 50300 20644 50356 20700
rect 50356 20644 50360 20700
rect 50296 20640 50360 20644
rect 50376 20700 50440 20704
rect 50376 20644 50380 20700
rect 50380 20644 50436 20700
rect 50436 20644 50440 20700
rect 50376 20640 50440 20644
rect 50456 20700 50520 20704
rect 50456 20644 50460 20700
rect 50460 20644 50516 20700
rect 50516 20644 50520 20700
rect 50456 20640 50520 20644
rect 50536 20700 50600 20704
rect 50536 20644 50540 20700
rect 50540 20644 50596 20700
rect 50596 20644 50600 20700
rect 50536 20640 50600 20644
rect 4216 20156 4280 20160
rect 4216 20100 4220 20156
rect 4220 20100 4276 20156
rect 4276 20100 4280 20156
rect 4216 20096 4280 20100
rect 4296 20156 4360 20160
rect 4296 20100 4300 20156
rect 4300 20100 4356 20156
rect 4356 20100 4360 20156
rect 4296 20096 4360 20100
rect 4376 20156 4440 20160
rect 4376 20100 4380 20156
rect 4380 20100 4436 20156
rect 4436 20100 4440 20156
rect 4376 20096 4440 20100
rect 4456 20156 4520 20160
rect 4456 20100 4460 20156
rect 4460 20100 4516 20156
rect 4516 20100 4520 20156
rect 4456 20096 4520 20100
rect 34936 20156 35000 20160
rect 34936 20100 34940 20156
rect 34940 20100 34996 20156
rect 34996 20100 35000 20156
rect 34936 20096 35000 20100
rect 35016 20156 35080 20160
rect 35016 20100 35020 20156
rect 35020 20100 35076 20156
rect 35076 20100 35080 20156
rect 35016 20096 35080 20100
rect 35096 20156 35160 20160
rect 35096 20100 35100 20156
rect 35100 20100 35156 20156
rect 35156 20100 35160 20156
rect 35096 20096 35160 20100
rect 35176 20156 35240 20160
rect 35176 20100 35180 20156
rect 35180 20100 35236 20156
rect 35236 20100 35240 20156
rect 35176 20096 35240 20100
rect 19576 19612 19640 19616
rect 19576 19556 19580 19612
rect 19580 19556 19636 19612
rect 19636 19556 19640 19612
rect 19576 19552 19640 19556
rect 19656 19612 19720 19616
rect 19656 19556 19660 19612
rect 19660 19556 19716 19612
rect 19716 19556 19720 19612
rect 19656 19552 19720 19556
rect 19736 19612 19800 19616
rect 19736 19556 19740 19612
rect 19740 19556 19796 19612
rect 19796 19556 19800 19612
rect 19736 19552 19800 19556
rect 19816 19612 19880 19616
rect 19816 19556 19820 19612
rect 19820 19556 19876 19612
rect 19876 19556 19880 19612
rect 19816 19552 19880 19556
rect 50296 19612 50360 19616
rect 50296 19556 50300 19612
rect 50300 19556 50356 19612
rect 50356 19556 50360 19612
rect 50296 19552 50360 19556
rect 50376 19612 50440 19616
rect 50376 19556 50380 19612
rect 50380 19556 50436 19612
rect 50436 19556 50440 19612
rect 50376 19552 50440 19556
rect 50456 19612 50520 19616
rect 50456 19556 50460 19612
rect 50460 19556 50516 19612
rect 50516 19556 50520 19612
rect 50456 19552 50520 19556
rect 50536 19612 50600 19616
rect 50536 19556 50540 19612
rect 50540 19556 50596 19612
rect 50596 19556 50600 19612
rect 50536 19552 50600 19556
rect 4216 19068 4280 19072
rect 4216 19012 4220 19068
rect 4220 19012 4276 19068
rect 4276 19012 4280 19068
rect 4216 19008 4280 19012
rect 4296 19068 4360 19072
rect 4296 19012 4300 19068
rect 4300 19012 4356 19068
rect 4356 19012 4360 19068
rect 4296 19008 4360 19012
rect 4376 19068 4440 19072
rect 4376 19012 4380 19068
rect 4380 19012 4436 19068
rect 4436 19012 4440 19068
rect 4376 19008 4440 19012
rect 4456 19068 4520 19072
rect 4456 19012 4460 19068
rect 4460 19012 4516 19068
rect 4516 19012 4520 19068
rect 4456 19008 4520 19012
rect 34936 19068 35000 19072
rect 34936 19012 34940 19068
rect 34940 19012 34996 19068
rect 34996 19012 35000 19068
rect 34936 19008 35000 19012
rect 35016 19068 35080 19072
rect 35016 19012 35020 19068
rect 35020 19012 35076 19068
rect 35076 19012 35080 19068
rect 35016 19008 35080 19012
rect 35096 19068 35160 19072
rect 35096 19012 35100 19068
rect 35100 19012 35156 19068
rect 35156 19012 35160 19068
rect 35096 19008 35160 19012
rect 35176 19068 35240 19072
rect 35176 19012 35180 19068
rect 35180 19012 35236 19068
rect 35236 19012 35240 19068
rect 35176 19008 35240 19012
rect 23612 18804 23676 18868
rect 19576 18524 19640 18528
rect 19576 18468 19580 18524
rect 19580 18468 19636 18524
rect 19636 18468 19640 18524
rect 19576 18464 19640 18468
rect 19656 18524 19720 18528
rect 19656 18468 19660 18524
rect 19660 18468 19716 18524
rect 19716 18468 19720 18524
rect 19656 18464 19720 18468
rect 19736 18524 19800 18528
rect 19736 18468 19740 18524
rect 19740 18468 19796 18524
rect 19796 18468 19800 18524
rect 19736 18464 19800 18468
rect 19816 18524 19880 18528
rect 19816 18468 19820 18524
rect 19820 18468 19876 18524
rect 19876 18468 19880 18524
rect 19816 18464 19880 18468
rect 50296 18524 50360 18528
rect 50296 18468 50300 18524
rect 50300 18468 50356 18524
rect 50356 18468 50360 18524
rect 50296 18464 50360 18468
rect 50376 18524 50440 18528
rect 50376 18468 50380 18524
rect 50380 18468 50436 18524
rect 50436 18468 50440 18524
rect 50376 18464 50440 18468
rect 50456 18524 50520 18528
rect 50456 18468 50460 18524
rect 50460 18468 50516 18524
rect 50516 18468 50520 18524
rect 50456 18464 50520 18468
rect 50536 18524 50600 18528
rect 50536 18468 50540 18524
rect 50540 18468 50596 18524
rect 50596 18468 50600 18524
rect 50536 18464 50600 18468
rect 4216 17980 4280 17984
rect 4216 17924 4220 17980
rect 4220 17924 4276 17980
rect 4276 17924 4280 17980
rect 4216 17920 4280 17924
rect 4296 17980 4360 17984
rect 4296 17924 4300 17980
rect 4300 17924 4356 17980
rect 4356 17924 4360 17980
rect 4296 17920 4360 17924
rect 4376 17980 4440 17984
rect 4376 17924 4380 17980
rect 4380 17924 4436 17980
rect 4436 17924 4440 17980
rect 4376 17920 4440 17924
rect 4456 17980 4520 17984
rect 4456 17924 4460 17980
rect 4460 17924 4516 17980
rect 4516 17924 4520 17980
rect 4456 17920 4520 17924
rect 34936 17980 35000 17984
rect 34936 17924 34940 17980
rect 34940 17924 34996 17980
rect 34996 17924 35000 17980
rect 34936 17920 35000 17924
rect 35016 17980 35080 17984
rect 35016 17924 35020 17980
rect 35020 17924 35076 17980
rect 35076 17924 35080 17980
rect 35016 17920 35080 17924
rect 35096 17980 35160 17984
rect 35096 17924 35100 17980
rect 35100 17924 35156 17980
rect 35156 17924 35160 17980
rect 35096 17920 35160 17924
rect 35176 17980 35240 17984
rect 35176 17924 35180 17980
rect 35180 17924 35236 17980
rect 35236 17924 35240 17980
rect 35176 17920 35240 17924
rect 19576 17436 19640 17440
rect 19576 17380 19580 17436
rect 19580 17380 19636 17436
rect 19636 17380 19640 17436
rect 19576 17376 19640 17380
rect 19656 17436 19720 17440
rect 19656 17380 19660 17436
rect 19660 17380 19716 17436
rect 19716 17380 19720 17436
rect 19656 17376 19720 17380
rect 19736 17436 19800 17440
rect 19736 17380 19740 17436
rect 19740 17380 19796 17436
rect 19796 17380 19800 17436
rect 19736 17376 19800 17380
rect 19816 17436 19880 17440
rect 19816 17380 19820 17436
rect 19820 17380 19876 17436
rect 19876 17380 19880 17436
rect 19816 17376 19880 17380
rect 50296 17436 50360 17440
rect 50296 17380 50300 17436
rect 50300 17380 50356 17436
rect 50356 17380 50360 17436
rect 50296 17376 50360 17380
rect 50376 17436 50440 17440
rect 50376 17380 50380 17436
rect 50380 17380 50436 17436
rect 50436 17380 50440 17436
rect 50376 17376 50440 17380
rect 50456 17436 50520 17440
rect 50456 17380 50460 17436
rect 50460 17380 50516 17436
rect 50516 17380 50520 17436
rect 50456 17376 50520 17380
rect 50536 17436 50600 17440
rect 50536 17380 50540 17436
rect 50540 17380 50596 17436
rect 50596 17380 50600 17436
rect 50536 17376 50600 17380
rect 4216 16892 4280 16896
rect 4216 16836 4220 16892
rect 4220 16836 4276 16892
rect 4276 16836 4280 16892
rect 4216 16832 4280 16836
rect 4296 16892 4360 16896
rect 4296 16836 4300 16892
rect 4300 16836 4356 16892
rect 4356 16836 4360 16892
rect 4296 16832 4360 16836
rect 4376 16892 4440 16896
rect 4376 16836 4380 16892
rect 4380 16836 4436 16892
rect 4436 16836 4440 16892
rect 4376 16832 4440 16836
rect 4456 16892 4520 16896
rect 4456 16836 4460 16892
rect 4460 16836 4516 16892
rect 4516 16836 4520 16892
rect 4456 16832 4520 16836
rect 34936 16892 35000 16896
rect 34936 16836 34940 16892
rect 34940 16836 34996 16892
rect 34996 16836 35000 16892
rect 34936 16832 35000 16836
rect 35016 16892 35080 16896
rect 35016 16836 35020 16892
rect 35020 16836 35076 16892
rect 35076 16836 35080 16892
rect 35016 16832 35080 16836
rect 35096 16892 35160 16896
rect 35096 16836 35100 16892
rect 35100 16836 35156 16892
rect 35156 16836 35160 16892
rect 35096 16832 35160 16836
rect 35176 16892 35240 16896
rect 35176 16836 35180 16892
rect 35180 16836 35236 16892
rect 35236 16836 35240 16892
rect 35176 16832 35240 16836
rect 23428 16764 23492 16828
rect 19576 16348 19640 16352
rect 19576 16292 19580 16348
rect 19580 16292 19636 16348
rect 19636 16292 19640 16348
rect 19576 16288 19640 16292
rect 19656 16348 19720 16352
rect 19656 16292 19660 16348
rect 19660 16292 19716 16348
rect 19716 16292 19720 16348
rect 19656 16288 19720 16292
rect 19736 16348 19800 16352
rect 19736 16292 19740 16348
rect 19740 16292 19796 16348
rect 19796 16292 19800 16348
rect 19736 16288 19800 16292
rect 19816 16348 19880 16352
rect 19816 16292 19820 16348
rect 19820 16292 19876 16348
rect 19876 16292 19880 16348
rect 19816 16288 19880 16292
rect 50296 16348 50360 16352
rect 50296 16292 50300 16348
rect 50300 16292 50356 16348
rect 50356 16292 50360 16348
rect 50296 16288 50360 16292
rect 50376 16348 50440 16352
rect 50376 16292 50380 16348
rect 50380 16292 50436 16348
rect 50436 16292 50440 16348
rect 50376 16288 50440 16292
rect 50456 16348 50520 16352
rect 50456 16292 50460 16348
rect 50460 16292 50516 16348
rect 50516 16292 50520 16348
rect 50456 16288 50520 16292
rect 50536 16348 50600 16352
rect 50536 16292 50540 16348
rect 50540 16292 50596 16348
rect 50596 16292 50600 16348
rect 50536 16288 50600 16292
rect 4216 15804 4280 15808
rect 4216 15748 4220 15804
rect 4220 15748 4276 15804
rect 4276 15748 4280 15804
rect 4216 15744 4280 15748
rect 4296 15804 4360 15808
rect 4296 15748 4300 15804
rect 4300 15748 4356 15804
rect 4356 15748 4360 15804
rect 4296 15744 4360 15748
rect 4376 15804 4440 15808
rect 4376 15748 4380 15804
rect 4380 15748 4436 15804
rect 4436 15748 4440 15804
rect 4376 15744 4440 15748
rect 4456 15804 4520 15808
rect 4456 15748 4460 15804
rect 4460 15748 4516 15804
rect 4516 15748 4520 15804
rect 4456 15744 4520 15748
rect 34936 15804 35000 15808
rect 34936 15748 34940 15804
rect 34940 15748 34996 15804
rect 34996 15748 35000 15804
rect 34936 15744 35000 15748
rect 35016 15804 35080 15808
rect 35016 15748 35020 15804
rect 35020 15748 35076 15804
rect 35076 15748 35080 15804
rect 35016 15744 35080 15748
rect 35096 15804 35160 15808
rect 35096 15748 35100 15804
rect 35100 15748 35156 15804
rect 35156 15748 35160 15804
rect 35096 15744 35160 15748
rect 35176 15804 35240 15808
rect 35176 15748 35180 15804
rect 35180 15748 35236 15804
rect 35236 15748 35240 15804
rect 35176 15744 35240 15748
rect 21220 15268 21284 15332
rect 19576 15260 19640 15264
rect 19576 15204 19580 15260
rect 19580 15204 19636 15260
rect 19636 15204 19640 15260
rect 19576 15200 19640 15204
rect 19656 15260 19720 15264
rect 19656 15204 19660 15260
rect 19660 15204 19716 15260
rect 19716 15204 19720 15260
rect 19656 15200 19720 15204
rect 19736 15260 19800 15264
rect 19736 15204 19740 15260
rect 19740 15204 19796 15260
rect 19796 15204 19800 15260
rect 19736 15200 19800 15204
rect 19816 15260 19880 15264
rect 19816 15204 19820 15260
rect 19820 15204 19876 15260
rect 19876 15204 19880 15260
rect 19816 15200 19880 15204
rect 50296 15260 50360 15264
rect 50296 15204 50300 15260
rect 50300 15204 50356 15260
rect 50356 15204 50360 15260
rect 50296 15200 50360 15204
rect 50376 15260 50440 15264
rect 50376 15204 50380 15260
rect 50380 15204 50436 15260
rect 50436 15204 50440 15260
rect 50376 15200 50440 15204
rect 50456 15260 50520 15264
rect 50456 15204 50460 15260
rect 50460 15204 50516 15260
rect 50516 15204 50520 15260
rect 50456 15200 50520 15204
rect 50536 15260 50600 15264
rect 50536 15204 50540 15260
rect 50540 15204 50596 15260
rect 50596 15204 50600 15260
rect 50536 15200 50600 15204
rect 4216 14716 4280 14720
rect 4216 14660 4220 14716
rect 4220 14660 4276 14716
rect 4276 14660 4280 14716
rect 4216 14656 4280 14660
rect 4296 14716 4360 14720
rect 4296 14660 4300 14716
rect 4300 14660 4356 14716
rect 4356 14660 4360 14716
rect 4296 14656 4360 14660
rect 4376 14716 4440 14720
rect 4376 14660 4380 14716
rect 4380 14660 4436 14716
rect 4436 14660 4440 14716
rect 4376 14656 4440 14660
rect 4456 14716 4520 14720
rect 4456 14660 4460 14716
rect 4460 14660 4516 14716
rect 4516 14660 4520 14716
rect 4456 14656 4520 14660
rect 34936 14716 35000 14720
rect 34936 14660 34940 14716
rect 34940 14660 34996 14716
rect 34996 14660 35000 14716
rect 34936 14656 35000 14660
rect 35016 14716 35080 14720
rect 35016 14660 35020 14716
rect 35020 14660 35076 14716
rect 35076 14660 35080 14716
rect 35016 14656 35080 14660
rect 35096 14716 35160 14720
rect 35096 14660 35100 14716
rect 35100 14660 35156 14716
rect 35156 14660 35160 14716
rect 35096 14656 35160 14660
rect 35176 14716 35240 14720
rect 35176 14660 35180 14716
rect 35180 14660 35236 14716
rect 35236 14660 35240 14716
rect 35176 14656 35240 14660
rect 19576 14172 19640 14176
rect 19576 14116 19580 14172
rect 19580 14116 19636 14172
rect 19636 14116 19640 14172
rect 19576 14112 19640 14116
rect 19656 14172 19720 14176
rect 19656 14116 19660 14172
rect 19660 14116 19716 14172
rect 19716 14116 19720 14172
rect 19656 14112 19720 14116
rect 19736 14172 19800 14176
rect 19736 14116 19740 14172
rect 19740 14116 19796 14172
rect 19796 14116 19800 14172
rect 19736 14112 19800 14116
rect 19816 14172 19880 14176
rect 19816 14116 19820 14172
rect 19820 14116 19876 14172
rect 19876 14116 19880 14172
rect 19816 14112 19880 14116
rect 50296 14172 50360 14176
rect 50296 14116 50300 14172
rect 50300 14116 50356 14172
rect 50356 14116 50360 14172
rect 50296 14112 50360 14116
rect 50376 14172 50440 14176
rect 50376 14116 50380 14172
rect 50380 14116 50436 14172
rect 50436 14116 50440 14172
rect 50376 14112 50440 14116
rect 50456 14172 50520 14176
rect 50456 14116 50460 14172
rect 50460 14116 50516 14172
rect 50516 14116 50520 14172
rect 50456 14112 50520 14116
rect 50536 14172 50600 14176
rect 50536 14116 50540 14172
rect 50540 14116 50596 14172
rect 50596 14116 50600 14172
rect 50536 14112 50600 14116
rect 4216 13628 4280 13632
rect 4216 13572 4220 13628
rect 4220 13572 4276 13628
rect 4276 13572 4280 13628
rect 4216 13568 4280 13572
rect 4296 13628 4360 13632
rect 4296 13572 4300 13628
rect 4300 13572 4356 13628
rect 4356 13572 4360 13628
rect 4296 13568 4360 13572
rect 4376 13628 4440 13632
rect 4376 13572 4380 13628
rect 4380 13572 4436 13628
rect 4436 13572 4440 13628
rect 4376 13568 4440 13572
rect 4456 13628 4520 13632
rect 4456 13572 4460 13628
rect 4460 13572 4516 13628
rect 4516 13572 4520 13628
rect 4456 13568 4520 13572
rect 34936 13628 35000 13632
rect 34936 13572 34940 13628
rect 34940 13572 34996 13628
rect 34996 13572 35000 13628
rect 34936 13568 35000 13572
rect 35016 13628 35080 13632
rect 35016 13572 35020 13628
rect 35020 13572 35076 13628
rect 35076 13572 35080 13628
rect 35016 13568 35080 13572
rect 35096 13628 35160 13632
rect 35096 13572 35100 13628
rect 35100 13572 35156 13628
rect 35156 13572 35160 13628
rect 35096 13568 35160 13572
rect 35176 13628 35240 13632
rect 35176 13572 35180 13628
rect 35180 13572 35236 13628
rect 35236 13572 35240 13628
rect 35176 13568 35240 13572
rect 19576 13084 19640 13088
rect 19576 13028 19580 13084
rect 19580 13028 19636 13084
rect 19636 13028 19640 13084
rect 19576 13024 19640 13028
rect 19656 13084 19720 13088
rect 19656 13028 19660 13084
rect 19660 13028 19716 13084
rect 19716 13028 19720 13084
rect 19656 13024 19720 13028
rect 19736 13084 19800 13088
rect 19736 13028 19740 13084
rect 19740 13028 19796 13084
rect 19796 13028 19800 13084
rect 19736 13024 19800 13028
rect 19816 13084 19880 13088
rect 19816 13028 19820 13084
rect 19820 13028 19876 13084
rect 19876 13028 19880 13084
rect 19816 13024 19880 13028
rect 50296 13084 50360 13088
rect 50296 13028 50300 13084
rect 50300 13028 50356 13084
rect 50356 13028 50360 13084
rect 50296 13024 50360 13028
rect 50376 13084 50440 13088
rect 50376 13028 50380 13084
rect 50380 13028 50436 13084
rect 50436 13028 50440 13084
rect 50376 13024 50440 13028
rect 50456 13084 50520 13088
rect 50456 13028 50460 13084
rect 50460 13028 50516 13084
rect 50516 13028 50520 13084
rect 50456 13024 50520 13028
rect 50536 13084 50600 13088
rect 50536 13028 50540 13084
rect 50540 13028 50596 13084
rect 50596 13028 50600 13084
rect 50536 13024 50600 13028
rect 4216 12540 4280 12544
rect 4216 12484 4220 12540
rect 4220 12484 4276 12540
rect 4276 12484 4280 12540
rect 4216 12480 4280 12484
rect 4296 12540 4360 12544
rect 4296 12484 4300 12540
rect 4300 12484 4356 12540
rect 4356 12484 4360 12540
rect 4296 12480 4360 12484
rect 4376 12540 4440 12544
rect 4376 12484 4380 12540
rect 4380 12484 4436 12540
rect 4436 12484 4440 12540
rect 4376 12480 4440 12484
rect 4456 12540 4520 12544
rect 4456 12484 4460 12540
rect 4460 12484 4516 12540
rect 4516 12484 4520 12540
rect 4456 12480 4520 12484
rect 34936 12540 35000 12544
rect 34936 12484 34940 12540
rect 34940 12484 34996 12540
rect 34996 12484 35000 12540
rect 34936 12480 35000 12484
rect 35016 12540 35080 12544
rect 35016 12484 35020 12540
rect 35020 12484 35076 12540
rect 35076 12484 35080 12540
rect 35016 12480 35080 12484
rect 35096 12540 35160 12544
rect 35096 12484 35100 12540
rect 35100 12484 35156 12540
rect 35156 12484 35160 12540
rect 35096 12480 35160 12484
rect 35176 12540 35240 12544
rect 35176 12484 35180 12540
rect 35180 12484 35236 12540
rect 35236 12484 35240 12540
rect 35176 12480 35240 12484
rect 19576 11996 19640 12000
rect 19576 11940 19580 11996
rect 19580 11940 19636 11996
rect 19636 11940 19640 11996
rect 19576 11936 19640 11940
rect 19656 11996 19720 12000
rect 19656 11940 19660 11996
rect 19660 11940 19716 11996
rect 19716 11940 19720 11996
rect 19656 11936 19720 11940
rect 19736 11996 19800 12000
rect 19736 11940 19740 11996
rect 19740 11940 19796 11996
rect 19796 11940 19800 11996
rect 19736 11936 19800 11940
rect 19816 11996 19880 12000
rect 19816 11940 19820 11996
rect 19820 11940 19876 11996
rect 19876 11940 19880 11996
rect 19816 11936 19880 11940
rect 50296 11996 50360 12000
rect 50296 11940 50300 11996
rect 50300 11940 50356 11996
rect 50356 11940 50360 11996
rect 50296 11936 50360 11940
rect 50376 11996 50440 12000
rect 50376 11940 50380 11996
rect 50380 11940 50436 11996
rect 50436 11940 50440 11996
rect 50376 11936 50440 11940
rect 50456 11996 50520 12000
rect 50456 11940 50460 11996
rect 50460 11940 50516 11996
rect 50516 11940 50520 11996
rect 50456 11936 50520 11940
rect 50536 11996 50600 12000
rect 50536 11940 50540 11996
rect 50540 11940 50596 11996
rect 50596 11940 50600 11996
rect 50536 11936 50600 11940
rect 4216 11452 4280 11456
rect 4216 11396 4220 11452
rect 4220 11396 4276 11452
rect 4276 11396 4280 11452
rect 4216 11392 4280 11396
rect 4296 11452 4360 11456
rect 4296 11396 4300 11452
rect 4300 11396 4356 11452
rect 4356 11396 4360 11452
rect 4296 11392 4360 11396
rect 4376 11452 4440 11456
rect 4376 11396 4380 11452
rect 4380 11396 4436 11452
rect 4436 11396 4440 11452
rect 4376 11392 4440 11396
rect 4456 11452 4520 11456
rect 4456 11396 4460 11452
rect 4460 11396 4516 11452
rect 4516 11396 4520 11452
rect 4456 11392 4520 11396
rect 34936 11452 35000 11456
rect 34936 11396 34940 11452
rect 34940 11396 34996 11452
rect 34996 11396 35000 11452
rect 34936 11392 35000 11396
rect 35016 11452 35080 11456
rect 35016 11396 35020 11452
rect 35020 11396 35076 11452
rect 35076 11396 35080 11452
rect 35016 11392 35080 11396
rect 35096 11452 35160 11456
rect 35096 11396 35100 11452
rect 35100 11396 35156 11452
rect 35156 11396 35160 11452
rect 35096 11392 35160 11396
rect 35176 11452 35240 11456
rect 35176 11396 35180 11452
rect 35180 11396 35236 11452
rect 35236 11396 35240 11452
rect 35176 11392 35240 11396
rect 19576 10908 19640 10912
rect 19576 10852 19580 10908
rect 19580 10852 19636 10908
rect 19636 10852 19640 10908
rect 19576 10848 19640 10852
rect 19656 10908 19720 10912
rect 19656 10852 19660 10908
rect 19660 10852 19716 10908
rect 19716 10852 19720 10908
rect 19656 10848 19720 10852
rect 19736 10908 19800 10912
rect 19736 10852 19740 10908
rect 19740 10852 19796 10908
rect 19796 10852 19800 10908
rect 19736 10848 19800 10852
rect 19816 10908 19880 10912
rect 19816 10852 19820 10908
rect 19820 10852 19876 10908
rect 19876 10852 19880 10908
rect 19816 10848 19880 10852
rect 50296 10908 50360 10912
rect 50296 10852 50300 10908
rect 50300 10852 50356 10908
rect 50356 10852 50360 10908
rect 50296 10848 50360 10852
rect 50376 10908 50440 10912
rect 50376 10852 50380 10908
rect 50380 10852 50436 10908
rect 50436 10852 50440 10908
rect 50376 10848 50440 10852
rect 50456 10908 50520 10912
rect 50456 10852 50460 10908
rect 50460 10852 50516 10908
rect 50516 10852 50520 10908
rect 50456 10848 50520 10852
rect 50536 10908 50600 10912
rect 50536 10852 50540 10908
rect 50540 10852 50596 10908
rect 50596 10852 50600 10908
rect 50536 10848 50600 10852
rect 4216 10364 4280 10368
rect 4216 10308 4220 10364
rect 4220 10308 4276 10364
rect 4276 10308 4280 10364
rect 4216 10304 4280 10308
rect 4296 10364 4360 10368
rect 4296 10308 4300 10364
rect 4300 10308 4356 10364
rect 4356 10308 4360 10364
rect 4296 10304 4360 10308
rect 4376 10364 4440 10368
rect 4376 10308 4380 10364
rect 4380 10308 4436 10364
rect 4436 10308 4440 10364
rect 4376 10304 4440 10308
rect 4456 10364 4520 10368
rect 4456 10308 4460 10364
rect 4460 10308 4516 10364
rect 4516 10308 4520 10364
rect 4456 10304 4520 10308
rect 34936 10364 35000 10368
rect 34936 10308 34940 10364
rect 34940 10308 34996 10364
rect 34996 10308 35000 10364
rect 34936 10304 35000 10308
rect 35016 10364 35080 10368
rect 35016 10308 35020 10364
rect 35020 10308 35076 10364
rect 35076 10308 35080 10364
rect 35016 10304 35080 10308
rect 35096 10364 35160 10368
rect 35096 10308 35100 10364
rect 35100 10308 35156 10364
rect 35156 10308 35160 10364
rect 35096 10304 35160 10308
rect 35176 10364 35240 10368
rect 35176 10308 35180 10364
rect 35180 10308 35236 10364
rect 35236 10308 35240 10364
rect 35176 10304 35240 10308
rect 19576 9820 19640 9824
rect 19576 9764 19580 9820
rect 19580 9764 19636 9820
rect 19636 9764 19640 9820
rect 19576 9760 19640 9764
rect 19656 9820 19720 9824
rect 19656 9764 19660 9820
rect 19660 9764 19716 9820
rect 19716 9764 19720 9820
rect 19656 9760 19720 9764
rect 19736 9820 19800 9824
rect 19736 9764 19740 9820
rect 19740 9764 19796 9820
rect 19796 9764 19800 9820
rect 19736 9760 19800 9764
rect 19816 9820 19880 9824
rect 19816 9764 19820 9820
rect 19820 9764 19876 9820
rect 19876 9764 19880 9820
rect 19816 9760 19880 9764
rect 50296 9820 50360 9824
rect 50296 9764 50300 9820
rect 50300 9764 50356 9820
rect 50356 9764 50360 9820
rect 50296 9760 50360 9764
rect 50376 9820 50440 9824
rect 50376 9764 50380 9820
rect 50380 9764 50436 9820
rect 50436 9764 50440 9820
rect 50376 9760 50440 9764
rect 50456 9820 50520 9824
rect 50456 9764 50460 9820
rect 50460 9764 50516 9820
rect 50516 9764 50520 9820
rect 50456 9760 50520 9764
rect 50536 9820 50600 9824
rect 50536 9764 50540 9820
rect 50540 9764 50596 9820
rect 50596 9764 50600 9820
rect 50536 9760 50600 9764
rect 4216 9276 4280 9280
rect 4216 9220 4220 9276
rect 4220 9220 4276 9276
rect 4276 9220 4280 9276
rect 4216 9216 4280 9220
rect 4296 9276 4360 9280
rect 4296 9220 4300 9276
rect 4300 9220 4356 9276
rect 4356 9220 4360 9276
rect 4296 9216 4360 9220
rect 4376 9276 4440 9280
rect 4376 9220 4380 9276
rect 4380 9220 4436 9276
rect 4436 9220 4440 9276
rect 4376 9216 4440 9220
rect 4456 9276 4520 9280
rect 4456 9220 4460 9276
rect 4460 9220 4516 9276
rect 4516 9220 4520 9276
rect 4456 9216 4520 9220
rect 34936 9276 35000 9280
rect 34936 9220 34940 9276
rect 34940 9220 34996 9276
rect 34996 9220 35000 9276
rect 34936 9216 35000 9220
rect 35016 9276 35080 9280
rect 35016 9220 35020 9276
rect 35020 9220 35076 9276
rect 35076 9220 35080 9276
rect 35016 9216 35080 9220
rect 35096 9276 35160 9280
rect 35096 9220 35100 9276
rect 35100 9220 35156 9276
rect 35156 9220 35160 9276
rect 35096 9216 35160 9220
rect 35176 9276 35240 9280
rect 35176 9220 35180 9276
rect 35180 9220 35236 9276
rect 35236 9220 35240 9276
rect 35176 9216 35240 9220
rect 19576 8732 19640 8736
rect 19576 8676 19580 8732
rect 19580 8676 19636 8732
rect 19636 8676 19640 8732
rect 19576 8672 19640 8676
rect 19656 8732 19720 8736
rect 19656 8676 19660 8732
rect 19660 8676 19716 8732
rect 19716 8676 19720 8732
rect 19656 8672 19720 8676
rect 19736 8732 19800 8736
rect 19736 8676 19740 8732
rect 19740 8676 19796 8732
rect 19796 8676 19800 8732
rect 19736 8672 19800 8676
rect 19816 8732 19880 8736
rect 19816 8676 19820 8732
rect 19820 8676 19876 8732
rect 19876 8676 19880 8732
rect 19816 8672 19880 8676
rect 50296 8732 50360 8736
rect 50296 8676 50300 8732
rect 50300 8676 50356 8732
rect 50356 8676 50360 8732
rect 50296 8672 50360 8676
rect 50376 8732 50440 8736
rect 50376 8676 50380 8732
rect 50380 8676 50436 8732
rect 50436 8676 50440 8732
rect 50376 8672 50440 8676
rect 50456 8732 50520 8736
rect 50456 8676 50460 8732
rect 50460 8676 50516 8732
rect 50516 8676 50520 8732
rect 50456 8672 50520 8676
rect 50536 8732 50600 8736
rect 50536 8676 50540 8732
rect 50540 8676 50596 8732
rect 50596 8676 50600 8732
rect 50536 8672 50600 8676
rect 4216 8188 4280 8192
rect 4216 8132 4220 8188
rect 4220 8132 4276 8188
rect 4276 8132 4280 8188
rect 4216 8128 4280 8132
rect 4296 8188 4360 8192
rect 4296 8132 4300 8188
rect 4300 8132 4356 8188
rect 4356 8132 4360 8188
rect 4296 8128 4360 8132
rect 4376 8188 4440 8192
rect 4376 8132 4380 8188
rect 4380 8132 4436 8188
rect 4436 8132 4440 8188
rect 4376 8128 4440 8132
rect 4456 8188 4520 8192
rect 4456 8132 4460 8188
rect 4460 8132 4516 8188
rect 4516 8132 4520 8188
rect 4456 8128 4520 8132
rect 34936 8188 35000 8192
rect 34936 8132 34940 8188
rect 34940 8132 34996 8188
rect 34996 8132 35000 8188
rect 34936 8128 35000 8132
rect 35016 8188 35080 8192
rect 35016 8132 35020 8188
rect 35020 8132 35076 8188
rect 35076 8132 35080 8188
rect 35016 8128 35080 8132
rect 35096 8188 35160 8192
rect 35096 8132 35100 8188
rect 35100 8132 35156 8188
rect 35156 8132 35160 8188
rect 35096 8128 35160 8132
rect 35176 8188 35240 8192
rect 35176 8132 35180 8188
rect 35180 8132 35236 8188
rect 35236 8132 35240 8188
rect 35176 8128 35240 8132
rect 19576 7644 19640 7648
rect 19576 7588 19580 7644
rect 19580 7588 19636 7644
rect 19636 7588 19640 7644
rect 19576 7584 19640 7588
rect 19656 7644 19720 7648
rect 19656 7588 19660 7644
rect 19660 7588 19716 7644
rect 19716 7588 19720 7644
rect 19656 7584 19720 7588
rect 19736 7644 19800 7648
rect 19736 7588 19740 7644
rect 19740 7588 19796 7644
rect 19796 7588 19800 7644
rect 19736 7584 19800 7588
rect 19816 7644 19880 7648
rect 19816 7588 19820 7644
rect 19820 7588 19876 7644
rect 19876 7588 19880 7644
rect 19816 7584 19880 7588
rect 50296 7644 50360 7648
rect 50296 7588 50300 7644
rect 50300 7588 50356 7644
rect 50356 7588 50360 7644
rect 50296 7584 50360 7588
rect 50376 7644 50440 7648
rect 50376 7588 50380 7644
rect 50380 7588 50436 7644
rect 50436 7588 50440 7644
rect 50376 7584 50440 7588
rect 50456 7644 50520 7648
rect 50456 7588 50460 7644
rect 50460 7588 50516 7644
rect 50516 7588 50520 7644
rect 50456 7584 50520 7588
rect 50536 7644 50600 7648
rect 50536 7588 50540 7644
rect 50540 7588 50596 7644
rect 50596 7588 50600 7644
rect 50536 7584 50600 7588
rect 4216 7100 4280 7104
rect 4216 7044 4220 7100
rect 4220 7044 4276 7100
rect 4276 7044 4280 7100
rect 4216 7040 4280 7044
rect 4296 7100 4360 7104
rect 4296 7044 4300 7100
rect 4300 7044 4356 7100
rect 4356 7044 4360 7100
rect 4296 7040 4360 7044
rect 4376 7100 4440 7104
rect 4376 7044 4380 7100
rect 4380 7044 4436 7100
rect 4436 7044 4440 7100
rect 4376 7040 4440 7044
rect 4456 7100 4520 7104
rect 4456 7044 4460 7100
rect 4460 7044 4516 7100
rect 4516 7044 4520 7100
rect 4456 7040 4520 7044
rect 34936 7100 35000 7104
rect 34936 7044 34940 7100
rect 34940 7044 34996 7100
rect 34996 7044 35000 7100
rect 34936 7040 35000 7044
rect 35016 7100 35080 7104
rect 35016 7044 35020 7100
rect 35020 7044 35076 7100
rect 35076 7044 35080 7100
rect 35016 7040 35080 7044
rect 35096 7100 35160 7104
rect 35096 7044 35100 7100
rect 35100 7044 35156 7100
rect 35156 7044 35160 7100
rect 35096 7040 35160 7044
rect 35176 7100 35240 7104
rect 35176 7044 35180 7100
rect 35180 7044 35236 7100
rect 35236 7044 35240 7100
rect 35176 7040 35240 7044
rect 19576 6556 19640 6560
rect 19576 6500 19580 6556
rect 19580 6500 19636 6556
rect 19636 6500 19640 6556
rect 19576 6496 19640 6500
rect 19656 6556 19720 6560
rect 19656 6500 19660 6556
rect 19660 6500 19716 6556
rect 19716 6500 19720 6556
rect 19656 6496 19720 6500
rect 19736 6556 19800 6560
rect 19736 6500 19740 6556
rect 19740 6500 19796 6556
rect 19796 6500 19800 6556
rect 19736 6496 19800 6500
rect 19816 6556 19880 6560
rect 19816 6500 19820 6556
rect 19820 6500 19876 6556
rect 19876 6500 19880 6556
rect 19816 6496 19880 6500
rect 50296 6556 50360 6560
rect 50296 6500 50300 6556
rect 50300 6500 50356 6556
rect 50356 6500 50360 6556
rect 50296 6496 50360 6500
rect 50376 6556 50440 6560
rect 50376 6500 50380 6556
rect 50380 6500 50436 6556
rect 50436 6500 50440 6556
rect 50376 6496 50440 6500
rect 50456 6556 50520 6560
rect 50456 6500 50460 6556
rect 50460 6500 50516 6556
rect 50516 6500 50520 6556
rect 50456 6496 50520 6500
rect 50536 6556 50600 6560
rect 50536 6500 50540 6556
rect 50540 6500 50596 6556
rect 50596 6500 50600 6556
rect 50536 6496 50600 6500
rect 4216 6012 4280 6016
rect 4216 5956 4220 6012
rect 4220 5956 4276 6012
rect 4276 5956 4280 6012
rect 4216 5952 4280 5956
rect 4296 6012 4360 6016
rect 4296 5956 4300 6012
rect 4300 5956 4356 6012
rect 4356 5956 4360 6012
rect 4296 5952 4360 5956
rect 4376 6012 4440 6016
rect 4376 5956 4380 6012
rect 4380 5956 4436 6012
rect 4436 5956 4440 6012
rect 4376 5952 4440 5956
rect 4456 6012 4520 6016
rect 4456 5956 4460 6012
rect 4460 5956 4516 6012
rect 4516 5956 4520 6012
rect 4456 5952 4520 5956
rect 34936 6012 35000 6016
rect 34936 5956 34940 6012
rect 34940 5956 34996 6012
rect 34996 5956 35000 6012
rect 34936 5952 35000 5956
rect 35016 6012 35080 6016
rect 35016 5956 35020 6012
rect 35020 5956 35076 6012
rect 35076 5956 35080 6012
rect 35016 5952 35080 5956
rect 35096 6012 35160 6016
rect 35096 5956 35100 6012
rect 35100 5956 35156 6012
rect 35156 5956 35160 6012
rect 35096 5952 35160 5956
rect 35176 6012 35240 6016
rect 35176 5956 35180 6012
rect 35180 5956 35236 6012
rect 35236 5956 35240 6012
rect 35176 5952 35240 5956
rect 19576 5468 19640 5472
rect 19576 5412 19580 5468
rect 19580 5412 19636 5468
rect 19636 5412 19640 5468
rect 19576 5408 19640 5412
rect 19656 5468 19720 5472
rect 19656 5412 19660 5468
rect 19660 5412 19716 5468
rect 19716 5412 19720 5468
rect 19656 5408 19720 5412
rect 19736 5468 19800 5472
rect 19736 5412 19740 5468
rect 19740 5412 19796 5468
rect 19796 5412 19800 5468
rect 19736 5408 19800 5412
rect 19816 5468 19880 5472
rect 19816 5412 19820 5468
rect 19820 5412 19876 5468
rect 19876 5412 19880 5468
rect 19816 5408 19880 5412
rect 50296 5468 50360 5472
rect 50296 5412 50300 5468
rect 50300 5412 50356 5468
rect 50356 5412 50360 5468
rect 50296 5408 50360 5412
rect 50376 5468 50440 5472
rect 50376 5412 50380 5468
rect 50380 5412 50436 5468
rect 50436 5412 50440 5468
rect 50376 5408 50440 5412
rect 50456 5468 50520 5472
rect 50456 5412 50460 5468
rect 50460 5412 50516 5468
rect 50516 5412 50520 5468
rect 50456 5408 50520 5412
rect 50536 5468 50600 5472
rect 50536 5412 50540 5468
rect 50540 5412 50596 5468
rect 50596 5412 50600 5468
rect 50536 5408 50600 5412
rect 4216 4924 4280 4928
rect 4216 4868 4220 4924
rect 4220 4868 4276 4924
rect 4276 4868 4280 4924
rect 4216 4864 4280 4868
rect 4296 4924 4360 4928
rect 4296 4868 4300 4924
rect 4300 4868 4356 4924
rect 4356 4868 4360 4924
rect 4296 4864 4360 4868
rect 4376 4924 4440 4928
rect 4376 4868 4380 4924
rect 4380 4868 4436 4924
rect 4436 4868 4440 4924
rect 4376 4864 4440 4868
rect 4456 4924 4520 4928
rect 4456 4868 4460 4924
rect 4460 4868 4516 4924
rect 4516 4868 4520 4924
rect 4456 4864 4520 4868
rect 34936 4924 35000 4928
rect 34936 4868 34940 4924
rect 34940 4868 34996 4924
rect 34996 4868 35000 4924
rect 34936 4864 35000 4868
rect 35016 4924 35080 4928
rect 35016 4868 35020 4924
rect 35020 4868 35076 4924
rect 35076 4868 35080 4924
rect 35016 4864 35080 4868
rect 35096 4924 35160 4928
rect 35096 4868 35100 4924
rect 35100 4868 35156 4924
rect 35156 4868 35160 4924
rect 35096 4864 35160 4868
rect 35176 4924 35240 4928
rect 35176 4868 35180 4924
rect 35180 4868 35236 4924
rect 35236 4868 35240 4924
rect 35176 4864 35240 4868
rect 19576 4380 19640 4384
rect 19576 4324 19580 4380
rect 19580 4324 19636 4380
rect 19636 4324 19640 4380
rect 19576 4320 19640 4324
rect 19656 4380 19720 4384
rect 19656 4324 19660 4380
rect 19660 4324 19716 4380
rect 19716 4324 19720 4380
rect 19656 4320 19720 4324
rect 19736 4380 19800 4384
rect 19736 4324 19740 4380
rect 19740 4324 19796 4380
rect 19796 4324 19800 4380
rect 19736 4320 19800 4324
rect 19816 4380 19880 4384
rect 19816 4324 19820 4380
rect 19820 4324 19876 4380
rect 19876 4324 19880 4380
rect 19816 4320 19880 4324
rect 50296 4380 50360 4384
rect 50296 4324 50300 4380
rect 50300 4324 50356 4380
rect 50356 4324 50360 4380
rect 50296 4320 50360 4324
rect 50376 4380 50440 4384
rect 50376 4324 50380 4380
rect 50380 4324 50436 4380
rect 50436 4324 50440 4380
rect 50376 4320 50440 4324
rect 50456 4380 50520 4384
rect 50456 4324 50460 4380
rect 50460 4324 50516 4380
rect 50516 4324 50520 4380
rect 50456 4320 50520 4324
rect 50536 4380 50600 4384
rect 50536 4324 50540 4380
rect 50540 4324 50596 4380
rect 50596 4324 50600 4380
rect 50536 4320 50600 4324
rect 4216 3836 4280 3840
rect 4216 3780 4220 3836
rect 4220 3780 4276 3836
rect 4276 3780 4280 3836
rect 4216 3776 4280 3780
rect 4296 3836 4360 3840
rect 4296 3780 4300 3836
rect 4300 3780 4356 3836
rect 4356 3780 4360 3836
rect 4296 3776 4360 3780
rect 4376 3836 4440 3840
rect 4376 3780 4380 3836
rect 4380 3780 4436 3836
rect 4436 3780 4440 3836
rect 4376 3776 4440 3780
rect 4456 3836 4520 3840
rect 4456 3780 4460 3836
rect 4460 3780 4516 3836
rect 4516 3780 4520 3836
rect 4456 3776 4520 3780
rect 34936 3836 35000 3840
rect 34936 3780 34940 3836
rect 34940 3780 34996 3836
rect 34996 3780 35000 3836
rect 34936 3776 35000 3780
rect 35016 3836 35080 3840
rect 35016 3780 35020 3836
rect 35020 3780 35076 3836
rect 35076 3780 35080 3836
rect 35016 3776 35080 3780
rect 35096 3836 35160 3840
rect 35096 3780 35100 3836
rect 35100 3780 35156 3836
rect 35156 3780 35160 3836
rect 35096 3776 35160 3780
rect 35176 3836 35240 3840
rect 35176 3780 35180 3836
rect 35180 3780 35236 3836
rect 35236 3780 35240 3836
rect 35176 3776 35240 3780
rect 19576 3292 19640 3296
rect 19576 3236 19580 3292
rect 19580 3236 19636 3292
rect 19636 3236 19640 3292
rect 19576 3232 19640 3236
rect 19656 3292 19720 3296
rect 19656 3236 19660 3292
rect 19660 3236 19716 3292
rect 19716 3236 19720 3292
rect 19656 3232 19720 3236
rect 19736 3292 19800 3296
rect 19736 3236 19740 3292
rect 19740 3236 19796 3292
rect 19796 3236 19800 3292
rect 19736 3232 19800 3236
rect 19816 3292 19880 3296
rect 19816 3236 19820 3292
rect 19820 3236 19876 3292
rect 19876 3236 19880 3292
rect 19816 3232 19880 3236
rect 50296 3292 50360 3296
rect 50296 3236 50300 3292
rect 50300 3236 50356 3292
rect 50356 3236 50360 3292
rect 50296 3232 50360 3236
rect 50376 3292 50440 3296
rect 50376 3236 50380 3292
rect 50380 3236 50436 3292
rect 50436 3236 50440 3292
rect 50376 3232 50440 3236
rect 50456 3292 50520 3296
rect 50456 3236 50460 3292
rect 50460 3236 50516 3292
rect 50516 3236 50520 3292
rect 50456 3232 50520 3236
rect 50536 3292 50600 3296
rect 50536 3236 50540 3292
rect 50540 3236 50596 3292
rect 50596 3236 50600 3292
rect 50536 3232 50600 3236
rect 4216 2748 4280 2752
rect 4216 2692 4220 2748
rect 4220 2692 4276 2748
rect 4276 2692 4280 2748
rect 4216 2688 4280 2692
rect 4296 2748 4360 2752
rect 4296 2692 4300 2748
rect 4300 2692 4356 2748
rect 4356 2692 4360 2748
rect 4296 2688 4360 2692
rect 4376 2748 4440 2752
rect 4376 2692 4380 2748
rect 4380 2692 4436 2748
rect 4436 2692 4440 2748
rect 4376 2688 4440 2692
rect 4456 2748 4520 2752
rect 4456 2692 4460 2748
rect 4460 2692 4516 2748
rect 4516 2692 4520 2748
rect 4456 2688 4520 2692
rect 34936 2748 35000 2752
rect 34936 2692 34940 2748
rect 34940 2692 34996 2748
rect 34996 2692 35000 2748
rect 34936 2688 35000 2692
rect 35016 2748 35080 2752
rect 35016 2692 35020 2748
rect 35020 2692 35076 2748
rect 35076 2692 35080 2748
rect 35016 2688 35080 2692
rect 35096 2748 35160 2752
rect 35096 2692 35100 2748
rect 35100 2692 35156 2748
rect 35156 2692 35160 2748
rect 35096 2688 35160 2692
rect 35176 2748 35240 2752
rect 35176 2692 35180 2748
rect 35180 2692 35236 2748
rect 35236 2692 35240 2748
rect 35176 2688 35240 2692
rect 19576 2204 19640 2208
rect 19576 2148 19580 2204
rect 19580 2148 19636 2204
rect 19636 2148 19640 2204
rect 19576 2144 19640 2148
rect 19656 2204 19720 2208
rect 19656 2148 19660 2204
rect 19660 2148 19716 2204
rect 19716 2148 19720 2204
rect 19656 2144 19720 2148
rect 19736 2204 19800 2208
rect 19736 2148 19740 2204
rect 19740 2148 19796 2204
rect 19796 2148 19800 2204
rect 19736 2144 19800 2148
rect 19816 2204 19880 2208
rect 19816 2148 19820 2204
rect 19820 2148 19876 2204
rect 19876 2148 19880 2204
rect 19816 2144 19880 2148
rect 50296 2204 50360 2208
rect 50296 2148 50300 2204
rect 50300 2148 50356 2204
rect 50356 2148 50360 2204
rect 50296 2144 50360 2148
rect 50376 2204 50440 2208
rect 50376 2148 50380 2204
rect 50380 2148 50436 2204
rect 50436 2148 50440 2204
rect 50376 2144 50440 2148
rect 50456 2204 50520 2208
rect 50456 2148 50460 2204
rect 50460 2148 50516 2204
rect 50516 2148 50520 2204
rect 50456 2144 50520 2148
rect 50536 2204 50600 2208
rect 50536 2148 50540 2204
rect 50540 2148 50596 2204
rect 50596 2148 50600 2204
rect 50536 2144 50600 2148
<< metal4 >>
rect 4208 37568 4528 37584
rect 4208 37504 4216 37568
rect 4280 37504 4296 37568
rect 4360 37504 4376 37568
rect 4440 37504 4456 37568
rect 4520 37504 4528 37568
rect 4208 36480 4528 37504
rect 4208 36416 4216 36480
rect 4280 36416 4296 36480
rect 4360 36416 4376 36480
rect 4440 36416 4456 36480
rect 4520 36416 4528 36480
rect 4208 35392 4528 36416
rect 4208 35328 4216 35392
rect 4280 35328 4296 35392
rect 4360 35328 4376 35392
rect 4440 35328 4456 35392
rect 4520 35328 4528 35392
rect 4208 34304 4528 35328
rect 4208 34240 4216 34304
rect 4280 34240 4296 34304
rect 4360 34240 4376 34304
rect 4440 34240 4456 34304
rect 4520 34240 4528 34304
rect 4208 33216 4528 34240
rect 4208 33152 4216 33216
rect 4280 33152 4296 33216
rect 4360 33152 4376 33216
rect 4440 33152 4456 33216
rect 4520 33152 4528 33216
rect 4208 32128 4528 33152
rect 4208 32064 4216 32128
rect 4280 32064 4296 32128
rect 4360 32064 4376 32128
rect 4440 32064 4456 32128
rect 4520 32064 4528 32128
rect 4208 31040 4528 32064
rect 4208 30976 4216 31040
rect 4280 30976 4296 31040
rect 4360 30976 4376 31040
rect 4440 30976 4456 31040
rect 4520 30976 4528 31040
rect 4208 29952 4528 30976
rect 4208 29888 4216 29952
rect 4280 29888 4296 29952
rect 4360 29888 4376 29952
rect 4440 29888 4456 29952
rect 4520 29888 4528 29952
rect 4208 28864 4528 29888
rect 4208 28800 4216 28864
rect 4280 28800 4296 28864
rect 4360 28800 4376 28864
rect 4440 28800 4456 28864
rect 4520 28800 4528 28864
rect 4208 27776 4528 28800
rect 4208 27712 4216 27776
rect 4280 27712 4296 27776
rect 4360 27712 4376 27776
rect 4440 27712 4456 27776
rect 4520 27712 4528 27776
rect 4208 26688 4528 27712
rect 4208 26624 4216 26688
rect 4280 26624 4296 26688
rect 4360 26624 4376 26688
rect 4440 26624 4456 26688
rect 4520 26624 4528 26688
rect 4208 25600 4528 26624
rect 4208 25536 4216 25600
rect 4280 25536 4296 25600
rect 4360 25536 4376 25600
rect 4440 25536 4456 25600
rect 4520 25536 4528 25600
rect 4208 24512 4528 25536
rect 4208 24448 4216 24512
rect 4280 24448 4296 24512
rect 4360 24448 4376 24512
rect 4440 24448 4456 24512
rect 4520 24448 4528 24512
rect 4208 23424 4528 24448
rect 4208 23360 4216 23424
rect 4280 23360 4296 23424
rect 4360 23360 4376 23424
rect 4440 23360 4456 23424
rect 4520 23360 4528 23424
rect 4208 22336 4528 23360
rect 4208 22272 4216 22336
rect 4280 22272 4296 22336
rect 4360 22272 4376 22336
rect 4440 22272 4456 22336
rect 4520 22272 4528 22336
rect 4208 21248 4528 22272
rect 4208 21184 4216 21248
rect 4280 21184 4296 21248
rect 4360 21184 4376 21248
rect 4440 21184 4456 21248
rect 4520 21184 4528 21248
rect 4208 20160 4528 21184
rect 4208 20096 4216 20160
rect 4280 20096 4296 20160
rect 4360 20096 4376 20160
rect 4440 20096 4456 20160
rect 4520 20096 4528 20160
rect 4208 19072 4528 20096
rect 4208 19008 4216 19072
rect 4280 19008 4296 19072
rect 4360 19008 4376 19072
rect 4440 19008 4456 19072
rect 4520 19008 4528 19072
rect 4208 17984 4528 19008
rect 4208 17920 4216 17984
rect 4280 17920 4296 17984
rect 4360 17920 4376 17984
rect 4440 17920 4456 17984
rect 4520 17920 4528 17984
rect 4208 16896 4528 17920
rect 4208 16832 4216 16896
rect 4280 16832 4296 16896
rect 4360 16832 4376 16896
rect 4440 16832 4456 16896
rect 4520 16832 4528 16896
rect 4208 15808 4528 16832
rect 4208 15744 4216 15808
rect 4280 15744 4296 15808
rect 4360 15744 4376 15808
rect 4440 15744 4456 15808
rect 4520 15744 4528 15808
rect 4208 14720 4528 15744
rect 4208 14656 4216 14720
rect 4280 14656 4296 14720
rect 4360 14656 4376 14720
rect 4440 14656 4456 14720
rect 4520 14656 4528 14720
rect 4208 13632 4528 14656
rect 4208 13568 4216 13632
rect 4280 13568 4296 13632
rect 4360 13568 4376 13632
rect 4440 13568 4456 13632
rect 4520 13568 4528 13632
rect 4208 12544 4528 13568
rect 4208 12480 4216 12544
rect 4280 12480 4296 12544
rect 4360 12480 4376 12544
rect 4440 12480 4456 12544
rect 4520 12480 4528 12544
rect 4208 11456 4528 12480
rect 4208 11392 4216 11456
rect 4280 11392 4296 11456
rect 4360 11392 4376 11456
rect 4440 11392 4456 11456
rect 4520 11392 4528 11456
rect 4208 10368 4528 11392
rect 4208 10304 4216 10368
rect 4280 10304 4296 10368
rect 4360 10304 4376 10368
rect 4440 10304 4456 10368
rect 4520 10304 4528 10368
rect 4208 9280 4528 10304
rect 4208 9216 4216 9280
rect 4280 9216 4296 9280
rect 4360 9216 4376 9280
rect 4440 9216 4456 9280
rect 4520 9216 4528 9280
rect 4208 8192 4528 9216
rect 4208 8128 4216 8192
rect 4280 8128 4296 8192
rect 4360 8128 4376 8192
rect 4440 8128 4456 8192
rect 4520 8128 4528 8192
rect 4208 7104 4528 8128
rect 4208 7040 4216 7104
rect 4280 7040 4296 7104
rect 4360 7040 4376 7104
rect 4440 7040 4456 7104
rect 4520 7040 4528 7104
rect 4208 6016 4528 7040
rect 4208 5952 4216 6016
rect 4280 5952 4296 6016
rect 4360 5952 4376 6016
rect 4440 5952 4456 6016
rect 4520 5952 4528 6016
rect 4208 4928 4528 5952
rect 4208 4864 4216 4928
rect 4280 4864 4296 4928
rect 4360 4864 4376 4928
rect 4440 4864 4456 4928
rect 4520 4864 4528 4928
rect 4208 3840 4528 4864
rect 4208 3776 4216 3840
rect 4280 3776 4296 3840
rect 4360 3776 4376 3840
rect 4440 3776 4456 3840
rect 4520 3776 4528 3840
rect 4208 2752 4528 3776
rect 4208 2688 4216 2752
rect 4280 2688 4296 2752
rect 4360 2688 4376 2752
rect 4440 2688 4456 2752
rect 4520 2688 4528 2752
rect 4208 2128 4528 2688
rect 19568 37024 19888 37584
rect 19568 36960 19576 37024
rect 19640 36960 19656 37024
rect 19720 36960 19736 37024
rect 19800 36960 19816 37024
rect 19880 36960 19888 37024
rect 19568 35936 19888 36960
rect 19568 35872 19576 35936
rect 19640 35872 19656 35936
rect 19720 35872 19736 35936
rect 19800 35872 19816 35936
rect 19880 35872 19888 35936
rect 19568 34848 19888 35872
rect 19568 34784 19576 34848
rect 19640 34784 19656 34848
rect 19720 34784 19736 34848
rect 19800 34784 19816 34848
rect 19880 34784 19888 34848
rect 19568 33760 19888 34784
rect 19568 33696 19576 33760
rect 19640 33696 19656 33760
rect 19720 33696 19736 33760
rect 19800 33696 19816 33760
rect 19880 33696 19888 33760
rect 19568 32672 19888 33696
rect 19568 32608 19576 32672
rect 19640 32608 19656 32672
rect 19720 32608 19736 32672
rect 19800 32608 19816 32672
rect 19880 32608 19888 32672
rect 19568 31584 19888 32608
rect 19568 31520 19576 31584
rect 19640 31520 19656 31584
rect 19720 31520 19736 31584
rect 19800 31520 19816 31584
rect 19880 31520 19888 31584
rect 19568 30496 19888 31520
rect 19568 30432 19576 30496
rect 19640 30432 19656 30496
rect 19720 30432 19736 30496
rect 19800 30432 19816 30496
rect 19880 30432 19888 30496
rect 19568 29408 19888 30432
rect 19568 29344 19576 29408
rect 19640 29344 19656 29408
rect 19720 29344 19736 29408
rect 19800 29344 19816 29408
rect 19880 29344 19888 29408
rect 19568 28320 19888 29344
rect 19568 28256 19576 28320
rect 19640 28256 19656 28320
rect 19720 28256 19736 28320
rect 19800 28256 19816 28320
rect 19880 28256 19888 28320
rect 19568 27232 19888 28256
rect 19568 27168 19576 27232
rect 19640 27168 19656 27232
rect 19720 27168 19736 27232
rect 19800 27168 19816 27232
rect 19880 27168 19888 27232
rect 19568 26144 19888 27168
rect 34928 37568 35248 37584
rect 34928 37504 34936 37568
rect 35000 37504 35016 37568
rect 35080 37504 35096 37568
rect 35160 37504 35176 37568
rect 35240 37504 35248 37568
rect 34928 36480 35248 37504
rect 34928 36416 34936 36480
rect 35000 36416 35016 36480
rect 35080 36416 35096 36480
rect 35160 36416 35176 36480
rect 35240 36416 35248 36480
rect 34928 35392 35248 36416
rect 34928 35328 34936 35392
rect 35000 35328 35016 35392
rect 35080 35328 35096 35392
rect 35160 35328 35176 35392
rect 35240 35328 35248 35392
rect 34928 34304 35248 35328
rect 34928 34240 34936 34304
rect 35000 34240 35016 34304
rect 35080 34240 35096 34304
rect 35160 34240 35176 34304
rect 35240 34240 35248 34304
rect 34928 33216 35248 34240
rect 34928 33152 34936 33216
rect 35000 33152 35016 33216
rect 35080 33152 35096 33216
rect 35160 33152 35176 33216
rect 35240 33152 35248 33216
rect 34928 32128 35248 33152
rect 34928 32064 34936 32128
rect 35000 32064 35016 32128
rect 35080 32064 35096 32128
rect 35160 32064 35176 32128
rect 35240 32064 35248 32128
rect 34928 31040 35248 32064
rect 34928 30976 34936 31040
rect 35000 30976 35016 31040
rect 35080 30976 35096 31040
rect 35160 30976 35176 31040
rect 35240 30976 35248 31040
rect 34928 29952 35248 30976
rect 34928 29888 34936 29952
rect 35000 29888 35016 29952
rect 35080 29888 35096 29952
rect 35160 29888 35176 29952
rect 35240 29888 35248 29952
rect 34928 28864 35248 29888
rect 34928 28800 34936 28864
rect 35000 28800 35016 28864
rect 35080 28800 35096 28864
rect 35160 28800 35176 28864
rect 35240 28800 35248 28864
rect 34928 27776 35248 28800
rect 34928 27712 34936 27776
rect 35000 27712 35016 27776
rect 35080 27712 35096 27776
rect 35160 27712 35176 27776
rect 35240 27712 35248 27776
rect 34928 26688 35248 27712
rect 34928 26624 34936 26688
rect 35000 26624 35016 26688
rect 35080 26624 35096 26688
rect 35160 26624 35176 26688
rect 35240 26624 35248 26688
rect 21219 26620 21285 26621
rect 21219 26556 21220 26620
rect 21284 26556 21285 26620
rect 21219 26555 21285 26556
rect 19568 26080 19576 26144
rect 19640 26080 19656 26144
rect 19720 26080 19736 26144
rect 19800 26080 19816 26144
rect 19880 26080 19888 26144
rect 19568 25056 19888 26080
rect 19568 24992 19576 25056
rect 19640 24992 19656 25056
rect 19720 24992 19736 25056
rect 19800 24992 19816 25056
rect 19880 24992 19888 25056
rect 19568 23968 19888 24992
rect 19568 23904 19576 23968
rect 19640 23904 19656 23968
rect 19720 23904 19736 23968
rect 19800 23904 19816 23968
rect 19880 23904 19888 23968
rect 19568 22880 19888 23904
rect 19568 22816 19576 22880
rect 19640 22816 19656 22880
rect 19720 22816 19736 22880
rect 19800 22816 19816 22880
rect 19880 22816 19888 22880
rect 19568 21792 19888 22816
rect 19568 21728 19576 21792
rect 19640 21728 19656 21792
rect 19720 21728 19736 21792
rect 19800 21728 19816 21792
rect 19880 21728 19888 21792
rect 19568 20704 19888 21728
rect 19568 20640 19576 20704
rect 19640 20640 19656 20704
rect 19720 20640 19736 20704
rect 19800 20640 19816 20704
rect 19880 20640 19888 20704
rect 19568 19616 19888 20640
rect 19568 19552 19576 19616
rect 19640 19552 19656 19616
rect 19720 19552 19736 19616
rect 19800 19552 19816 19616
rect 19880 19552 19888 19616
rect 19568 18528 19888 19552
rect 19568 18464 19576 18528
rect 19640 18464 19656 18528
rect 19720 18464 19736 18528
rect 19800 18464 19816 18528
rect 19880 18464 19888 18528
rect 19568 17440 19888 18464
rect 19568 17376 19576 17440
rect 19640 17376 19656 17440
rect 19720 17376 19736 17440
rect 19800 17376 19816 17440
rect 19880 17376 19888 17440
rect 19568 16352 19888 17376
rect 19568 16288 19576 16352
rect 19640 16288 19656 16352
rect 19720 16288 19736 16352
rect 19800 16288 19816 16352
rect 19880 16288 19888 16352
rect 19568 15264 19888 16288
rect 21222 15333 21282 26555
rect 23611 25940 23677 25941
rect 23611 25876 23612 25940
rect 23676 25876 23677 25940
rect 23611 25875 23677 25876
rect 23427 23492 23493 23493
rect 23427 23428 23428 23492
rect 23492 23428 23493 23492
rect 23427 23427 23493 23428
rect 23430 16829 23490 23427
rect 23614 18869 23674 25875
rect 34928 25600 35248 26624
rect 34928 25536 34936 25600
rect 35000 25536 35016 25600
rect 35080 25536 35096 25600
rect 35160 25536 35176 25600
rect 35240 25536 35248 25600
rect 34928 24512 35248 25536
rect 34928 24448 34936 24512
rect 35000 24448 35016 24512
rect 35080 24448 35096 24512
rect 35160 24448 35176 24512
rect 35240 24448 35248 24512
rect 34928 23424 35248 24448
rect 34928 23360 34936 23424
rect 35000 23360 35016 23424
rect 35080 23360 35096 23424
rect 35160 23360 35176 23424
rect 35240 23360 35248 23424
rect 34928 22336 35248 23360
rect 34928 22272 34936 22336
rect 35000 22272 35016 22336
rect 35080 22272 35096 22336
rect 35160 22272 35176 22336
rect 35240 22272 35248 22336
rect 34928 21248 35248 22272
rect 34928 21184 34936 21248
rect 35000 21184 35016 21248
rect 35080 21184 35096 21248
rect 35160 21184 35176 21248
rect 35240 21184 35248 21248
rect 34928 20160 35248 21184
rect 34928 20096 34936 20160
rect 35000 20096 35016 20160
rect 35080 20096 35096 20160
rect 35160 20096 35176 20160
rect 35240 20096 35248 20160
rect 34928 19072 35248 20096
rect 34928 19008 34936 19072
rect 35000 19008 35016 19072
rect 35080 19008 35096 19072
rect 35160 19008 35176 19072
rect 35240 19008 35248 19072
rect 23611 18868 23677 18869
rect 23611 18804 23612 18868
rect 23676 18804 23677 18868
rect 23611 18803 23677 18804
rect 34928 17984 35248 19008
rect 34928 17920 34936 17984
rect 35000 17920 35016 17984
rect 35080 17920 35096 17984
rect 35160 17920 35176 17984
rect 35240 17920 35248 17984
rect 34928 16896 35248 17920
rect 34928 16832 34936 16896
rect 35000 16832 35016 16896
rect 35080 16832 35096 16896
rect 35160 16832 35176 16896
rect 35240 16832 35248 16896
rect 23427 16828 23493 16829
rect 23427 16764 23428 16828
rect 23492 16764 23493 16828
rect 23427 16763 23493 16764
rect 34928 15808 35248 16832
rect 34928 15744 34936 15808
rect 35000 15744 35016 15808
rect 35080 15744 35096 15808
rect 35160 15744 35176 15808
rect 35240 15744 35248 15808
rect 21219 15332 21285 15333
rect 21219 15268 21220 15332
rect 21284 15268 21285 15332
rect 21219 15267 21285 15268
rect 19568 15200 19576 15264
rect 19640 15200 19656 15264
rect 19720 15200 19736 15264
rect 19800 15200 19816 15264
rect 19880 15200 19888 15264
rect 19568 14176 19888 15200
rect 19568 14112 19576 14176
rect 19640 14112 19656 14176
rect 19720 14112 19736 14176
rect 19800 14112 19816 14176
rect 19880 14112 19888 14176
rect 19568 13088 19888 14112
rect 19568 13024 19576 13088
rect 19640 13024 19656 13088
rect 19720 13024 19736 13088
rect 19800 13024 19816 13088
rect 19880 13024 19888 13088
rect 19568 12000 19888 13024
rect 19568 11936 19576 12000
rect 19640 11936 19656 12000
rect 19720 11936 19736 12000
rect 19800 11936 19816 12000
rect 19880 11936 19888 12000
rect 19568 10912 19888 11936
rect 19568 10848 19576 10912
rect 19640 10848 19656 10912
rect 19720 10848 19736 10912
rect 19800 10848 19816 10912
rect 19880 10848 19888 10912
rect 19568 9824 19888 10848
rect 19568 9760 19576 9824
rect 19640 9760 19656 9824
rect 19720 9760 19736 9824
rect 19800 9760 19816 9824
rect 19880 9760 19888 9824
rect 19568 8736 19888 9760
rect 19568 8672 19576 8736
rect 19640 8672 19656 8736
rect 19720 8672 19736 8736
rect 19800 8672 19816 8736
rect 19880 8672 19888 8736
rect 19568 7648 19888 8672
rect 19568 7584 19576 7648
rect 19640 7584 19656 7648
rect 19720 7584 19736 7648
rect 19800 7584 19816 7648
rect 19880 7584 19888 7648
rect 19568 6560 19888 7584
rect 19568 6496 19576 6560
rect 19640 6496 19656 6560
rect 19720 6496 19736 6560
rect 19800 6496 19816 6560
rect 19880 6496 19888 6560
rect 19568 5472 19888 6496
rect 19568 5408 19576 5472
rect 19640 5408 19656 5472
rect 19720 5408 19736 5472
rect 19800 5408 19816 5472
rect 19880 5408 19888 5472
rect 19568 4384 19888 5408
rect 19568 4320 19576 4384
rect 19640 4320 19656 4384
rect 19720 4320 19736 4384
rect 19800 4320 19816 4384
rect 19880 4320 19888 4384
rect 19568 3296 19888 4320
rect 19568 3232 19576 3296
rect 19640 3232 19656 3296
rect 19720 3232 19736 3296
rect 19800 3232 19816 3296
rect 19880 3232 19888 3296
rect 19568 2208 19888 3232
rect 19568 2144 19576 2208
rect 19640 2144 19656 2208
rect 19720 2144 19736 2208
rect 19800 2144 19816 2208
rect 19880 2144 19888 2208
rect 19568 2128 19888 2144
rect 34928 14720 35248 15744
rect 34928 14656 34936 14720
rect 35000 14656 35016 14720
rect 35080 14656 35096 14720
rect 35160 14656 35176 14720
rect 35240 14656 35248 14720
rect 34928 13632 35248 14656
rect 34928 13568 34936 13632
rect 35000 13568 35016 13632
rect 35080 13568 35096 13632
rect 35160 13568 35176 13632
rect 35240 13568 35248 13632
rect 34928 12544 35248 13568
rect 34928 12480 34936 12544
rect 35000 12480 35016 12544
rect 35080 12480 35096 12544
rect 35160 12480 35176 12544
rect 35240 12480 35248 12544
rect 34928 11456 35248 12480
rect 34928 11392 34936 11456
rect 35000 11392 35016 11456
rect 35080 11392 35096 11456
rect 35160 11392 35176 11456
rect 35240 11392 35248 11456
rect 34928 10368 35248 11392
rect 34928 10304 34936 10368
rect 35000 10304 35016 10368
rect 35080 10304 35096 10368
rect 35160 10304 35176 10368
rect 35240 10304 35248 10368
rect 34928 9280 35248 10304
rect 34928 9216 34936 9280
rect 35000 9216 35016 9280
rect 35080 9216 35096 9280
rect 35160 9216 35176 9280
rect 35240 9216 35248 9280
rect 34928 8192 35248 9216
rect 34928 8128 34936 8192
rect 35000 8128 35016 8192
rect 35080 8128 35096 8192
rect 35160 8128 35176 8192
rect 35240 8128 35248 8192
rect 34928 7104 35248 8128
rect 34928 7040 34936 7104
rect 35000 7040 35016 7104
rect 35080 7040 35096 7104
rect 35160 7040 35176 7104
rect 35240 7040 35248 7104
rect 34928 6016 35248 7040
rect 34928 5952 34936 6016
rect 35000 5952 35016 6016
rect 35080 5952 35096 6016
rect 35160 5952 35176 6016
rect 35240 5952 35248 6016
rect 34928 4928 35248 5952
rect 34928 4864 34936 4928
rect 35000 4864 35016 4928
rect 35080 4864 35096 4928
rect 35160 4864 35176 4928
rect 35240 4864 35248 4928
rect 34928 3840 35248 4864
rect 34928 3776 34936 3840
rect 35000 3776 35016 3840
rect 35080 3776 35096 3840
rect 35160 3776 35176 3840
rect 35240 3776 35248 3840
rect 34928 2752 35248 3776
rect 34928 2688 34936 2752
rect 35000 2688 35016 2752
rect 35080 2688 35096 2752
rect 35160 2688 35176 2752
rect 35240 2688 35248 2752
rect 34928 2128 35248 2688
rect 50288 37024 50608 37584
rect 50288 36960 50296 37024
rect 50360 36960 50376 37024
rect 50440 36960 50456 37024
rect 50520 36960 50536 37024
rect 50600 36960 50608 37024
rect 50288 35936 50608 36960
rect 50288 35872 50296 35936
rect 50360 35872 50376 35936
rect 50440 35872 50456 35936
rect 50520 35872 50536 35936
rect 50600 35872 50608 35936
rect 50288 34848 50608 35872
rect 50288 34784 50296 34848
rect 50360 34784 50376 34848
rect 50440 34784 50456 34848
rect 50520 34784 50536 34848
rect 50600 34784 50608 34848
rect 50288 33760 50608 34784
rect 50288 33696 50296 33760
rect 50360 33696 50376 33760
rect 50440 33696 50456 33760
rect 50520 33696 50536 33760
rect 50600 33696 50608 33760
rect 50288 32672 50608 33696
rect 50288 32608 50296 32672
rect 50360 32608 50376 32672
rect 50440 32608 50456 32672
rect 50520 32608 50536 32672
rect 50600 32608 50608 32672
rect 50288 31584 50608 32608
rect 50288 31520 50296 31584
rect 50360 31520 50376 31584
rect 50440 31520 50456 31584
rect 50520 31520 50536 31584
rect 50600 31520 50608 31584
rect 50288 30496 50608 31520
rect 50288 30432 50296 30496
rect 50360 30432 50376 30496
rect 50440 30432 50456 30496
rect 50520 30432 50536 30496
rect 50600 30432 50608 30496
rect 50288 29408 50608 30432
rect 50288 29344 50296 29408
rect 50360 29344 50376 29408
rect 50440 29344 50456 29408
rect 50520 29344 50536 29408
rect 50600 29344 50608 29408
rect 50288 28320 50608 29344
rect 50288 28256 50296 28320
rect 50360 28256 50376 28320
rect 50440 28256 50456 28320
rect 50520 28256 50536 28320
rect 50600 28256 50608 28320
rect 50288 27232 50608 28256
rect 50288 27168 50296 27232
rect 50360 27168 50376 27232
rect 50440 27168 50456 27232
rect 50520 27168 50536 27232
rect 50600 27168 50608 27232
rect 50288 26144 50608 27168
rect 50288 26080 50296 26144
rect 50360 26080 50376 26144
rect 50440 26080 50456 26144
rect 50520 26080 50536 26144
rect 50600 26080 50608 26144
rect 50288 25056 50608 26080
rect 50288 24992 50296 25056
rect 50360 24992 50376 25056
rect 50440 24992 50456 25056
rect 50520 24992 50536 25056
rect 50600 24992 50608 25056
rect 50288 23968 50608 24992
rect 50288 23904 50296 23968
rect 50360 23904 50376 23968
rect 50440 23904 50456 23968
rect 50520 23904 50536 23968
rect 50600 23904 50608 23968
rect 50288 22880 50608 23904
rect 50288 22816 50296 22880
rect 50360 22816 50376 22880
rect 50440 22816 50456 22880
rect 50520 22816 50536 22880
rect 50600 22816 50608 22880
rect 50288 21792 50608 22816
rect 50288 21728 50296 21792
rect 50360 21728 50376 21792
rect 50440 21728 50456 21792
rect 50520 21728 50536 21792
rect 50600 21728 50608 21792
rect 50288 20704 50608 21728
rect 50288 20640 50296 20704
rect 50360 20640 50376 20704
rect 50440 20640 50456 20704
rect 50520 20640 50536 20704
rect 50600 20640 50608 20704
rect 50288 19616 50608 20640
rect 50288 19552 50296 19616
rect 50360 19552 50376 19616
rect 50440 19552 50456 19616
rect 50520 19552 50536 19616
rect 50600 19552 50608 19616
rect 50288 18528 50608 19552
rect 50288 18464 50296 18528
rect 50360 18464 50376 18528
rect 50440 18464 50456 18528
rect 50520 18464 50536 18528
rect 50600 18464 50608 18528
rect 50288 17440 50608 18464
rect 50288 17376 50296 17440
rect 50360 17376 50376 17440
rect 50440 17376 50456 17440
rect 50520 17376 50536 17440
rect 50600 17376 50608 17440
rect 50288 16352 50608 17376
rect 50288 16288 50296 16352
rect 50360 16288 50376 16352
rect 50440 16288 50456 16352
rect 50520 16288 50536 16352
rect 50600 16288 50608 16352
rect 50288 15264 50608 16288
rect 50288 15200 50296 15264
rect 50360 15200 50376 15264
rect 50440 15200 50456 15264
rect 50520 15200 50536 15264
rect 50600 15200 50608 15264
rect 50288 14176 50608 15200
rect 50288 14112 50296 14176
rect 50360 14112 50376 14176
rect 50440 14112 50456 14176
rect 50520 14112 50536 14176
rect 50600 14112 50608 14176
rect 50288 13088 50608 14112
rect 50288 13024 50296 13088
rect 50360 13024 50376 13088
rect 50440 13024 50456 13088
rect 50520 13024 50536 13088
rect 50600 13024 50608 13088
rect 50288 12000 50608 13024
rect 50288 11936 50296 12000
rect 50360 11936 50376 12000
rect 50440 11936 50456 12000
rect 50520 11936 50536 12000
rect 50600 11936 50608 12000
rect 50288 10912 50608 11936
rect 50288 10848 50296 10912
rect 50360 10848 50376 10912
rect 50440 10848 50456 10912
rect 50520 10848 50536 10912
rect 50600 10848 50608 10912
rect 50288 9824 50608 10848
rect 50288 9760 50296 9824
rect 50360 9760 50376 9824
rect 50440 9760 50456 9824
rect 50520 9760 50536 9824
rect 50600 9760 50608 9824
rect 50288 8736 50608 9760
rect 50288 8672 50296 8736
rect 50360 8672 50376 8736
rect 50440 8672 50456 8736
rect 50520 8672 50536 8736
rect 50600 8672 50608 8736
rect 50288 7648 50608 8672
rect 50288 7584 50296 7648
rect 50360 7584 50376 7648
rect 50440 7584 50456 7648
rect 50520 7584 50536 7648
rect 50600 7584 50608 7648
rect 50288 6560 50608 7584
rect 50288 6496 50296 6560
rect 50360 6496 50376 6560
rect 50440 6496 50456 6560
rect 50520 6496 50536 6560
rect 50600 6496 50608 6560
rect 50288 5472 50608 6496
rect 50288 5408 50296 5472
rect 50360 5408 50376 5472
rect 50440 5408 50456 5472
rect 50520 5408 50536 5472
rect 50600 5408 50608 5472
rect 50288 4384 50608 5408
rect 50288 4320 50296 4384
rect 50360 4320 50376 4384
rect 50440 4320 50456 4384
rect 50520 4320 50536 4384
rect 50600 4320 50608 4384
rect 50288 3296 50608 4320
rect 50288 3232 50296 3296
rect 50360 3232 50376 3296
rect 50440 3232 50456 3296
rect 50520 3232 50536 3296
rect 50600 3232 50608 3296
rect 50288 2208 50608 3232
rect 50288 2144 50296 2208
rect 50360 2144 50376 2208
rect 50440 2144 50456 2208
rect 50520 2144 50536 2208
rect 50600 2144 50608 2208
rect 50288 2128 50608 2144
use sky130_fd_sc_hd__diode_2  ANTENNA__1478__B pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 8188 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1479__A
timestamp 1644511149
transform 1 0 8924 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1479__B
timestamp 1644511149
transform 1 0 7084 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1480__A2
timestamp 1644511149
transform 1 0 9016 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1482__A2
timestamp 1644511149
transform 1 0 9384 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1482__B1
timestamp 1644511149
transform -1 0 10120 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1482__B2
timestamp 1644511149
transform 1 0 9476 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1483__A1
timestamp 1644511149
transform -1 0 8648 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1483__A2
timestamp 1644511149
transform 1 0 9016 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1484__A2
timestamp 1644511149
transform 1 0 6992 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1485__A1
timestamp 1644511149
transform 1 0 10028 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1485__A2
timestamp 1644511149
transform 1 0 9752 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1486__A1
timestamp 1644511149
transform 1 0 10304 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1486__A2
timestamp 1644511149
transform 1 0 10856 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1487__B
timestamp 1644511149
transform -1 0 8648 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1488__A
timestamp 1644511149
transform 1 0 9476 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1489__A
timestamp 1644511149
transform 1 0 11224 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1490__A1_N
timestamp 1644511149
transform -1 0 11684 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1491__B
timestamp 1644511149
transform -1 0 17480 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1495__A1
timestamp 1644511149
transform -1 0 14444 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1495__A2
timestamp 1644511149
transform 1 0 14996 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1501__A
timestamp 1644511149
transform 1 0 16652 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1503__B
timestamp 1644511149
transform 1 0 20792 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1506__A
timestamp 1644511149
transform -1 0 20700 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1521__A
timestamp 1644511149
transform 1 0 3772 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1528__A1
timestamp 1644511149
transform -1 0 15456 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1528__A2
timestamp 1644511149
transform 1 0 15548 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1532__A
timestamp 1644511149
transform -1 0 23736 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1533__A0
timestamp 1644511149
transform 1 0 22908 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1533__A1
timestamp 1644511149
transform -1 0 24104 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1534__A
timestamp 1644511149
transform -1 0 26220 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1538__A
timestamp 1644511149
transform 1 0 23736 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1540__A
timestamp 1644511149
transform 1 0 12144 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1556__B2
timestamp 1644511149
transform 1 0 6992 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1560__A1
timestamp 1644511149
transform 1 0 4048 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1565__A
timestamp 1644511149
transform 1 0 21620 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1570__B
timestamp 1644511149
transform -1 0 19320 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1577__A
timestamp 1644511149
transform 1 0 34684 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1577__B
timestamp 1644511149
transform 1 0 33304 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1580__A1
timestamp 1644511149
transform -1 0 29624 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1582__A
timestamp 1644511149
transform -1 0 31648 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1601__A
timestamp 1644511149
transform -1 0 1840 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1603__A1
timestamp 1644511149
transform -1 0 3956 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1611__A
timestamp 1644511149
transform 1 0 24380 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1611__B
timestamp 1644511149
transform 1 0 24472 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1618__A
timestamp 1644511149
transform 1 0 27416 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1621__A
timestamp 1644511149
transform 1 0 32292 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1639__A
timestamp 1644511149
transform 1 0 5244 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1640__A1
timestamp 1644511149
transform 1 0 3036 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1642__A
timestamp 1644511149
transform 1 0 4600 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1643__A1
timestamp 1644511149
transform -1 0 2208 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1643__B2
timestamp 1644511149
transform 1 0 4692 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1649__A1_N
timestamp 1644511149
transform -1 0 24656 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1655__B
timestamp 1644511149
transform -1 0 27140 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1656__A0
timestamp 1644511149
transform 1 0 26312 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1656__A1
timestamp 1644511149
transform 1 0 27508 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1679__A
timestamp 1644511149
transform -1 0 4692 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1682__A1
timestamp 1644511149
transform 1 0 30084 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1686__A
timestamp 1644511149
transform -1 0 39008 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1706__A
timestamp 1644511149
transform 1 0 14536 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1707__A
timestamp 1644511149
transform 1 0 15548 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1711__A1
timestamp 1644511149
transform -1 0 11040 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1715__A1
timestamp 1644511149
transform 1 0 39192 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1717__A1
timestamp 1644511149
transform 1 0 31372 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1730__A
timestamp 1644511149
transform 1 0 18584 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1731__A
timestamp 1644511149
transform -1 0 19872 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1733__B2
timestamp 1644511149
transform 1 0 13340 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1734__A1
timestamp 1644511149
transform 1 0 11776 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1746__A
timestamp 1644511149
transform 1 0 43332 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1752__A2
timestamp 1644511149
transform 1 0 28336 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1752__B1
timestamp 1644511149
transform -1 0 28704 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1754__A
timestamp 1644511149
transform -1 0 5888 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1757__A
timestamp 1644511149
transform 1 0 27416 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1759__A
timestamp 1644511149
transform 1 0 22080 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1762__C
timestamp 1644511149
transform 1 0 27140 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1763__A
timestamp 1644511149
transform 1 0 19872 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1765__A
timestamp 1644511149
transform 1 0 8188 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1767__B
timestamp 1644511149
transform -1 0 25208 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1768__A
timestamp 1644511149
transform -1 0 5244 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1771__A
timestamp 1644511149
transform 1 0 24104 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1780__A
timestamp 1644511149
transform 1 0 8924 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1783__A
timestamp 1644511149
transform 1 0 17940 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1788__A
timestamp 1644511149
transform 1 0 4508 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1791__A
timestamp 1644511149
transform -1 0 26128 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1792__C1
timestamp 1644511149
transform 1 0 22816 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1794__B
timestamp 1644511149
transform -1 0 24564 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1795__A1
timestamp 1644511149
transform -1 0 25116 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1796__A
timestamp 1644511149
transform 1 0 29440 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1797__A
timestamp 1644511149
transform -1 0 26496 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1802__A
timestamp 1644511149
transform -1 0 43976 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1804__A
timestamp 1644511149
transform 1 0 12512 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1811__A
timestamp 1644511149
transform 1 0 20516 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1811__B
timestamp 1644511149
transform 1 0 18584 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1814__A_N
timestamp 1644511149
transform -1 0 10672 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1824__A
timestamp 1644511149
transform 1 0 22448 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1825__A1
timestamp 1644511149
transform -1 0 22264 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1830__A
timestamp 1644511149
transform 1 0 27416 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1834__A
timestamp 1644511149
transform -1 0 3312 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1835__A
timestamp 1644511149
transform -1 0 28796 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1844__A_N
timestamp 1644511149
transform 1 0 17480 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1844__B
timestamp 1644511149
transform 1 0 18032 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1848__A2_N
timestamp 1644511149
transform 1 0 15456 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1849__A
timestamp 1644511149
transform 1 0 4784 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1863__A
timestamp 1644511149
transform 1 0 26956 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1867__A
timestamp 1644511149
transform 1 0 2852 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1871__A
timestamp 1644511149
transform 1 0 37812 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1872__A
timestamp 1644511149
transform -1 0 9200 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1873__A
timestamp 1644511149
transform -1 0 7176 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1873__B
timestamp 1644511149
transform 1 0 7544 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1877__A
timestamp 1644511149
transform 1 0 19228 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1877__B
timestamp 1644511149
transform 1 0 17480 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1880__A1
timestamp 1644511149
transform -1 0 17388 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1880__A2
timestamp 1644511149
transform -1 0 17756 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1880__B1
timestamp 1644511149
transform 1 0 17020 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1882__B
timestamp 1644511149
transform 1 0 14444 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1891__B
timestamp 1644511149
transform 1 0 4692 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1894__A
timestamp 1644511149
transform -1 0 20424 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1903__A
timestamp 1644511149
transform 1 0 28428 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1904__B1
timestamp 1644511149
transform -1 0 27140 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1905__A1
timestamp 1644511149
transform 1 0 27600 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1909__A
timestamp 1644511149
transform -1 0 52164 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1910__A
timestamp 1644511149
transform 1 0 27140 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1913__A
timestamp 1644511149
transform 1 0 9384 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1917__B1
timestamp 1644511149
transform -1 0 8832 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1918__A1
timestamp 1644511149
transform 1 0 10764 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1920__A
timestamp 1644511149
transform 1 0 16468 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1920__B
timestamp 1644511149
transform 1 0 17020 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1924__A
timestamp 1644511149
transform 1 0 13156 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1928__B1
timestamp 1644511149
transform 1 0 15456 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1929__A
timestamp 1644511149
transform -1 0 19964 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1930__A
timestamp 1644511149
transform 1 0 20148 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1931__A
timestamp 1644511149
transform 1 0 33304 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1933__A1
timestamp 1644511149
transform 1 0 22816 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1933__A2
timestamp 1644511149
transform 1 0 21160 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1937__A
timestamp 1644511149
transform -1 0 20792 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1937__B
timestamp 1644511149
transform 1 0 21068 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1941__A
timestamp 1644511149
transform 1 0 5336 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1941__B
timestamp 1644511149
transform 1 0 6532 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1946__A
timestamp 1644511149
transform 1 0 23276 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1955__A
timestamp 1644511149
transform 1 0 30084 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1964__A
timestamp 1644511149
transform -1 0 23460 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1968__A
timestamp 1644511149
transform 1 0 13432 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1968__B
timestamp 1644511149
transform 1 0 12880 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1970__A1
timestamp 1644511149
transform 1 0 15732 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1970__B1
timestamp 1644511149
transform 1 0 15916 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1971__A1
timestamp 1644511149
transform 1 0 16008 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1972__A
timestamp 1644511149
transform 1 0 10764 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1980__A2
timestamp 1644511149
transform 1 0 14076 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1982__A2
timestamp 1644511149
transform 1 0 15180 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1984__A
timestamp 1644511149
transform -1 0 29072 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__1991__A1_N
timestamp 1644511149
transform 1 0 22908 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2005__A1
timestamp 1644511149
transform -1 0 30360 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2011__A
timestamp 1644511149
transform 1 0 29072 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2012__A
timestamp 1644511149
transform 1 0 29624 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2013__A
timestamp 1644511149
transform 1 0 5060 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2018__B
timestamp 1644511149
transform 1 0 30268 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2021__A
timestamp 1644511149
transform -1 0 9752 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2021__B
timestamp 1644511149
transform 1 0 8924 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2027__B1
timestamp 1644511149
transform 1 0 12972 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2028__A
timestamp 1644511149
transform 1 0 30176 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2028__B
timestamp 1644511149
transform -1 0 30544 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2032__A
timestamp 1644511149
transform -1 0 22080 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2032__B
timestamp 1644511149
transform -1 0 22264 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2038__A1
timestamp 1644511149
transform 1 0 18216 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2039__A
timestamp 1644511149
transform 1 0 31372 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2063__A
timestamp 1644511149
transform 1 0 5612 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2065__A
timestamp 1644511149
transform 1 0 22908 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2065__B
timestamp 1644511149
transform 1 0 23092 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2066__A1
timestamp 1644511149
transform 1 0 24564 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2066__B1
timestamp 1644511149
transform 1 0 25116 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2067__A1
timestamp 1644511149
transform -1 0 23828 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2071__A2
timestamp 1644511149
transform 1 0 9476 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2075__B1
timestamp 1644511149
transform 1 0 14076 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2076__A
timestamp 1644511149
transform 1 0 30636 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2078__B
timestamp 1644511149
transform -1 0 30820 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2084__A1
timestamp 1644511149
transform -1 0 22172 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2084__A2
timestamp 1644511149
transform 1 0 20424 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2085__A
timestamp 1644511149
transform 1 0 34868 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2086__A
timestamp 1644511149
transform 1 0 21068 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2086__B
timestamp 1644511149
transform 1 0 20884 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2089__A
timestamp 1644511149
transform -1 0 22816 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2089__B
timestamp 1644511149
transform 1 0 25116 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2093__A
timestamp 1644511149
transform 1 0 23368 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2112__A
timestamp 1644511149
transform 1 0 39008 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2113__A
timestamp 1644511149
transform -1 0 40296 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2124__A
timestamp 1644511149
transform -1 0 26312 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2128__A
timestamp 1644511149
transform 1 0 23736 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2128__B
timestamp 1644511149
transform -1 0 24196 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2129__A
timestamp 1644511149
transform -1 0 26864 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2130__A1
timestamp 1644511149
transform 1 0 25300 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2132__A
timestamp 1644511149
transform 1 0 34040 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2133__B
timestamp 1644511149
transform -1 0 1932 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2134__B
timestamp 1644511149
transform 1 0 2944 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2139__A2
timestamp 1644511149
transform -1 0 12420 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2140__B1
timestamp 1644511149
transform 1 0 12696 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2141__B
timestamp 1644511149
transform -1 0 36800 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2147__A1_N
timestamp 1644511149
transform 1 0 23000 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2150__B
timestamp 1644511149
transform 1 0 20516 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2153__A
timestamp 1644511149
transform 1 0 33488 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2177__A1
timestamp 1644511149
transform -1 0 11684 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2177__A2
timestamp 1644511149
transform -1 0 10396 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2177__B1
timestamp 1644511149
transform -1 0 9568 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2178__A1
timestamp 1644511149
transform -1 0 8464 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2179__A
timestamp 1644511149
transform 1 0 32936 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2179__B
timestamp 1644511149
transform 1 0 33304 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2182__A
timestamp 1644511149
transform 1 0 5152 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2182__B
timestamp 1644511149
transform -1 0 6348 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2188__A2
timestamp 1644511149
transform 1 0 14076 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2190__B
timestamp 1644511149
transform 1 0 35420 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2190__C
timestamp 1644511149
transform -1 0 35788 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2191__A1
timestamp 1644511149
transform -1 0 34224 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2191__A2
timestamp 1644511149
transform -1 0 33672 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2191__B1
timestamp 1644511149
transform -1 0 34500 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2198__B1
timestamp 1644511149
transform 1 0 18492 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2199__A
timestamp 1644511149
transform -1 0 35880 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2199__B
timestamp 1644511149
transform -1 0 34224 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2202__A1
timestamp 1644511149
transform 1 0 19044 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2205__A
timestamp 1644511149
transform 1 0 32660 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2206__A
timestamp 1644511149
transform 1 0 11868 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2206__B
timestamp 1644511149
transform 1 0 10672 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2237__A2
timestamp 1644511149
transform 1 0 36616 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2239__A
timestamp 1644511149
transform 1 0 26956 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2242__A2
timestamp 1644511149
transform 1 0 28888 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2248__A2
timestamp 1644511149
transform -1 0 14812 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2249__A2
timestamp 1644511149
transform 1 0 15640 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2249__B1
timestamp 1644511149
transform -1 0 17204 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2250__B
timestamp 1644511149
transform -1 0 38364 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2254__B1
timestamp 1644511149
transform 1 0 14260 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2255__B
timestamp 1644511149
transform 1 0 33212 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2257__A1
timestamp 1644511149
transform 1 0 17848 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2262__A
timestamp 1644511149
transform 1 0 10856 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2262__B
timestamp 1644511149
transform 1 0 13064 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2264__A
timestamp 1644511149
transform 1 0 10120 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2264__B
timestamp 1644511149
transform -1 0 11868 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2267__A
timestamp 1644511149
transform 1 0 17940 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2269__B
timestamp 1644511149
transform 1 0 39376 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2299__A
timestamp 1644511149
transform -1 0 28980 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2300__A0
timestamp 1644511149
transform 1 0 26312 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2300__A1
timestamp 1644511149
transform -1 0 25944 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2300__S
timestamp 1644511149
transform 1 0 26312 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2303__A
timestamp 1644511149
transform -1 0 27140 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2304__A1
timestamp 1644511149
transform 1 0 28244 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2312__B1
timestamp 1644511149
transform -1 0 13616 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2313__A2
timestamp 1644511149
transform 1 0 30360 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2313__B1
timestamp 1644511149
transform 1 0 30728 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2314__A
timestamp 1644511149
transform 1 0 30544 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2314__C
timestamp 1644511149
transform -1 0 30084 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2321__A
timestamp 1644511149
transform 1 0 19964 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2321__B
timestamp 1644511149
transform 1 0 20976 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2327__B1
timestamp 1644511149
transform 1 0 18584 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2327__B2
timestamp 1644511149
transform 1 0 19228 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2333__B
timestamp 1644511149
transform 1 0 18308 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2335__A1_N
timestamp 1644511149
transform 1 0 18492 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2355__A
timestamp 1644511149
transform 1 0 47840 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2357__A
timestamp 1644511149
transform -1 0 49588 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2362__B
timestamp 1644511149
transform -1 0 7360 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2367__A
timestamp 1644511149
transform 1 0 32844 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2367__B
timestamp 1644511149
transform 1 0 31740 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2367__C
timestamp 1644511149
transform -1 0 34040 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2370__B2
timestamp 1644511149
transform 1 0 28888 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2371__A2
timestamp 1644511149
transform 1 0 26588 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2372__B1
timestamp 1644511149
transform 1 0 32936 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2373__A
timestamp 1644511149
transform -1 0 35236 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2377__A
timestamp 1644511149
transform -1 0 32016 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2389__A1
timestamp 1644511149
transform 1 0 21804 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2395__A
timestamp 1644511149
transform 1 0 25024 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2395__B
timestamp 1644511149
transform 1 0 23736 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2405__A1
timestamp 1644511149
transform -1 0 20608 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2406__B
timestamp 1644511149
transform 1 0 39744 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2415__A
timestamp 1644511149
transform 1 0 5704 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2415__B
timestamp 1644511149
transform 1 0 7452 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2417__A
timestamp 1644511149
transform -1 0 30544 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2417__C
timestamp 1644511149
transform -1 0 29992 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2418__A1
timestamp 1644511149
transform 1 0 30176 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2418__A2
timestamp 1644511149
transform 1 0 29624 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2419__A
timestamp 1644511149
transform -1 0 46460 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2427__A
timestamp 1644511149
transform -1 0 50324 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2428__A
timestamp 1644511149
transform 1 0 48668 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2437__C
timestamp 1644511149
transform 1 0 36800 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2438__A
timestamp 1644511149
transform 1 0 35880 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2446__A
timestamp 1644511149
transform 1 0 11224 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2446__B
timestamp 1644511149
transform 1 0 11776 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2447__A
timestamp 1644511149
transform -1 0 9844 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2452__A
timestamp 1644511149
transform 1 0 27508 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2454__A2
timestamp 1644511149
transform 1 0 28888 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2455__A1
timestamp 1644511149
transform 1 0 29808 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2455__A2
timestamp 1644511149
transform 1 0 29992 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2461__B1
timestamp 1644511149
transform -1 0 25576 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2461__B2
timestamp 1644511149
transform 1 0 22908 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2465__A1
timestamp 1644511149
transform 1 0 21620 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2472__A1
timestamp 1644511149
transform 1 0 20056 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2473__B
timestamp 1644511149
transform -1 0 40388 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2482__B
timestamp 1644511149
transform 1 0 11868 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2484__A1
timestamp 1644511149
transform 1 0 8280 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2485__A1
timestamp 1644511149
transform 1 0 8924 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2486__B
timestamp 1644511149
transform 1 0 13524 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2487__A
timestamp 1644511149
transform 1 0 14720 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2488__B2
timestamp 1644511149
transform -1 0 16836 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2489__B1
timestamp 1644511149
transform -1 0 43424 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2490__C
timestamp 1644511149
transform -1 0 44344 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2494__A
timestamp 1644511149
transform 1 0 49496 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2502__B1
timestamp 1644511149
transform -1 0 54280 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2503__A
timestamp 1644511149
transform -1 0 52256 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2510__A
timestamp 1644511149
transform -1 0 51796 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2518__A
timestamp 1644511149
transform 1 0 27600 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2518__B
timestamp 1644511149
transform 1 0 27232 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2519__A
timestamp 1644511149
transform 1 0 25668 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2519__B
timestamp 1644511149
transform 1 0 26680 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2523__A1
timestamp 1644511149
transform 1 0 12144 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2524__A
timestamp 1644511149
transform 1 0 13064 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2526__A
timestamp 1644511149
transform -1 0 32292 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2529__B
timestamp 1644511149
transform -1 0 42504 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2530__A1
timestamp 1644511149
transform 1 0 41952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2542__B1
timestamp 1644511149
transform 1 0 25852 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2542__B2
timestamp 1644511149
transform 1 0 26220 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2548__A2
timestamp 1644511149
transform 1 0 22448 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2552__A
timestamp 1644511149
transform -1 0 21344 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2557__B
timestamp 1644511149
transform 1 0 40020 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2565__A
timestamp 1644511149
transform 1 0 20976 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2566__A
timestamp 1644511149
transform 1 0 14904 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2566__B
timestamp 1644511149
transform -1 0 15272 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2567__A1_N
timestamp 1644511149
transform -1 0 13616 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2567__B2
timestamp 1644511149
transform 1 0 15272 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2569__B1
timestamp 1644511149
transform 1 0 41768 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2570__C
timestamp 1644511149
transform -1 0 42596 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2585__A
timestamp 1644511149
transform -1 0 53728 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2586__B1
timestamp 1644511149
transform -1 0 52440 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2588__B1
timestamp 1644511149
transform 1 0 50692 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2595__A
timestamp 1644511149
transform 1 0 31464 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2595__B
timestamp 1644511149
transform -1 0 33488 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2595__C
timestamp 1644511149
transform 1 0 31648 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2599__B1
timestamp 1644511149
transform 1 0 38364 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2600__A
timestamp 1644511149
transform -1 0 39100 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2604__A1
timestamp 1644511149
transform 1 0 24196 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2604__A2
timestamp 1644511149
transform -1 0 24932 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2609__A1
timestamp 1644511149
transform 1 0 19044 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2610__B
timestamp 1644511149
transform 1 0 39836 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2614__A
timestamp 1644511149
transform 1 0 32476 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2614__B
timestamp 1644511149
transform -1 0 34776 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2615__A
timestamp 1644511149
transform -1 0 31740 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2615__C
timestamp 1644511149
transform -1 0 31188 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2616__A1
timestamp 1644511149
transform 1 0 31464 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2616__A3
timestamp 1644511149
transform 1 0 30912 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2617__B1
timestamp 1644511149
transform -1 0 31096 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2618__A1
timestamp 1644511149
transform 1 0 34224 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2632__B
timestamp 1644511149
transform 1 0 13432 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2633__A1
timestamp 1644511149
transform -1 0 13708 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2635__B1
timestamp 1644511149
transform -1 0 50324 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2636__C
timestamp 1644511149
transform -1 0 51244 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2664__A1
timestamp 1644511149
transform 1 0 29808 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2664__A2
timestamp 1644511149
transform 1 0 29624 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2668__B1
timestamp 1644511149
transform 1 0 23460 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2675__A1
timestamp 1644511149
transform 1 0 19504 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2676__B
timestamp 1644511149
transform 1 0 40020 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2679__A
timestamp 1644511149
transform -1 0 34132 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2679__C
timestamp 1644511149
transform -1 0 33120 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2681__A1
timestamp 1644511149
transform -1 0 33672 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2681__A2
timestamp 1644511149
transform -1 0 34224 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2682__D1
timestamp 1644511149
transform -1 0 35144 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2692__A1
timestamp 1644511149
transform -1 0 13616 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2694__B1
timestamp 1644511149
transform 1 0 53544 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2695__C
timestamp 1644511149
transform 1 0 52808 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2705__A
timestamp 1644511149
transform 1 0 56120 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2712__A
timestamp 1644511149
transform -1 0 3312 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2723__A
timestamp 1644511149
transform 1 0 14260 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2727__A1
timestamp 1644511149
transform -1 0 37720 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2728__B
timestamp 1644511149
transform 1 0 38456 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2732__B1
timestamp 1644511149
transform 1 0 25116 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2733__A
timestamp 1644511149
transform 1 0 25760 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2741__A1
timestamp 1644511149
transform 1 0 22356 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2742__B
timestamp 1644511149
transform 1 0 40388 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2755__A
timestamp 1644511149
transform 1 0 16284 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2755__B
timestamp 1644511149
transform -1 0 17020 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2758__B
timestamp 1644511149
transform 1 0 50416 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2780__A1
timestamp 1644511149
transform -1 0 56396 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2787__B
timestamp 1644511149
transform -1 0 50416 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2791__B
timestamp 1644511149
transform -1 0 40020 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2793__B1
timestamp 1644511149
transform 1 0 31096 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2799__A
timestamp 1644511149
transform 1 0 31924 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2799__B
timestamp 1644511149
transform -1 0 32292 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2799__C
timestamp 1644511149
transform 1 0 31372 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2808__A
timestamp 1644511149
transform -1 0 19504 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2812__B
timestamp 1644511149
transform 1 0 40296 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2824__A1
timestamp 1644511149
transform -1 0 18216 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2824__A2
timestamp 1644511149
transform 1 0 18400 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2826__B
timestamp 1644511149
transform -1 0 48116 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2835__A
timestamp 1644511149
transform 1 0 55384 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2836__A1
timestamp 1644511149
transform 1 0 57040 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2838__B
timestamp 1644511149
transform -1 0 56396 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2840__B1
timestamp 1644511149
transform 1 0 47656 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2846__A1
timestamp 1644511149
transform 1 0 21804 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2848__A
timestamp 1644511149
transform -1 0 13800 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2851__A1
timestamp 1644511149
transform 1 0 30636 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2851__A2
timestamp 1644511149
transform 1 0 30820 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2852__A
timestamp 1644511149
transform 1 0 32016 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2856__A1
timestamp 1644511149
transform -1 0 28704 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2857__A
timestamp 1644511149
transform 1 0 33212 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2863__A1
timestamp 1644511149
transform -1 0 15180 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2865__B1
timestamp 1644511149
transform 1 0 42412 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2866__C
timestamp 1644511149
transform -1 0 42964 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2882__A
timestamp 1644511149
transform 1 0 53176 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2883__A
timestamp 1644511149
transform -1 0 55936 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2884__A2
timestamp 1644511149
transform 1 0 57224 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2896__A1
timestamp 1644511149
transform -1 0 15548 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2898__B1_N
timestamp 1644511149
transform -1 0 35512 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2899__C_N
timestamp 1644511149
transform 1 0 35604 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2900__A_N
timestamp 1644511149
transform -1 0 36432 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2907__A1
timestamp 1644511149
transform 1 0 23092 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2908__A
timestamp 1644511149
transform 1 0 13340 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2909__A
timestamp 1644511149
transform 1 0 13432 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2910__A0
timestamp 1644511149
transform -1 0 14352 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2910__A1
timestamp 1644511149
transform -1 0 11868 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2918__A2
timestamp 1644511149
transform 1 0 18584 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2919__A
timestamp 1644511149
transform 1 0 15824 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2921__B
timestamp 1644511149
transform -1 0 39836 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2930__A_N
timestamp 1644511149
transform -1 0 10304 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2930__B
timestamp 1644511149
transform 1 0 10672 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2931__A
timestamp 1644511149
transform 1 0 11500 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2932__B
timestamp 1644511149
transform -1 0 9936 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2933__B
timestamp 1644511149
transform -1 0 7820 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2935__A
timestamp 1644511149
transform 1 0 53544 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2936__B2
timestamp 1644511149
transform 1 0 54556 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2938__A2
timestamp 1644511149
transform -1 0 57960 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2939__B
timestamp 1644511149
transform 1 0 6348 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2943__A
timestamp 1644511149
transform 1 0 14444 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2943__B
timestamp 1644511149
transform 1 0 14812 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2950__A
timestamp 1644511149
transform 1 0 18308 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2956__B
timestamp 1644511149
transform 1 0 17572 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2957__A
timestamp 1644511149
transform 1 0 19596 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2957__B
timestamp 1644511149
transform -1 0 18952 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2963__A
timestamp 1644511149
transform 1 0 15732 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2966__A
timestamp 1644511149
transform -1 0 12236 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2966__B
timestamp 1644511149
transform 1 0 11684 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2969__A
timestamp 1644511149
transform -1 0 38824 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2971__A3
timestamp 1644511149
transform 1 0 38824 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2972__B
timestamp 1644511149
transform -1 0 10120 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2973__A
timestamp 1644511149
transform -1 0 10120 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2975__B
timestamp 1644511149
transform 1 0 10580 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2976__B
timestamp 1644511149
transform -1 0 9752 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2978__A
timestamp 1644511149
transform -1 0 8004 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2979__A
timestamp 1644511149
transform -1 0 7912 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA__2981__B
timestamp 1644511149
transform -1 0 53636 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input1_A
timestamp 1644511149
transform -1 0 1748 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input2_A
timestamp 1644511149
transform -1 0 57408 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input3_A
timestamp 1644511149
transform -1 0 57500 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input4_A
timestamp 1644511149
transform -1 0 58236 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input5_A
timestamp 1644511149
transform -1 0 41952 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input6_A
timestamp 1644511149
transform -1 0 28060 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input7_A
timestamp 1644511149
transform -1 0 29992 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input8_A
timestamp 1644511149
transform -1 0 1564 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input9_A
timestamp 1644511149
transform -1 0 56856 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input10_A
timestamp 1644511149
transform -1 0 57408 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input11_A
timestamp 1644511149
transform -1 0 58236 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input12_A
timestamp 1644511149
transform -1 0 25484 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input13_A
timestamp 1644511149
transform -1 0 35788 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input14_A
timestamp 1644511149
transform -1 0 1564 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input15_A
timestamp 1644511149
transform -1 0 7452 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input16_A
timestamp 1644511149
transform -1 0 58236 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input17_A
timestamp 1644511149
transform -1 0 23920 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input18_A
timestamp 1644511149
transform -1 0 1748 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input19_A
timestamp 1644511149
transform -1 0 1748 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input20_A
timestamp 1644511149
transform -1 0 58236 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input21_A
timestamp 1644511149
transform -1 0 9384 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input22_A
timestamp 1644511149
transform -1 0 58236 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input23_A
timestamp 1644511149
transform -1 0 58236 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input24_A
timestamp 1644511149
transform -1 0 1748 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input25_A
timestamp 1644511149
transform -1 0 19596 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input26_A
timestamp 1644511149
transform -1 0 58236 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input27_A
timestamp 1644511149
transform -1 0 32292 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input28_A
timestamp 1644511149
transform -1 0 56672 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input29_A
timestamp 1644511149
transform -1 0 58236 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input30_A
timestamp 1644511149
transform -1 0 43424 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input31_A
timestamp 1644511149
transform -1 0 33580 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input32_A
timestamp 1644511149
transform -1 0 9384 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input33_A
timestamp 1644511149
transform 1 0 58052 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input34_A
timestamp 1644511149
transform -1 0 19688 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input35_A
timestamp 1644511149
transform -1 0 1748 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input36_A
timestamp 1644511149
transform -1 0 23184 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input37_A
timestamp 1644511149
transform -1 0 2484 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input38_A
timestamp 1644511149
transform -1 0 29072 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input39_A
timestamp 1644511149
transform -1 0 1564 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input40_A
timestamp 1644511149
transform -1 0 37628 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input41_A
timestamp 1644511149
transform -1 0 1748 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input42_A
timestamp 1644511149
transform -1 0 11960 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input43_A
timestamp 1644511149
transform -1 0 1748 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input44_A
timestamp 1644511149
transform -1 0 3036 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input45_A
timestamp 1644511149
transform -1 0 55752 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input46_A
timestamp 1644511149
transform -1 0 48576 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input47_A
timestamp 1644511149
transform -1 0 21988 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input48_A
timestamp 1644511149
transform -1 0 58236 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input49_A
timestamp 1644511149
transform -1 0 55476 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input50_A
timestamp 1644511149
transform -1 0 1564 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input51_A
timestamp 1644511149
transform -1 0 1564 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input52_A
timestamp 1644511149
transform -1 0 8648 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input53_A
timestamp 1644511149
transform -1 0 16836 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input54_A
timestamp 1644511149
transform -1 0 27048 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input55_A
timestamp 1644511149
transform -1 0 58236 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input56_A
timestamp 1644511149
transform -1 0 27784 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input57_A
timestamp 1644511149
transform -1 0 50508 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input58_A
timestamp 1644511149
transform -1 0 49128 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input59_A
timestamp 1644511149
transform -1 0 14260 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input60_A
timestamp 1644511149
transform -1 0 23092 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input61_A
timestamp 1644511149
transform -1 0 34224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input62_A
timestamp 1644511149
transform -1 0 2208 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input63_A
timestamp 1644511149
transform -1 0 4140 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_input64_A
timestamp 1644511149
transform -1 0 58236 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output65_A
timestamp 1644511149
transform -1 0 52256 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output66_A
timestamp 1644511149
transform 1 0 12420 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output67_A
timestamp 1644511149
transform 1 0 51060 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output68_A
timestamp 1644511149
transform 1 0 46552 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output72_A
timestamp 1644511149
transform 1 0 48484 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output75_A
timestamp 1644511149
transform 1 0 40940 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output76_A
timestamp 1644511149
transform -1 0 17756 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output82_A
timestamp 1644511149
transform 1 0 37536 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output83_A
timestamp 1644511149
transform -1 0 3036 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output84_A
timestamp 1644511149
transform -1 0 16192 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output88_A
timestamp 1644511149
transform 1 0 57684 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output89_A
timestamp 1644511149
transform -1 0 57316 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output90_A
timestamp 1644511149
transform -1 0 2300 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output94_A
timestamp 1644511149
transform -1 0 57868 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output95_A
timestamp 1644511149
transform 1 0 2116 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_output96_A
timestamp 1644511149
transform 1 0 41492 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12 pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2208 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20 pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 2944 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29 pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3772 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_35 pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 4324 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47
timestamp 1644511149
transform 1 0 5428 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55 pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6164 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_57
timestamp 1644511149
transform 1 0 6348 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69
timestamp 1644511149
transform 1 0 7452 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_80
timestamp 1644511149
transform 1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_85 pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8924 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_90
timestamp 1644511149
transform 1 0 9384 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_104
timestamp 1644511149
transform 1 0 10672 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_113
timestamp 1644511149
transform 1 0 11500 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_119
timestamp 1644511149
transform 1 0 12052 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_125
timestamp 1644511149
transform 1 0 12604 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_137
timestamp 1644511149
transform 1 0 13708 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_145
timestamp 1644511149
transform 1 0 14444 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_153
timestamp 1644511149
transform 1 0 15180 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_164
timestamp 1644511149
transform 1 0 16192 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_171
timestamp 1644511149
transform 1 0 16836 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_181
timestamp 1644511149
transform 1 0 17756 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_189 pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 18492 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_195
timestamp 1644511149
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_197
timestamp 1644511149
transform 1 0 19228 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_201
timestamp 1644511149
transform 1 0 19596 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_209
timestamp 1644511149
transform 1 0 20332 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_218
timestamp 1644511149
transform 1 0 21160 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_225
timestamp 1644511149
transform 1 0 21804 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_231
timestamp 1644511149
transform 1 0 22356 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_237
timestamp 1644511149
transform 1 0 22908 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_240
timestamp 1644511149
transform 1 0 23184 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_247
timestamp 1644511149
transform 1 0 23828 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_251
timestamp 1644511149
transform 1 0 24196 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_253
timestamp 1644511149
transform 1 0 24380 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_263
timestamp 1644511149
transform 1 0 25300 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_276
timestamp 1644511149
transform 1 0 26496 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_285
timestamp 1644511149
transform 1 0 27324 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_289
timestamp 1644511149
transform 1 0 27692 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_296
timestamp 1644511149
transform 1 0 28336 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_304
timestamp 1644511149
transform 1 0 29072 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_309
timestamp 1644511149
transform 1 0 29532 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_319
timestamp 1644511149
transform 1 0 30452 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_327
timestamp 1644511149
transform 1 0 31188 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_332
timestamp 1644511149
transform 1 0 31648 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_337
timestamp 1644511149
transform 1 0 32108 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_343
timestamp 1644511149
transform 1 0 32660 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_352
timestamp 1644511149
transform 1 0 33488 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_360
timestamp 1644511149
transform 1 0 34224 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_371
timestamp 1644511149
transform 1 0 35236 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_377
timestamp 1644511149
transform 1 0 35788 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_385
timestamp 1644511149
transform 1 0 36524 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_391
timestamp 1644511149
transform 1 0 37076 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_393
timestamp 1644511149
transform 1 0 37260 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_398
timestamp 1644511149
transform 1 0 37720 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_406
timestamp 1644511149
transform 1 0 38456 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_418
timestamp 1644511149
transform 1 0 39560 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_421
timestamp 1644511149
transform 1 0 39836 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_427
timestamp 1644511149
transform 1 0 40388 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_435
timestamp 1644511149
transform 1 0 41124 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_441
timestamp 1644511149
transform 1 0 41676 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_444
timestamp 1644511149
transform 1 0 41952 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_455
timestamp 1644511149
transform 1 0 42964 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_461
timestamp 1644511149
transform 1 0 43516 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_469
timestamp 1644511149
transform 1 0 44252 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_475
timestamp 1644511149
transform 1 0 44804 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_477
timestamp 1644511149
transform 1 0 44988 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_485
timestamp 1644511149
transform 1 0 45724 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_490
timestamp 1644511149
transform 1 0 46184 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_496
timestamp 1644511149
transform 1 0 46736 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_505
timestamp 1644511149
transform 1 0 47564 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_511
timestamp 1644511149
transform 1 0 48116 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_517
timestamp 1644511149
transform 1 0 48668 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_529
timestamp 1644511149
transform 1 0 49772 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_533
timestamp 1644511149
transform 1 0 50140 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_539
timestamp 1644511149
transform 1 0 50692 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_0_545
timestamp 1644511149
transform 1 0 51244 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_557
timestamp 1644511149
transform 1 0 52348 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_565
timestamp 1644511149
transform 1 0 53084 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_573
timestamp 1644511149
transform 1 0 53820 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_584
timestamp 1644511149
transform 1 0 54832 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_591
timestamp 1644511149
transform 1 0 55476 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_595
timestamp 1644511149
transform 1 0 55844 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_602
timestamp 1644511149
transform 1 0 56488 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_612
timestamp 1644511149
transform 1 0 57408 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_621
timestamp 1644511149
transform 1 0 58236 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_9
timestamp 1644511149
transform 1 0 1932 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_15
timestamp 1644511149
transform 1 0 2484 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_21
timestamp 1644511149
transform 1 0 3036 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_33
timestamp 1644511149
transform 1 0 4140 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_39
timestamp 1644511149
transform 1 0 4692 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_50
timestamp 1644511149
transform 1 0 5704 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_57
timestamp 1644511149
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_69
timestamp 1644511149
transform 1 0 7452 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_1_77
timestamp 1644511149
transform 1 0 8188 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_1_82
timestamp 1644511149
transform 1 0 8648 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_88
timestamp 1644511149
transform 1 0 9200 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_102
timestamp 1644511149
transform 1 0 10488 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_108
timestamp 1644511149
transform 1 0 11040 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_121
timestamp 1644511149
transform 1 0 12236 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_127
timestamp 1644511149
transform 1 0 12788 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_135
timestamp 1644511149
transform 1 0 13524 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_144
timestamp 1644511149
transform 1 0 14352 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_156
timestamp 1644511149
transform 1 0 15456 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_176
timestamp 1644511149
transform 1 0 17296 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_183
timestamp 1644511149
transform 1 0 17940 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_198
timestamp 1644511149
transform 1 0 19320 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_204
timestamp 1644511149
transform 1 0 19872 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_1_218
timestamp 1644511149
transform 1 0 21160 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_1_227
timestamp 1644511149
transform 1 0 21988 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_239
timestamp 1644511149
transform 1 0 23092 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_248
timestamp 1644511149
transform 1 0 23920 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_257
timestamp 1644511149
transform 1 0 24748 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_261
timestamp 1644511149
transform 1 0 25116 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_265
timestamp 1644511149
transform 1 0 25484 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_276
timestamp 1644511149
transform 1 0 26496 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_284
timestamp 1644511149
transform 1 0 27232 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_301
timestamp 1644511149
transform 1 0 28796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_1_327
timestamp 1644511149
transform 1 0 31188 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_1_335
timestamp 1644511149
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_339
timestamp 1644511149
transform 1 0 32292 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_352
timestamp 1644511149
transform 1 0 33488 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_361
timestamp 1644511149
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_373
timestamp 1644511149
transform 1 0 35420 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_388
timestamp 1644511149
transform 1 0 36800 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_400
timestamp 1644511149
transform 1 0 37904 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_1_412
timestamp 1644511149
transform 1 0 39008 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_1_426
timestamp 1644511149
transform 1 0 40296 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_435
timestamp 1644511149
transform 1 0 41124 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_439
timestamp 1644511149
transform 1 0 41492 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_444
timestamp 1644511149
transform 1 0 41952 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_454
timestamp 1644511149
transform 1 0 42872 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_460
timestamp 1644511149
transform 1 0 43424 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_468
timestamp 1644511149
transform 1 0 44160 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_1_485
timestamp 1644511149
transform 1 0 45724 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_1_497
timestamp 1644511149
transform 1 0 46828 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_1_503
timestamp 1644511149
transform 1 0 47380 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_505
timestamp 1644511149
transform 1 0 47564 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_517
timestamp 1644511149
transform 1 0 48668 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_529
timestamp 1644511149
transform 1 0 49772 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_541
timestamp 1644511149
transform 1 0 50876 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_545
timestamp 1644511149
transform 1 0 51244 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_549
timestamp 1644511149
transform 1 0 51612 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_555
timestamp 1644511149
transform 1 0 52164 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_559
timestamp 1644511149
transform 1 0 52532 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_1_561
timestamp 1644511149
transform 1 0 52716 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_573
timestamp 1644511149
transform 1 0 53820 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_585
timestamp 1644511149
transform 1 0 54924 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_597
timestamp 1644511149
transform 1 0 56028 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_601
timestamp 1644511149
transform 1 0 56396 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_1_604
timestamp 1644511149
transform 1 0 56672 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_612
timestamp 1644511149
transform 1 0 57408 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_621
timestamp 1644511149
transform 1 0 58236 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_5
timestamp 1644511149
transform 1 0 1564 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_17
timestamp 1644511149
transform 1 0 2668 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_25
timestamp 1644511149
transform 1 0 3404 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_2_29
timestamp 1644511149
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_41
timestamp 1644511149
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_53
timestamp 1644511149
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_65
timestamp 1644511149
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_77
timestamp 1644511149
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_83
timestamp 1644511149
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_85
timestamp 1644511149
transform 1 0 8924 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_98
timestamp 1644511149
transform 1 0 10120 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_102
timestamp 1644511149
transform 1 0 10488 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_106
timestamp 1644511149
transform 1 0 10856 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_113
timestamp 1644511149
transform 1 0 11500 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_132
timestamp 1644511149
transform 1 0 13248 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_146
timestamp 1644511149
transform 1 0 14536 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_153
timestamp 1644511149
transform 1 0 15180 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_159
timestamp 1644511149
transform 1 0 15732 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_167
timestamp 1644511149
transform 1 0 16468 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_2_172
timestamp 1644511149
transform 1 0 16928 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_184
timestamp 1644511149
transform 1 0 18032 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_192
timestamp 1644511149
transform 1 0 18768 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_200
timestamp 1644511149
transform 1 0 19504 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_209
timestamp 1644511149
transform 1 0 20332 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_2_217
timestamp 1644511149
transform 1 0 21068 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_240
timestamp 1644511149
transform 1 0 23184 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_258
timestamp 1644511149
transform 1 0 24840 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_276
timestamp 1644511149
transform 1 0 26496 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_282
timestamp 1644511149
transform 1 0 27048 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_2_290
timestamp 1644511149
transform 1 0 27784 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_296
timestamp 1644511149
transform 1 0 28336 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_304
timestamp 1644511149
transform 1 0 29072 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_309
timestamp 1644511149
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_321
timestamp 1644511149
transform 1 0 30636 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_327
timestamp 1644511149
transform 1 0 31188 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_331
timestamp 1644511149
transform 1 0 31556 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_340
timestamp 1644511149
transform 1 0 32384 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_347
timestamp 1644511149
transform 1 0 33028 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_351
timestamp 1644511149
transform 1 0 33396 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_357
timestamp 1644511149
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_363
timestamp 1644511149
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_365
timestamp 1644511149
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_377
timestamp 1644511149
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_2_389
timestamp 1644511149
transform 1 0 36892 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_2_398
timestamp 1644511149
transform 1 0 37720 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_410
timestamp 1644511149
transform 1 0 38824 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_418
timestamp 1644511149
transform 1 0 39560 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_421
timestamp 1644511149
transform 1 0 39836 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_2_426
timestamp 1644511149
transform 1 0 40296 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_2_435
timestamp 1644511149
transform 1 0 41124 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_441
timestamp 1644511149
transform 1 0 41676 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_2_450
timestamp 1644511149
transform 1 0 42504 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_456
timestamp 1644511149
transform 1 0 43056 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_460
timestamp 1644511149
transform 1 0 43424 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_2_466
timestamp 1644511149
transform 1 0 43976 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_2_474
timestamp 1644511149
transform 1 0 44712 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_2_477
timestamp 1644511149
transform 1 0 44988 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_2_492
timestamp 1644511149
transform 1 0 46368 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_504
timestamp 1644511149
transform 1 0 47472 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_516
timestamp 1644511149
transform 1 0 48576 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_2_528
timestamp 1644511149
transform 1 0 49680 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_2_533
timestamp 1644511149
transform 1 0 50140 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_545
timestamp 1644511149
transform 1 0 51244 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_557
timestamp 1644511149
transform 1 0 52348 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_2_569
timestamp 1644511149
transform 1 0 53452 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_2_581
timestamp 1644511149
transform 1 0 54556 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_587
timestamp 1644511149
transform 1 0 55108 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_2_589
timestamp 1644511149
transform 1 0 55292 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_2_601
timestamp 1644511149
transform 1 0 56396 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_2_611
timestamp 1644511149
transform 1 0 57316 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_2_621
timestamp 1644511149
transform 1 0 58236 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1644511149
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_15
timestamp 1644511149
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_27
timestamp 1644511149
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_39
timestamp 1644511149
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_51
timestamp 1644511149
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_55
timestamp 1644511149
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_62
timestamp 1644511149
transform 1 0 6808 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_74
timestamp 1644511149
transform 1 0 7912 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_86
timestamp 1644511149
transform 1 0 9016 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_103
timestamp 1644511149
transform 1 0 10580 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_3_111
timestamp 1644511149
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_3_113
timestamp 1644511149
transform 1 0 11500 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_118
timestamp 1644511149
transform 1 0 11960 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_3_129
timestamp 1644511149
transform 1 0 12972 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_135
timestamp 1644511149
transform 1 0 13524 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_3_143
timestamp 1644511149
transform 1 0 14260 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_148
timestamp 1644511149
transform 1 0 14720 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_160
timestamp 1644511149
transform 1 0 15824 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_164
timestamp 1644511149
transform 1 0 16192 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_174
timestamp 1644511149
transform 1 0 17112 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_186
timestamp 1644511149
transform 1 0 18216 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_198
timestamp 1644511149
transform 1 0 19320 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_210
timestamp 1644511149
transform 1 0 20424 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_3_216
timestamp 1644511149
transform 1 0 20976 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_3_225
timestamp 1644511149
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_237
timestamp 1644511149
transform 1 0 22908 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_3_250
timestamp 1644511149
transform 1 0 24104 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_262
timestamp 1644511149
transform 1 0 25208 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_274
timestamp 1644511149
transform 1 0 26312 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_3_281
timestamp 1644511149
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_293
timestamp 1644511149
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_305
timestamp 1644511149
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_317
timestamp 1644511149
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_329
timestamp 1644511149
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_335
timestamp 1644511149
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_337
timestamp 1644511149
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_349
timestamp 1644511149
transform 1 0 33212 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_355
timestamp 1644511149
transform 1 0 33764 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_367
timestamp 1644511149
transform 1 0 34868 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_379
timestamp 1644511149
transform 1 0 35972 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_3_387
timestamp 1644511149
transform 1 0 36708 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_3_391
timestamp 1644511149
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_400
timestamp 1644511149
transform 1 0 37904 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_412
timestamp 1644511149
transform 1 0 39008 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_3_424
timestamp 1644511149
transform 1 0 40112 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_433
timestamp 1644511149
transform 1 0 40940 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_3_440
timestamp 1644511149
transform 1 0 41584 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_3_449
timestamp 1644511149
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_461
timestamp 1644511149
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_3_473
timestamp 1644511149
transform 1 0 44620 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_3_481
timestamp 1644511149
transform 1 0 45356 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_3_494
timestamp 1644511149
transform 1 0 46552 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_502
timestamp 1644511149
transform 1 0 47288 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_3_505
timestamp 1644511149
transform 1 0 47564 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_517
timestamp 1644511149
transform 1 0 48668 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_529
timestamp 1644511149
transform 1 0 49772 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_541
timestamp 1644511149
transform 1 0 50876 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_553
timestamp 1644511149
transform 1 0 51980 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_559
timestamp 1644511149
transform 1 0 52532 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_561
timestamp 1644511149
transform 1 0 52716 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_573
timestamp 1644511149
transform 1 0 53820 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_585
timestamp 1644511149
transform 1 0 54924 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_597
timestamp 1644511149
transform 1 0 56028 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_3_609
timestamp 1644511149
transform 1 0 57132 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_3_615
timestamp 1644511149
transform 1 0 57684 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_3_617
timestamp 1644511149
transform 1 0 57868 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_3_621
timestamp 1644511149
transform 1 0 58236 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_7
timestamp 1644511149
transform 1 0 1748 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_11
timestamp 1644511149
transform 1 0 2116 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_15
timestamp 1644511149
transform 1 0 2484 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_21
timestamp 1644511149
transform 1 0 3036 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_27
timestamp 1644511149
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_32
timestamp 1644511149
transform 1 0 4048 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_44
timestamp 1644511149
transform 1 0 5152 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_62
timestamp 1644511149
transform 1 0 6808 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_69
timestamp 1644511149
transform 1 0 7452 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_4_81
timestamp 1644511149
transform 1 0 8556 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_85
timestamp 1644511149
transform 1 0 8924 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_89
timestamp 1644511149
transform 1 0 9292 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_111
timestamp 1644511149
transform 1 0 11316 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_123
timestamp 1644511149
transform 1 0 12420 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_4_135
timestamp 1644511149
transform 1 0 13524 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_139
timestamp 1644511149
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_141
timestamp 1644511149
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_153
timestamp 1644511149
transform 1 0 15180 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_161
timestamp 1644511149
transform 1 0 15916 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_165
timestamp 1644511149
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_177
timestamp 1644511149
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_189
timestamp 1644511149
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_195
timestamp 1644511149
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_197
timestamp 1644511149
transform 1 0 19228 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_204
timestamp 1644511149
transform 1 0 19872 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_216
timestamp 1644511149
transform 1 0 20976 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_228
timestamp 1644511149
transform 1 0 22080 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_240
timestamp 1644511149
transform 1 0 23184 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_258
timestamp 1644511149
transform 1 0 24840 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_270
timestamp 1644511149
transform 1 0 25944 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_278
timestamp 1644511149
transform 1 0 26680 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_288
timestamp 1644511149
transform 1 0 27600 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_300
timestamp 1644511149
transform 1 0 28704 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_309
timestamp 1644511149
transform 1 0 29532 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_324
timestamp 1644511149
transform 1 0 30912 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_336
timestamp 1644511149
transform 1 0 32016 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_344
timestamp 1644511149
transform 1 0 32752 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_355
timestamp 1644511149
transform 1 0 33764 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_363
timestamp 1644511149
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_365
timestamp 1644511149
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_377
timestamp 1644511149
transform 1 0 35788 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_385
timestamp 1644511149
transform 1 0 36524 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_4_392
timestamp 1644511149
transform 1 0 37168 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_396
timestamp 1644511149
transform 1 0 37536 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_400
timestamp 1644511149
transform 1 0 37904 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_412
timestamp 1644511149
transform 1 0 39008 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_421
timestamp 1644511149
transform 1 0 39836 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_432
timestamp 1644511149
transform 1 0 40848 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_4_441
timestamp 1644511149
transform 1 0 41676 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_453
timestamp 1644511149
transform 1 0 42780 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_465
timestamp 1644511149
transform 1 0 43884 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_473
timestamp 1644511149
transform 1 0 44620 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_480
timestamp 1644511149
transform 1 0 45264 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_488
timestamp 1644511149
transform 1 0 46000 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_4_497
timestamp 1644511149
transform 1 0 46828 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_509
timestamp 1644511149
transform 1 0 47932 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_4_521
timestamp 1644511149
transform 1 0 49036 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_529
timestamp 1644511149
transform 1 0 49772 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_4_533
timestamp 1644511149
transform 1 0 50140 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_545
timestamp 1644511149
transform 1 0 51244 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_557
timestamp 1644511149
transform 1 0 52348 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_569
timestamp 1644511149
transform 1 0 53452 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_4_581
timestamp 1644511149
transform 1 0 54556 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_4_587
timestamp 1644511149
transform 1 0 55108 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_4_589
timestamp 1644511149
transform 1 0 55292 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_601
timestamp 1644511149
transform 1 0 56396 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_4_613
timestamp 1644511149
transform 1 0 57500 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_3
timestamp 1644511149
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_15
timestamp 1644511149
transform 1 0 2484 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_24
timestamp 1644511149
transform 1 0 3312 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_37
timestamp 1644511149
transform 1 0 4508 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_49
timestamp 1644511149
transform 1 0 5612 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_55
timestamp 1644511149
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_63
timestamp 1644511149
transform 1 0 6900 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_75
timestamp 1644511149
transform 1 0 8004 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_5_87
timestamp 1644511149
transform 1 0 9108 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_92
timestamp 1644511149
transform 1 0 9568 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_104
timestamp 1644511149
transform 1 0 10672 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_113
timestamp 1644511149
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_125
timestamp 1644511149
transform 1 0 12604 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_131
timestamp 1644511149
transform 1 0 13156 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_137
timestamp 1644511149
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_149
timestamp 1644511149
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_161
timestamp 1644511149
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_167
timestamp 1644511149
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_175
timestamp 1644511149
transform 1 0 17204 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_183
timestamp 1644511149
transform 1 0 17940 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_195
timestamp 1644511149
transform 1 0 19044 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_201
timestamp 1644511149
transform 1 0 19596 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_207
timestamp 1644511149
transform 1 0 20148 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_219
timestamp 1644511149
transform 1 0 21252 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_223
timestamp 1644511149
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_225
timestamp 1644511149
transform 1 0 21804 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_5_240
timestamp 1644511149
transform 1 0 23184 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_5_254
timestamp 1644511149
transform 1 0 24472 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_265
timestamp 1644511149
transform 1 0 25484 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_277
timestamp 1644511149
transform 1 0 26588 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_281
timestamp 1644511149
transform 1 0 26956 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_292
timestamp 1644511149
transform 1 0 27968 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_304
timestamp 1644511149
transform 1 0 29072 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_316
timestamp 1644511149
transform 1 0 30176 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_324
timestamp 1644511149
transform 1 0 30912 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_332
timestamp 1644511149
transform 1 0 31648 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_337
timestamp 1644511149
transform 1 0 32108 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_358
timestamp 1644511149
transform 1 0 34040 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_370
timestamp 1644511149
transform 1 0 35144 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_382
timestamp 1644511149
transform 1 0 36248 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_5_390
timestamp 1644511149
transform 1 0 36984 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_5_393
timestamp 1644511149
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_405
timestamp 1644511149
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_417
timestamp 1644511149
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_429
timestamp 1644511149
transform 1 0 40572 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_433
timestamp 1644511149
transform 1 0 40940 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_445
timestamp 1644511149
transform 1 0 42044 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_449
timestamp 1644511149
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_461
timestamp 1644511149
transform 1 0 43516 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_5_465
timestamp 1644511149
transform 1 0 43884 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_473
timestamp 1644511149
transform 1 0 44620 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_5_484
timestamp 1644511149
transform 1 0 45632 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_496
timestamp 1644511149
transform 1 0 46736 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_505
timestamp 1644511149
transform 1 0 47564 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_517
timestamp 1644511149
transform 1 0 48668 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_529
timestamp 1644511149
transform 1 0 49772 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_5_541
timestamp 1644511149
transform 1 0 50876 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_5_553
timestamp 1644511149
transform 1 0 51980 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_559
timestamp 1644511149
transform 1 0 52532 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_561
timestamp 1644511149
transform 1 0 52716 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_5_573
timestamp 1644511149
transform 1 0 53820 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_5_583
timestamp 1644511149
transform 1 0 54740 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_5_595
timestamp 1644511149
transform 1 0 55844 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_601
timestamp 1644511149
transform 1 0 56396 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_612
timestamp 1644511149
transform 1 0 57408 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_5_617
timestamp 1644511149
transform 1 0 57868 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_3
timestamp 1644511149
transform 1 0 1380 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_7
timestamp 1644511149
transform 1 0 1748 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_19
timestamp 1644511149
transform 1 0 2852 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_27
timestamp 1644511149
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_29
timestamp 1644511149
transform 1 0 3772 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_33
timestamp 1644511149
transform 1 0 4140 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_47
timestamp 1644511149
transform 1 0 5428 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_59
timestamp 1644511149
transform 1 0 6532 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_67
timestamp 1644511149
transform 1 0 7268 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_79
timestamp 1644511149
transform 1 0 8372 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_83
timestamp 1644511149
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_85
timestamp 1644511149
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_104
timestamp 1644511149
transform 1 0 10672 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_116
timestamp 1644511149
transform 1 0 11776 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_124
timestamp 1644511149
transform 1 0 12512 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_6_133
timestamp 1644511149
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_139
timestamp 1644511149
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_146
timestamp 1644511149
transform 1 0 14536 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_6_158
timestamp 1644511149
transform 1 0 15640 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_166
timestamp 1644511149
transform 1 0 16376 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_175
timestamp 1644511149
transform 1 0 17204 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_182
timestamp 1644511149
transform 1 0 17848 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_6_194
timestamp 1644511149
transform 1 0 18952 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_197
timestamp 1644511149
transform 1 0 19228 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_205
timestamp 1644511149
transform 1 0 19964 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_212
timestamp 1644511149
transform 1 0 20608 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_219
timestamp 1644511149
transform 1 0 21252 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_225
timestamp 1644511149
transform 1 0 21804 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_237
timestamp 1644511149
transform 1 0 22908 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_244
timestamp 1644511149
transform 1 0 23552 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_6_258
timestamp 1644511149
transform 1 0 24840 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_270
timestamp 1644511149
transform 1 0 25944 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_278
timestamp 1644511149
transform 1 0 26680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_286
timestamp 1644511149
transform 1 0 27416 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_298
timestamp 1644511149
transform 1 0 28520 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_306
timestamp 1644511149
transform 1 0 29256 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_309
timestamp 1644511149
transform 1 0 29532 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_317
timestamp 1644511149
transform 1 0 30268 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_323
timestamp 1644511149
transform 1 0 30820 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_6_332
timestamp 1644511149
transform 1 0 31648 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_341
timestamp 1644511149
transform 1 0 32476 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_6_354
timestamp 1644511149
transform 1 0 33672 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_362
timestamp 1644511149
transform 1 0 34408 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_365
timestamp 1644511149
transform 1 0 34684 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_369
timestamp 1644511149
transform 1 0 35052 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_383
timestamp 1644511149
transform 1 0 36340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_389
timestamp 1644511149
transform 1 0 36892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_393
timestamp 1644511149
transform 1 0 37260 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_400
timestamp 1644511149
transform 1 0 37904 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_412
timestamp 1644511149
transform 1 0 39008 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_421
timestamp 1644511149
transform 1 0 39836 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_6_429
timestamp 1644511149
transform 1 0 40572 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_437
timestamp 1644511149
transform 1 0 41308 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_6_449
timestamp 1644511149
transform 1 0 42412 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_457
timestamp 1644511149
transform 1 0 43148 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_6_466
timestamp 1644511149
transform 1 0 43976 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_6_474
timestamp 1644511149
transform 1 0 44712 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_6_477
timestamp 1644511149
transform 1 0 44988 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_489
timestamp 1644511149
transform 1 0 46092 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_501
timestamp 1644511149
transform 1 0 47196 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_513
timestamp 1644511149
transform 1 0 48300 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_6_525
timestamp 1644511149
transform 1 0 49404 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_531
timestamp 1644511149
transform 1 0 49956 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_6_533
timestamp 1644511149
transform 1 0 50140 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_545
timestamp 1644511149
transform 1 0 51244 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_6_557
timestamp 1644511149
transform 1 0 52348 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_6_569
timestamp 1644511149
transform 1 0 53452 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_572
timestamp 1644511149
transform 1 0 53728 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_6_579
timestamp 1644511149
transform 1 0 54372 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_587
timestamp 1644511149
transform 1 0 55108 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_6_589
timestamp 1644511149
transform 1 0 55292 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_592
timestamp 1644511149
transform 1 0 55568 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_6_609
timestamp 1644511149
transform 1 0 57132 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_6_617
timestamp 1644511149
transform 1 0 57868 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_7_3
timestamp 1644511149
transform 1 0 1380 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_11
timestamp 1644511149
transform 1 0 2116 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_41
timestamp 1644511149
transform 1 0 4876 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_7_53
timestamp 1644511149
transform 1 0 5980 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_57
timestamp 1644511149
transform 1 0 6348 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_61
timestamp 1644511149
transform 1 0 6716 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_69
timestamp 1644511149
transform 1 0 7452 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_79
timestamp 1644511149
transform 1 0 8372 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_91
timestamp 1644511149
transform 1 0 9476 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_7_105
timestamp 1644511149
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_111
timestamp 1644511149
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_7_113
timestamp 1644511149
transform 1 0 11500 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_119
timestamp 1644511149
transform 1 0 12052 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_122
timestamp 1644511149
transform 1 0 12328 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_129
timestamp 1644511149
transform 1 0 12972 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_133
timestamp 1644511149
transform 1 0 13340 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_137
timestamp 1644511149
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_149
timestamp 1644511149
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_161
timestamp 1644511149
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_167
timestamp 1644511149
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_174
timestamp 1644511149
transform 1 0 17112 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_181
timestamp 1644511149
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_193
timestamp 1644511149
transform 1 0 18860 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_201
timestamp 1644511149
transform 1 0 19596 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_7_216
timestamp 1644511149
transform 1 0 20976 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_225
timestamp 1644511149
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_237
timestamp 1644511149
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_255
timestamp 1644511149
transform 1 0 24564 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_267
timestamp 1644511149
transform 1 0 25668 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_273
timestamp 1644511149
transform 1 0 26220 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_276
timestamp 1644511149
transform 1 0 26496 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_281
timestamp 1644511149
transform 1 0 26956 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_294
timestamp 1644511149
transform 1 0 28152 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_306
timestamp 1644511149
transform 1 0 29256 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_318
timestamp 1644511149
transform 1 0 30360 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_7_326
timestamp 1644511149
transform 1 0 31096 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_332
timestamp 1644511149
transform 1 0 31648 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_337
timestamp 1644511149
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_349
timestamp 1644511149
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_7_361
timestamp 1644511149
transform 1 0 34316 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_7_369
timestamp 1644511149
transform 1 0 35052 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_376
timestamp 1644511149
transform 1 0 35696 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_384
timestamp 1644511149
transform 1 0 36432 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_398
timestamp 1644511149
transform 1 0 37720 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_412
timestamp 1644511149
transform 1 0 39008 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_7_429
timestamp 1644511149
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_7_441
timestamp 1644511149
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_7_447
timestamp 1644511149
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_449
timestamp 1644511149
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_467
timestamp 1644511149
transform 1 0 44068 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_479
timestamp 1644511149
transform 1 0 45172 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_491
timestamp 1644511149
transform 1 0 46276 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_503
timestamp 1644511149
transform 1 0 47380 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_518
timestamp 1644511149
transform 1 0 48760 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_522
timestamp 1644511149
transform 1 0 49128 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_7_536
timestamp 1644511149
transform 1 0 50416 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_7_548
timestamp 1644511149
transform 1 0 51520 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_7_561
timestamp 1644511149
transform 1 0 52716 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_565
timestamp 1644511149
transform 1 0 53084 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_568
timestamp 1644511149
transform 1 0 53360 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_579
timestamp 1644511149
transform 1 0 54372 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_591
timestamp 1644511149
transform 1 0 55476 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_595
timestamp 1644511149
transform 1 0 55844 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_601
timestamp 1644511149
transform 1 0 56396 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_611
timestamp 1644511149
transform 1 0 57316 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_615
timestamp 1644511149
transform 1 0 57684 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_621
timestamp 1644511149
transform 1 0 58236 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1644511149
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_15
timestamp 1644511149
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_8_27
timestamp 1644511149
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_29
timestamp 1644511149
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_41
timestamp 1644511149
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_53
timestamp 1644511149
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_65
timestamp 1644511149
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_77
timestamp 1644511149
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_83
timestamp 1644511149
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_85
timestamp 1644511149
transform 1 0 8924 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_91
timestamp 1644511149
transform 1 0 9476 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_99
timestamp 1644511149
transform 1 0 10212 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_106
timestamp 1644511149
transform 1 0 10856 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_112
timestamp 1644511149
transform 1 0 11408 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_124
timestamp 1644511149
transform 1 0 12512 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_135
timestamp 1644511149
transform 1 0 13524 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_139
timestamp 1644511149
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_145
timestamp 1644511149
transform 1 0 14444 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_157
timestamp 1644511149
transform 1 0 15548 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_165
timestamp 1644511149
transform 1 0 16284 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_172
timestamp 1644511149
transform 1 0 16928 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_178
timestamp 1644511149
transform 1 0 17480 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_190
timestamp 1644511149
transform 1 0 18584 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_8_197
timestamp 1644511149
transform 1 0 19228 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_8_209
timestamp 1644511149
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_221
timestamp 1644511149
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_233
timestamp 1644511149
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_245
timestamp 1644511149
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_251
timestamp 1644511149
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_8_253
timestamp 1644511149
transform 1 0 24380 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_276
timestamp 1644511149
transform 1 0 26496 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_280
timestamp 1644511149
transform 1 0 26864 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_8_283
timestamp 1644511149
transform 1 0 27140 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_289
timestamp 1644511149
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_8_301
timestamp 1644511149
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_307
timestamp 1644511149
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_309
timestamp 1644511149
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_321
timestamp 1644511149
transform 1 0 30636 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_325
timestamp 1644511149
transform 1 0 31004 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_329
timestamp 1644511149
transform 1 0 31372 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_341
timestamp 1644511149
transform 1 0 32476 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_353
timestamp 1644511149
transform 1 0 33580 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_361
timestamp 1644511149
transform 1 0 34316 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_8_365
timestamp 1644511149
transform 1 0 34684 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_373
timestamp 1644511149
transform 1 0 35420 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_380
timestamp 1644511149
transform 1 0 36064 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_392
timestamp 1644511149
transform 1 0 37168 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_8_404
timestamp 1644511149
transform 1 0 38272 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_410
timestamp 1644511149
transform 1 0 38824 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_416
timestamp 1644511149
transform 1 0 39376 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_8_425
timestamp 1644511149
transform 1 0 40204 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_437
timestamp 1644511149
transform 1 0 41308 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_449
timestamp 1644511149
transform 1 0 42412 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_461
timestamp 1644511149
transform 1 0 43516 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_8_473
timestamp 1644511149
transform 1 0 44620 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_8_477
timestamp 1644511149
transform 1 0 44988 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_8_484
timestamp 1644511149
transform 1 0 45632 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_8_496
timestamp 1644511149
transform 1 0 46736 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_504
timestamp 1644511149
transform 1 0 47472 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_513
timestamp 1644511149
transform 1 0 48300 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_523
timestamp 1644511149
transform 1 0 49220 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_531
timestamp 1644511149
transform 1 0 49956 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_8_533
timestamp 1644511149
transform 1 0 50140 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_545
timestamp 1644511149
transform 1 0 51244 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_557
timestamp 1644511149
transform 1 0 52348 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_8_569
timestamp 1644511149
transform 1 0 53452 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_8_584
timestamp 1644511149
transform 1 0 54832 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_606
timestamp 1644511149
transform 1 0 56856 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_8_612
timestamp 1644511149
transform 1 0 57408 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_8_618
timestamp 1644511149
transform 1 0 57960 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_624
timestamp 1644511149
transform 1 0 58512 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1644511149
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1644511149
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_27
timestamp 1644511149
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_39
timestamp 1644511149
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_51
timestamp 1644511149
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_55
timestamp 1644511149
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_64
timestamp 1644511149
transform 1 0 6992 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_76
timestamp 1644511149
transform 1 0 8096 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_88
timestamp 1644511149
transform 1 0 9200 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_96
timestamp 1644511149
transform 1 0 9936 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_106
timestamp 1644511149
transform 1 0 10856 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_9_115
timestamp 1644511149
transform 1 0 11684 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_127
timestamp 1644511149
transform 1 0 12788 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_134
timestamp 1644511149
transform 1 0 13432 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_144
timestamp 1644511149
transform 1 0 14352 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_156
timestamp 1644511149
transform 1 0 15456 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_9_174
timestamp 1644511149
transform 1 0 17112 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_183
timestamp 1644511149
transform 1 0 17940 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_9_196
timestamp 1644511149
transform 1 0 19136 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_208
timestamp 1644511149
transform 1 0 20240 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_213
timestamp 1644511149
transform 1 0 20700 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_221
timestamp 1644511149
transform 1 0 21436 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_225
timestamp 1644511149
transform 1 0 21804 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_233
timestamp 1644511149
transform 1 0 22540 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_241
timestamp 1644511149
transform 1 0 23276 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_267
timestamp 1644511149
transform 1 0 25668 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_273
timestamp 1644511149
transform 1 0 26220 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_279
timestamp 1644511149
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_281
timestamp 1644511149
transform 1 0 26956 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_286
timestamp 1644511149
transform 1 0 27416 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_297
timestamp 1644511149
transform 1 0 28428 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_304
timestamp 1644511149
transform 1 0 29072 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_316
timestamp 1644511149
transform 1 0 30176 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_326
timestamp 1644511149
transform 1 0 31096 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_332
timestamp 1644511149
transform 1 0 31648 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_337
timestamp 1644511149
transform 1 0 32108 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_341
timestamp 1644511149
transform 1 0 32476 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_358
timestamp 1644511149
transform 1 0 34040 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_369
timestamp 1644511149
transform 1 0 35052 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_373
timestamp 1644511149
transform 1 0 35420 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_381
timestamp 1644511149
transform 1 0 36156 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_389
timestamp 1644511149
transform 1 0 36892 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_393
timestamp 1644511149
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_409
timestamp 1644511149
transform 1 0 38732 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_417
timestamp 1644511149
transform 1 0 39468 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_9_421
timestamp 1644511149
transform 1 0 39836 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_433
timestamp 1644511149
transform 1 0 40940 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_445
timestamp 1644511149
transform 1 0 42044 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_9_449
timestamp 1644511149
transform 1 0 42412 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_463
timestamp 1644511149
transform 1 0 43700 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_9_475
timestamp 1644511149
transform 1 0 44804 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_489
timestamp 1644511149
transform 1 0 46092 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_9_501
timestamp 1644511149
transform 1 0 47196 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_505
timestamp 1644511149
transform 1 0 47564 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_517
timestamp 1644511149
transform 1 0 48668 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_529
timestamp 1644511149
transform 1 0 49772 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_541
timestamp 1644511149
transform 1 0 50876 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_556
timestamp 1644511149
transform 1 0 52256 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_9_561
timestamp 1644511149
transform 1 0 52716 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_573
timestamp 1644511149
transform 1 0 53820 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_9_585
timestamp 1644511149
transform 1 0 54924 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_593
timestamp 1644511149
transform 1 0 55660 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_596
timestamp 1644511149
transform 1 0 55936 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_9_604
timestamp 1644511149
transform 1 0 56672 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_612
timestamp 1644511149
transform 1 0 57408 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_9_617
timestamp 1644511149
transform 1 0 57868 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_9_621
timestamp 1644511149
transform 1 0 58236 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1644511149
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1644511149
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_10_27
timestamp 1644511149
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_35
timestamp 1644511149
transform 1 0 4324 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_47
timestamp 1644511149
transform 1 0 5428 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_10_59
timestamp 1644511149
transform 1 0 6532 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_67
timestamp 1644511149
transform 1 0 7268 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_77
timestamp 1644511149
transform 1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_83
timestamp 1644511149
transform 1 0 8740 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_85
timestamp 1644511149
transform 1 0 8924 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_10_97
timestamp 1644511149
transform 1 0 10028 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_108
timestamp 1644511149
transform 1 0 11040 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_115
timestamp 1644511149
transform 1 0 11684 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_121
timestamp 1644511149
transform 1 0 12236 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_133
timestamp 1644511149
transform 1 0 13340 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_139
timestamp 1644511149
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_154
timestamp 1644511149
transform 1 0 15272 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_179
timestamp 1644511149
transform 1 0 17572 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_187
timestamp 1644511149
transform 1 0 18308 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_195
timestamp 1644511149
transform 1 0 19044 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_197
timestamp 1644511149
transform 1 0 19228 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_203
timestamp 1644511149
transform 1 0 19780 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_211
timestamp 1644511149
transform 1 0 20516 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_217
timestamp 1644511149
transform 1 0 21068 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_224
timestamp 1644511149
transform 1 0 21712 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_228
timestamp 1644511149
transform 1 0 22080 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_242
timestamp 1644511149
transform 1 0 23368 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_248
timestamp 1644511149
transform 1 0 23920 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_253
timestamp 1644511149
transform 1 0 24380 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_265
timestamp 1644511149
transform 1 0 25484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_277
timestamp 1644511149
transform 1 0 26588 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_291
timestamp 1644511149
transform 1 0 27876 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_302
timestamp 1644511149
transform 1 0 28888 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_10_309
timestamp 1644511149
transform 1 0 29532 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_10_317
timestamp 1644511149
transform 1 0 30268 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_327
timestamp 1644511149
transform 1 0 31188 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_338
timestamp 1644511149
transform 1 0 32200 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_352
timestamp 1644511149
transform 1 0 33488 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_10_359
timestamp 1644511149
transform 1 0 34132 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_363
timestamp 1644511149
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_10_367
timestamp 1644511149
transform 1 0 34868 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_375
timestamp 1644511149
transform 1 0 35604 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_381
timestamp 1644511149
transform 1 0 36156 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_393
timestamp 1644511149
transform 1 0 37260 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_405
timestamp 1644511149
transform 1 0 38364 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_416
timestamp 1644511149
transform 1 0 39376 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_10_434
timestamp 1644511149
transform 1 0 41032 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_440
timestamp 1644511149
transform 1 0 41584 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_444
timestamp 1644511149
transform 1 0 41952 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_456
timestamp 1644511149
transform 1 0 43056 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_468
timestamp 1644511149
transform 1 0 44160 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_10_477
timestamp 1644511149
transform 1 0 44988 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_494
timestamp 1644511149
transform 1 0 46552 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_10_506
timestamp 1644511149
transform 1 0 47656 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_512
timestamp 1644511149
transform 1 0 48208 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_520
timestamp 1644511149
transform 1 0 48944 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_533
timestamp 1644511149
transform 1 0 50140 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_545
timestamp 1644511149
transform 1 0 51244 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_10_559
timestamp 1644511149
transform 1 0 52532 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_571
timestamp 1644511149
transform 1 0 53636 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_10_583
timestamp 1644511149
transform 1 0 54740 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_587
timestamp 1644511149
transform 1 0 55108 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_10_589
timestamp 1644511149
transform 1 0 55292 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_10_601
timestamp 1644511149
transform 1 0 56396 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_10_609
timestamp 1644511149
transform 1 0 57132 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_10_621
timestamp 1644511149
transform 1 0 58236 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_7
timestamp 1644511149
transform 1 0 1748 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_13
timestamp 1644511149
transform 1 0 2300 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_22
timestamp 1644511149
transform 1 0 3128 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_32
timestamp 1644511149
transform 1 0 4048 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_39
timestamp 1644511149
transform 1 0 4692 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_51
timestamp 1644511149
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_55
timestamp 1644511149
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_65
timestamp 1644511149
transform 1 0 7084 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_77
timestamp 1644511149
transform 1 0 8188 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_82
timestamp 1644511149
transform 1 0 8648 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_94
timestamp 1644511149
transform 1 0 9752 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_106
timestamp 1644511149
transform 1 0 10856 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_11_113
timestamp 1644511149
transform 1 0 11500 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_11_117
timestamp 1644511149
transform 1 0 11868 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_129
timestamp 1644511149
transform 1 0 12972 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_141
timestamp 1644511149
transform 1 0 14076 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_153
timestamp 1644511149
transform 1 0 15180 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_165
timestamp 1644511149
transform 1 0 16284 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_169
timestamp 1644511149
transform 1 0 16652 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_177
timestamp 1644511149
transform 1 0 17388 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_11_181
timestamp 1644511149
transform 1 0 17756 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_11_189
timestamp 1644511149
transform 1 0 18492 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_195
timestamp 1644511149
transform 1 0 19044 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_198
timestamp 1644511149
transform 1 0 19320 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_210
timestamp 1644511149
transform 1 0 20424 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_11_218
timestamp 1644511149
transform 1 0 21160 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_11_225
timestamp 1644511149
transform 1 0 21804 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_237
timestamp 1644511149
transform 1 0 22908 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_249
timestamp 1644511149
transform 1 0 24012 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_253
timestamp 1644511149
transform 1 0 24380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_256
timestamp 1644511149
transform 1 0 24656 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_268
timestamp 1644511149
transform 1 0 25760 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_281
timestamp 1644511149
transform 1 0 26956 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_293
timestamp 1644511149
transform 1 0 28060 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_304
timestamp 1644511149
transform 1 0 29072 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_310
timestamp 1644511149
transform 1 0 29624 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_322
timestamp 1644511149
transform 1 0 30728 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_11_328
timestamp 1644511149
transform 1 0 31280 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_331
timestamp 1644511149
transform 1 0 31556 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_335
timestamp 1644511149
transform 1 0 31924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_337
timestamp 1644511149
transform 1 0 32108 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_349
timestamp 1644511149
transform 1 0 33212 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_361
timestamp 1644511149
transform 1 0 34316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_367
timestamp 1644511149
transform 1 0 34868 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_11_379
timestamp 1644511149
transform 1 0 35972 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_384
timestamp 1644511149
transform 1 0 36432 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_393
timestamp 1644511149
transform 1 0 37260 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_408
timestamp 1644511149
transform 1 0 38640 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_11_420
timestamp 1644511149
transform 1 0 39744 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_427
timestamp 1644511149
transform 1 0 40388 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_11_439
timestamp 1644511149
transform 1 0 41492 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_447
timestamp 1644511149
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_456
timestamp 1644511149
transform 1 0 43056 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_468
timestamp 1644511149
transform 1 0 44160 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_11_480
timestamp 1644511149
transform 1 0 45264 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_11_493
timestamp 1644511149
transform 1 0 46460 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_501
timestamp 1644511149
transform 1 0 47196 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_505
timestamp 1644511149
transform 1 0 47564 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_513
timestamp 1644511149
transform 1 0 48300 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_11_522
timestamp 1644511149
transform 1 0 49128 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_534
timestamp 1644511149
transform 1 0 50232 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_11_546
timestamp 1644511149
transform 1 0 51336 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_550
timestamp 1644511149
transform 1 0 51704 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_558
timestamp 1644511149
transform 1 0 52440 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_574
timestamp 1644511149
transform 1 0 53912 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_11_585
timestamp 1644511149
transform 1 0 54924 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_597
timestamp 1644511149
transform 1 0 56028 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_612
timestamp 1644511149
transform 1 0 57408 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_11_617
timestamp 1644511149
transform 1 0 57868 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1644511149
transform 1 0 1380 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_15
timestamp 1644511149
transform 1 0 2484 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_24
timestamp 1644511149
transform 1 0 3312 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_34
timestamp 1644511149
transform 1 0 4232 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_46
timestamp 1644511149
transform 1 0 5336 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_54
timestamp 1644511149
transform 1 0 6072 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_60
timestamp 1644511149
transform 1 0 6624 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_72
timestamp 1644511149
transform 1 0 7728 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_12_76
timestamp 1644511149
transform 1 0 8096 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_80
timestamp 1644511149
transform 1 0 8464 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_92
timestamp 1644511149
transform 1 0 9568 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_98
timestamp 1644511149
transform 1 0 10120 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_109
timestamp 1644511149
transform 1 0 11132 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_121
timestamp 1644511149
transform 1 0 12236 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_133
timestamp 1644511149
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_139
timestamp 1644511149
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_12_141
timestamp 1644511149
transform 1 0 14076 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_155
timestamp 1644511149
transform 1 0 15364 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_161
timestamp 1644511149
transform 1 0 15916 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_12_171
timestamp 1644511149
transform 1 0 16836 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_182
timestamp 1644511149
transform 1 0 17848 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_194
timestamp 1644511149
transform 1 0 18952 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_12_197
timestamp 1644511149
transform 1 0 19228 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_201
timestamp 1644511149
transform 1 0 19596 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_210
timestamp 1644511149
transform 1 0 20424 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_216
timestamp 1644511149
transform 1 0 20976 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_228
timestamp 1644511149
transform 1 0 22080 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_239
timestamp 1644511149
transform 1 0 23092 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_251
timestamp 1644511149
transform 1 0 24196 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_255
timestamp 1644511149
transform 1 0 24564 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_269
timestamp 1644511149
transform 1 0 25852 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_280
timestamp 1644511149
transform 1 0 26864 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_12_291
timestamp 1644511149
transform 1 0 27876 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_304
timestamp 1644511149
transform 1 0 29072 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_316
timestamp 1644511149
transform 1 0 30176 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_324
timestamp 1644511149
transform 1 0 30912 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_336
timestamp 1644511149
transform 1 0 32016 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_12_345
timestamp 1644511149
transform 1 0 32844 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_351
timestamp 1644511149
transform 1 0 33396 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_363
timestamp 1644511149
transform 1 0 34500 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_378
timestamp 1644511149
transform 1 0 35880 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_391
timestamp 1644511149
transform 1 0 37076 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_12_400
timestamp 1644511149
transform 1 0 37904 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_12_408
timestamp 1644511149
transform 1 0 38640 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_12_412
timestamp 1644511149
transform 1 0 39008 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_12_421
timestamp 1644511149
transform 1 0 39836 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_12_449
timestamp 1644511149
transform 1 0 42412 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_455
timestamp 1644511149
transform 1 0 42964 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_467
timestamp 1644511149
transform 1 0 44068 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_475
timestamp 1644511149
transform 1 0 44804 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_490
timestamp 1644511149
transform 1 0 46184 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_502
timestamp 1644511149
transform 1 0 47288 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_12_514
timestamp 1644511149
transform 1 0 48392 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_520
timestamp 1644511149
transform 1 0 48944 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_528
timestamp 1644511149
transform 1 0 49680 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_533
timestamp 1644511149
transform 1 0 50140 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_12_545
timestamp 1644511149
transform 1 0 51244 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_555
timestamp 1644511149
transform 1 0 52164 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_12_567
timestamp 1644511149
transform 1 0 53268 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_12_575
timestamp 1644511149
transform 1 0 54004 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_12_581
timestamp 1644511149
transform 1 0 54556 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_587
timestamp 1644511149
transform 1 0 55108 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_589
timestamp 1644511149
transform 1 0 55292 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_597
timestamp 1644511149
transform 1 0 56028 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_611
timestamp 1644511149
transform 1 0 57316 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_12_623
timestamp 1644511149
transform 1 0 58420 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1644511149
transform 1 0 1380 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_15
timestamp 1644511149
transform 1 0 2484 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_13_38
timestamp 1644511149
transform 1 0 4600 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_50
timestamp 1644511149
transform 1 0 5704 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_13_64
timestamp 1644511149
transform 1 0 6992 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_76
timestamp 1644511149
transform 1 0 8096 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_87
timestamp 1644511149
transform 1 0 9108 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_93
timestamp 1644511149
transform 1 0 9660 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_105
timestamp 1644511149
transform 1 0 10764 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_111
timestamp 1644511149
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_116
timestamp 1644511149
transform 1 0 11776 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_142
timestamp 1644511149
transform 1 0 14168 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_156
timestamp 1644511149
transform 1 0 15456 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_162
timestamp 1644511149
transform 1 0 16008 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_13_169
timestamp 1644511149
transform 1 0 16652 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_13_181
timestamp 1644511149
transform 1 0 17756 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_186
timestamp 1644511149
transform 1 0 18216 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_190
timestamp 1644511149
transform 1 0 18584 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_198
timestamp 1644511149
transform 1 0 19320 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_206
timestamp 1644511149
transform 1 0 20056 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_214
timestamp 1644511149
transform 1 0 20792 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_222
timestamp 1644511149
transform 1 0 21528 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_13_225
timestamp 1644511149
transform 1 0 21804 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_13_240
timestamp 1644511149
transform 1 0 23184 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_251
timestamp 1644511149
transform 1 0 24196 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_255
timestamp 1644511149
transform 1 0 24564 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_259
timestamp 1644511149
transform 1 0 24932 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_270
timestamp 1644511149
transform 1 0 25944 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_13_278
timestamp 1644511149
transform 1 0 26680 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_13_281
timestamp 1644511149
transform 1 0 26956 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_285
timestamp 1644511149
transform 1 0 27324 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_288
timestamp 1644511149
transform 1 0 27600 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_13_302
timestamp 1644511149
transform 1 0 28888 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_13_318
timestamp 1644511149
transform 1 0 30360 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_330
timestamp 1644511149
transform 1 0 31464 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_13_337
timestamp 1644511149
transform 1 0 32108 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_349
timestamp 1644511149
transform 1 0 33212 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_13_361
timestamp 1644511149
transform 1 0 34316 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_369
timestamp 1644511149
transform 1 0 35052 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_374
timestamp 1644511149
transform 1 0 35512 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_386
timestamp 1644511149
transform 1 0 36616 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_13_393
timestamp 1644511149
transform 1 0 37260 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_405
timestamp 1644511149
transform 1 0 38364 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_417
timestamp 1644511149
transform 1 0 39468 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_429
timestamp 1644511149
transform 1 0 40572 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_444
timestamp 1644511149
transform 1 0 41952 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_13_449
timestamp 1644511149
transform 1 0 42412 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_457
timestamp 1644511149
transform 1 0 43148 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_465
timestamp 1644511149
transform 1 0 43884 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_471
timestamp 1644511149
transform 1 0 44436 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_13_492
timestamp 1644511149
transform 1 0 46368 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_505
timestamp 1644511149
transform 1 0 47564 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_517
timestamp 1644511149
transform 1 0 48668 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_529
timestamp 1644511149
transform 1 0 49772 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_541
timestamp 1644511149
transform 1 0 50876 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_13_553
timestamp 1644511149
transform 1 0 51980 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_13_559
timestamp 1644511149
transform 1 0 52532 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_561
timestamp 1644511149
transform 1 0 52716 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_573
timestamp 1644511149
transform 1 0 53820 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_13_581
timestamp 1644511149
transform 1 0 54556 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_13_590
timestamp 1644511149
transform 1 0 55384 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_594
timestamp 1644511149
transform 1 0 55752 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_601
timestamp 1644511149
transform 1 0 56396 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_13_613
timestamp 1644511149
transform 1 0 57500 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_13_617
timestamp 1644511149
transform 1 0 57868 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_14_5
timestamp 1644511149
transform 1 0 1564 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_17
timestamp 1644511149
transform 1 0 2668 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_23
timestamp 1644511149
transform 1 0 3220 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_27
timestamp 1644511149
transform 1 0 3588 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_32
timestamp 1644511149
transform 1 0 4048 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_44
timestamp 1644511149
transform 1 0 5152 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_54
timestamp 1644511149
transform 1 0 6072 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_63
timestamp 1644511149
transform 1 0 6900 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_75
timestamp 1644511149
transform 1 0 8004 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_83
timestamp 1644511149
transform 1 0 8740 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_92
timestamp 1644511149
transform 1 0 9568 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_98
timestamp 1644511149
transform 1 0 10120 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_110
timestamp 1644511149
transform 1 0 11224 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_118
timestamp 1644511149
transform 1 0 11960 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_126
timestamp 1644511149
transform 1 0 12696 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_138
timestamp 1644511149
transform 1 0 13800 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_154
timestamp 1644511149
transform 1 0 15272 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_164
timestamp 1644511149
transform 1 0 16192 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_174
timestamp 1644511149
transform 1 0 17112 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_186
timestamp 1644511149
transform 1 0 18216 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_194
timestamp 1644511149
transform 1 0 18952 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_14_200
timestamp 1644511149
transform 1 0 19504 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_14_212
timestamp 1644511149
transform 1 0 20608 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_14_219
timestamp 1644511149
transform 1 0 21252 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_226
timestamp 1644511149
transform 1 0 21896 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_230
timestamp 1644511149
transform 1 0 22264 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_238
timestamp 1644511149
transform 1 0 23000 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_14_250
timestamp 1644511149
transform 1 0 24104 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_14_253
timestamp 1644511149
transform 1 0 24380 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_256
timestamp 1644511149
transform 1 0 24656 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_264
timestamp 1644511149
transform 1 0 25392 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_277
timestamp 1644511149
transform 1 0 26588 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_289
timestamp 1644511149
transform 1 0 27692 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_293
timestamp 1644511149
transform 1 0 28060 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_304
timestamp 1644511149
transform 1 0 29072 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_309
timestamp 1644511149
transform 1 0 29532 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_317
timestamp 1644511149
transform 1 0 30268 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_329
timestamp 1644511149
transform 1 0 31372 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_335
timestamp 1644511149
transform 1 0 31924 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_338
timestamp 1644511149
transform 1 0 32200 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_355
timestamp 1644511149
transform 1 0 33764 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_363
timestamp 1644511149
transform 1 0 34500 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_365
timestamp 1644511149
transform 1 0 34684 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_373
timestamp 1644511149
transform 1 0 35420 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_377
timestamp 1644511149
transform 1 0 35788 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_388
timestamp 1644511149
transform 1 0 36800 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_400
timestamp 1644511149
transform 1 0 37904 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_406
timestamp 1644511149
transform 1 0 38456 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_412
timestamp 1644511149
transform 1 0 39008 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_14_423
timestamp 1644511149
transform 1 0 40020 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_14_431
timestamp 1644511149
transform 1 0 40756 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_14_437
timestamp 1644511149
transform 1 0 41308 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_447
timestamp 1644511149
transform 1 0 42228 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_14_458
timestamp 1644511149
transform 1 0 43240 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_470
timestamp 1644511149
transform 1 0 44344 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_477
timestamp 1644511149
transform 1 0 44988 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_481
timestamp 1644511149
transform 1 0 45356 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_14_489
timestamp 1644511149
transform 1 0 46092 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_501
timestamp 1644511149
transform 1 0 47196 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_14_516
timestamp 1644511149
transform 1 0 48576 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_527
timestamp 1644511149
transform 1 0 49588 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_531
timestamp 1644511149
transform 1 0 49956 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_533
timestamp 1644511149
transform 1 0 50140 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_14_541
timestamp 1644511149
transform 1 0 50876 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_551
timestamp 1644511149
transform 1 0 51796 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_14_563
timestamp 1644511149
transform 1 0 52900 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_14_571
timestamp 1644511149
transform 1 0 53636 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_14_583
timestamp 1644511149
transform 1 0 54740 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_587
timestamp 1644511149
transform 1 0 55108 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_14_589
timestamp 1644511149
transform 1 0 55292 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_14_596
timestamp 1644511149
transform 1 0 55936 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_604
timestamp 1644511149
transform 1 0 56672 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_610
timestamp 1644511149
transform 1 0 57224 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_614
timestamp 1644511149
transform 1 0 57592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_14_617
timestamp 1644511149
transform 1 0 57868 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_15_6
timestamp 1644511149
transform 1 0 1656 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_14
timestamp 1644511149
transform 1 0 2392 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_28
timestamp 1644511149
transform 1 0 3680 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_37
timestamp 1644511149
transform 1 0 4508 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_15_49
timestamp 1644511149
transform 1 0 5612 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_55
timestamp 1644511149
transform 1 0 6164 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_62
timestamp 1644511149
transform 1 0 6808 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_74
timestamp 1644511149
transform 1 0 7912 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_86
timestamp 1644511149
transform 1 0 9016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_92
timestamp 1644511149
transform 1 0 9568 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_99
timestamp 1644511149
transform 1 0 10212 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_105
timestamp 1644511149
transform 1 0 10764 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_111
timestamp 1644511149
transform 1 0 11316 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_15_113
timestamp 1644511149
transform 1 0 11500 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_123
timestamp 1644511149
transform 1 0 12420 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_132
timestamp 1644511149
transform 1 0 13248 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_140
timestamp 1644511149
transform 1 0 13984 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_145
timestamp 1644511149
transform 1 0 14444 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_153
timestamp 1644511149
transform 1 0 15180 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_15_159
timestamp 1644511149
transform 1 0 15732 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_167
timestamp 1644511149
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_169
timestamp 1644511149
transform 1 0 16652 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_181
timestamp 1644511149
transform 1 0 17756 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_189
timestamp 1644511149
transform 1 0 18492 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_192
timestamp 1644511149
transform 1 0 18768 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_204
timestamp 1644511149
transform 1 0 19872 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_216
timestamp 1644511149
transform 1 0 20976 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_15_225
timestamp 1644511149
transform 1 0 21804 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_233
timestamp 1644511149
transform 1 0 22540 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_15_242
timestamp 1644511149
transform 1 0 23368 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_250
timestamp 1644511149
transform 1 0 24104 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_255
timestamp 1644511149
transform 1 0 24564 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_266
timestamp 1644511149
transform 1 0 25576 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_274
timestamp 1644511149
transform 1 0 26312 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_281
timestamp 1644511149
transform 1 0 26956 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_292
timestamp 1644511149
transform 1 0 27968 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_15_304
timestamp 1644511149
transform 1 0 29072 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_15_316
timestamp 1644511149
transform 1 0 30176 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_322
timestamp 1644511149
transform 1 0 30728 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_325
timestamp 1644511149
transform 1 0 31004 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_15_333
timestamp 1644511149
transform 1 0 31740 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_15_359
timestamp 1644511149
transform 1 0 34132 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_15_374
timestamp 1644511149
transform 1 0 35512 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_380
timestamp 1644511149
transform 1 0 36064 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_387
timestamp 1644511149
transform 1 0 36708 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_391
timestamp 1644511149
transform 1 0 37076 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_406
timestamp 1644511149
transform 1 0 38456 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_415
timestamp 1644511149
transform 1 0 39284 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_424
timestamp 1644511149
transform 1 0 40112 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_435
timestamp 1644511149
transform 1 0 41124 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_447
timestamp 1644511149
transform 1 0 42228 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_451
timestamp 1644511149
transform 1 0 42596 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_463
timestamp 1644511149
transform 1 0 43700 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_475
timestamp 1644511149
transform 1 0 44804 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_487
timestamp 1644511149
transform 1 0 45908 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_499
timestamp 1644511149
transform 1 0 47012 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_503
timestamp 1644511149
transform 1 0 47380 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_505
timestamp 1644511149
transform 1 0 47564 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_511
timestamp 1644511149
transform 1 0 48116 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_528
timestamp 1644511149
transform 1 0 49680 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_15_540
timestamp 1644511149
transform 1 0 50784 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_15_556
timestamp 1644511149
transform 1 0 52256 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_567
timestamp 1644511149
transform 1 0 53268 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_15_576
timestamp 1644511149
transform 1 0 54096 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_583
timestamp 1644511149
transform 1 0 54740 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_15_595
timestamp 1644511149
transform 1 0 55844 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_601
timestamp 1644511149
transform 1 0 56396 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_610
timestamp 1644511149
transform 1 0 57224 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_621
timestamp 1644511149
transform 1 0 58236 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1644511149
transform 1 0 1380 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_15
timestamp 1644511149
transform 1 0 2484 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_23
timestamp 1644511149
transform 1 0 3220 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_27
timestamp 1644511149
transform 1 0 3588 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_32
timestamp 1644511149
transform 1 0 4048 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_44
timestamp 1644511149
transform 1 0 5152 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_56
timestamp 1644511149
transform 1 0 6256 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_68
timestamp 1644511149
transform 1 0 7360 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_80
timestamp 1644511149
transform 1 0 8464 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_85
timestamp 1644511149
transform 1 0 8924 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_91
timestamp 1644511149
transform 1 0 9476 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_94
timestamp 1644511149
transform 1 0 9752 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_106
timestamp 1644511149
transform 1 0 10856 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_123
timestamp 1644511149
transform 1 0 12420 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_135
timestamp 1644511149
transform 1 0 13524 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_139
timestamp 1644511149
transform 1 0 13892 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_141
timestamp 1644511149
transform 1 0 14076 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_151
timestamp 1644511149
transform 1 0 14996 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_157
timestamp 1644511149
transform 1 0 15548 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_164
timestamp 1644511149
transform 1 0 16192 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_175
timestamp 1644511149
transform 1 0 17204 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_183
timestamp 1644511149
transform 1 0 17940 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_195
timestamp 1644511149
transform 1 0 19044 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_197
timestamp 1644511149
transform 1 0 19228 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_209
timestamp 1644511149
transform 1 0 20332 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_16_221
timestamp 1644511149
transform 1 0 21436 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_231
timestamp 1644511149
transform 1 0 22356 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_239
timestamp 1644511149
transform 1 0 23092 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_251
timestamp 1644511149
transform 1 0 24196 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_253
timestamp 1644511149
transform 1 0 24380 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_261
timestamp 1644511149
transform 1 0 25116 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_267
timestamp 1644511149
transform 1 0 25668 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_279
timestamp 1644511149
transform 1 0 26772 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_294
timestamp 1644511149
transform 1 0 28152 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_306
timestamp 1644511149
transform 1 0 29256 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_309
timestamp 1644511149
transform 1 0 29532 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_323
timestamp 1644511149
transform 1 0 30820 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_333
timestamp 1644511149
transform 1 0 31740 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_16_345
timestamp 1644511149
transform 1 0 32844 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_353
timestamp 1644511149
transform 1 0 33580 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_358
timestamp 1644511149
transform 1 0 34040 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_375
timestamp 1644511149
transform 1 0 35604 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_16_382
timestamp 1644511149
transform 1 0 36248 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_394
timestamp 1644511149
transform 1 0 37352 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_406
timestamp 1644511149
transform 1 0 38456 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_414
timestamp 1644511149
transform 1 0 39192 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_421
timestamp 1644511149
transform 1 0 39836 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_425
timestamp 1644511149
transform 1 0 40204 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_428
timestamp 1644511149
transform 1 0 40480 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_16_440
timestamp 1644511149
transform 1 0 41584 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_16_449
timestamp 1644511149
transform 1 0 42412 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_463
timestamp 1644511149
transform 1 0 43700 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_16_475
timestamp 1644511149
transform 1 0 44804 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_477
timestamp 1644511149
transform 1 0 44988 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_485
timestamp 1644511149
transform 1 0 45724 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_16_492
timestamp 1644511149
transform 1 0 46368 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_504
timestamp 1644511149
transform 1 0 47472 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_508
timestamp 1644511149
transform 1 0 47840 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_518
timestamp 1644511149
transform 1 0 48760 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_525
timestamp 1644511149
transform 1 0 49404 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_531
timestamp 1644511149
transform 1 0 49956 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_533
timestamp 1644511149
transform 1 0 50140 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_16_545
timestamp 1644511149
transform 1 0 51244 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_549
timestamp 1644511149
transform 1 0 51612 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_553
timestamp 1644511149
transform 1 0 51980 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_16_578
timestamp 1644511149
transform 1 0 54280 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_586
timestamp 1644511149
transform 1 0 55016 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_16_589
timestamp 1644511149
transform 1 0 55292 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_597
timestamp 1644511149
transform 1 0 56028 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_607
timestamp 1644511149
transform 1 0 56948 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_614
timestamp 1644511149
transform 1 0 57592 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_621
timestamp 1644511149
transform 1 0 58236 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_3
timestamp 1644511149
transform 1 0 1380 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_15
timestamp 1644511149
transform 1 0 2484 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_26
timestamp 1644511149
transform 1 0 3496 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_33
timestamp 1644511149
transform 1 0 4140 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_45
timestamp 1644511149
transform 1 0 5244 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_52
timestamp 1644511149
transform 1 0 5888 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_60
timestamp 1644511149
transform 1 0 6624 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_17_66
timestamp 1644511149
transform 1 0 7176 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_17_74
timestamp 1644511149
transform 1 0 7912 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_81
timestamp 1644511149
transform 1 0 8556 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_90
timestamp 1644511149
transform 1 0 9384 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_96
timestamp 1644511149
transform 1 0 9936 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_108
timestamp 1644511149
transform 1 0 11040 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_113
timestamp 1644511149
transform 1 0 11500 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_136
timestamp 1644511149
transform 1 0 13616 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_148
timestamp 1644511149
transform 1 0 14720 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_152
timestamp 1644511149
transform 1 0 15088 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_160
timestamp 1644511149
transform 1 0 15824 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_17_176
timestamp 1644511149
transform 1 0 17296 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_188
timestamp 1644511149
transform 1 0 18400 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_194
timestamp 1644511149
transform 1 0 18952 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_200
timestamp 1644511149
transform 1 0 19504 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_207
timestamp 1644511149
transform 1 0 20148 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_215
timestamp 1644511149
transform 1 0 20884 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_220
timestamp 1644511149
transform 1 0 21344 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_227
timestamp 1644511149
transform 1 0 21988 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_240
timestamp 1644511149
transform 1 0 23184 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_248
timestamp 1644511149
transform 1 0 23920 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_260
timestamp 1644511149
transform 1 0 25024 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_271
timestamp 1644511149
transform 1 0 26036 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_17_279
timestamp 1644511149
transform 1 0 26772 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_281
timestamp 1644511149
transform 1 0 26956 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_293
timestamp 1644511149
transform 1 0 28060 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_301
timestamp 1644511149
transform 1 0 28796 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_312
timestamp 1644511149
transform 1 0 29808 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_320
timestamp 1644511149
transform 1 0 30544 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_17_332
timestamp 1644511149
transform 1 0 31648 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_339
timestamp 1644511149
transform 1 0 32292 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_351
timestamp 1644511149
transform 1 0 33396 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_358
timestamp 1644511149
transform 1 0 34040 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_362
timestamp 1644511149
transform 1 0 34408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_17_367
timestamp 1644511149
transform 1 0 34868 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_379
timestamp 1644511149
transform 1 0 35972 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_391
timestamp 1644511149
transform 1 0 37076 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_393
timestamp 1644511149
transform 1 0 37260 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_401
timestamp 1644511149
transform 1 0 37996 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_409
timestamp 1644511149
transform 1 0 38732 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_17_417
timestamp 1644511149
transform 1 0 39468 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_429
timestamp 1644511149
transform 1 0 40572 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_17_441
timestamp 1644511149
transform 1 0 41676 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_17_447
timestamp 1644511149
transform 1 0 42228 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_449
timestamp 1644511149
transform 1 0 42412 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_17_465
timestamp 1644511149
transform 1 0 43884 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_473
timestamp 1644511149
transform 1 0 44620 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_482
timestamp 1644511149
transform 1 0 45448 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_17_493
timestamp 1644511149
transform 1 0 46460 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_501
timestamp 1644511149
transform 1 0 47196 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_505
timestamp 1644511149
transform 1 0 47564 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_513
timestamp 1644511149
transform 1 0 48300 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_17_522
timestamp 1644511149
transform 1 0 49128 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_534
timestamp 1644511149
transform 1 0 50232 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_546
timestamp 1644511149
transform 1 0 51336 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_17_558
timestamp 1644511149
transform 1 0 52440 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_17_561
timestamp 1644511149
transform 1 0 52716 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_17_572
timestamp 1644511149
transform 1 0 53728 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_17_584
timestamp 1644511149
transform 1 0 54832 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_17_596
timestamp 1644511149
transform 1 0 55936 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_611
timestamp 1644511149
transform 1 0 57316 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_615
timestamp 1644511149
transform 1 0 57684 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_17_617
timestamp 1644511149
transform 1 0 57868 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_17_621
timestamp 1644511149
transform 1 0 58236 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_5
timestamp 1644511149
transform 1 0 1564 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_17
timestamp 1644511149
transform 1 0 2668 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_25
timestamp 1644511149
transform 1 0 3404 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_35
timestamp 1644511149
transform 1 0 4324 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_18_43
timestamp 1644511149
transform 1 0 5060 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_47
timestamp 1644511149
transform 1 0 5428 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_59
timestamp 1644511149
transform 1 0 6532 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_18_68
timestamp 1644511149
transform 1 0 7360 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_74
timestamp 1644511149
transform 1 0 7912 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_80
timestamp 1644511149
transform 1 0 8464 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_18_85
timestamp 1644511149
transform 1 0 8924 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_93
timestamp 1644511149
transform 1 0 9660 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_99
timestamp 1644511149
transform 1 0 10212 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_18_111
timestamp 1644511149
transform 1 0 11316 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_115
timestamp 1644511149
transform 1 0 11684 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_129
timestamp 1644511149
transform 1 0 12972 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_135
timestamp 1644511149
transform 1 0 13524 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_139
timestamp 1644511149
transform 1 0 13892 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_141
timestamp 1644511149
transform 1 0 14076 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_147
timestamp 1644511149
transform 1 0 14628 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_154
timestamp 1644511149
transform 1 0 15272 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_158
timestamp 1644511149
transform 1 0 15640 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_163
timestamp 1644511149
transform 1 0 16100 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_174
timestamp 1644511149
transform 1 0 17112 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_186
timestamp 1644511149
transform 1 0 18216 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_18_190
timestamp 1644511149
transform 1 0 18584 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_202
timestamp 1644511149
transform 1 0 19688 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_214
timestamp 1644511149
transform 1 0 20792 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_225
timestamp 1644511149
transform 1 0 21804 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_235
timestamp 1644511149
transform 1 0 22724 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_18_241
timestamp 1644511149
transform 1 0 23276 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_249
timestamp 1644511149
transform 1 0 24012 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_18_253
timestamp 1644511149
transform 1 0 24380 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_18_263
timestamp 1644511149
transform 1 0 25300 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_275
timestamp 1644511149
transform 1 0 26404 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_287
timestamp 1644511149
transform 1 0 27508 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_18_299
timestamp 1644511149
transform 1 0 28612 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_304
timestamp 1644511149
transform 1 0 29072 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_316
timestamp 1644511149
transform 1 0 30176 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_324
timestamp 1644511149
transform 1 0 30912 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_328
timestamp 1644511149
transform 1 0 31280 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_331
timestamp 1644511149
transform 1 0 31556 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_337
timestamp 1644511149
transform 1 0 32108 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_346
timestamp 1644511149
transform 1 0 32936 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_358
timestamp 1644511149
transform 1 0 34040 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_18_370
timestamp 1644511149
transform 1 0 35144 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_382
timestamp 1644511149
transform 1 0 36248 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_18_394
timestamp 1644511149
transform 1 0 37352 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_398
timestamp 1644511149
transform 1 0 37720 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_402
timestamp 1644511149
transform 1 0 38088 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_409
timestamp 1644511149
transform 1 0 38732 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_417
timestamp 1644511149
transform 1 0 39468 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_18_421
timestamp 1644511149
transform 1 0 39836 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_18_429
timestamp 1644511149
transform 1 0 40572 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_440
timestamp 1644511149
transform 1 0 41584 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_452
timestamp 1644511149
transform 1 0 42688 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_464
timestamp 1644511149
transform 1 0 43792 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_18_477
timestamp 1644511149
transform 1 0 44988 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_18_489
timestamp 1644511149
transform 1 0 46092 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_501
timestamp 1644511149
transform 1 0 47196 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_18_513
timestamp 1644511149
transform 1 0 48300 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_18_524
timestamp 1644511149
transform 1 0 49312 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_18_533
timestamp 1644511149
transform 1 0 50140 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_541
timestamp 1644511149
transform 1 0 50876 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_548
timestamp 1644511149
transform 1 0 51520 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_18_557
timestamp 1644511149
transform 1 0 52348 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_18_569
timestamp 1644511149
transform 1 0 53452 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_18_581
timestamp 1644511149
transform 1 0 54556 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_18_587
timestamp 1644511149
transform 1 0 55108 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_18_589
timestamp 1644511149
transform 1 0 55292 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_18_597
timestamp 1644511149
transform 1 0 56028 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_18_604
timestamp 1644511149
transform 1 0 56672 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_611
timestamp 1644511149
transform 1 0 57316 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_621
timestamp 1644511149
transform 1 0 58236 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_6
timestamp 1644511149
transform 1 0 1656 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_19_34
timestamp 1644511149
transform 1 0 4232 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_46
timestamp 1644511149
transform 1 0 5336 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_54
timestamp 1644511149
transform 1 0 6072 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_19_62
timestamp 1644511149
transform 1 0 6808 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_70
timestamp 1644511149
transform 1 0 7544 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_75
timestamp 1644511149
transform 1 0 8004 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_96
timestamp 1644511149
transform 1 0 9936 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_102
timestamp 1644511149
transform 1 0 10488 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_108
timestamp 1644511149
transform 1 0 11040 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_113
timestamp 1644511149
transform 1 0 11500 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_125
timestamp 1644511149
transform 1 0 12604 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_132
timestamp 1644511149
transform 1 0 13248 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_138
timestamp 1644511149
transform 1 0 13800 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_144
timestamp 1644511149
transform 1 0 14352 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_148
timestamp 1644511149
transform 1 0 14720 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_151
timestamp 1644511149
transform 1 0 14996 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_157
timestamp 1644511149
transform 1 0 15548 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_165
timestamp 1644511149
transform 1 0 16284 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_174
timestamp 1644511149
transform 1 0 17112 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_182
timestamp 1644511149
transform 1 0 17848 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_186
timestamp 1644511149
transform 1 0 18216 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_197
timestamp 1644511149
transform 1 0 19228 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_203
timestamp 1644511149
transform 1 0 19780 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_215
timestamp 1644511149
transform 1 0 20884 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_223
timestamp 1644511149
transform 1 0 21620 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_225
timestamp 1644511149
transform 1 0 21804 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_239
timestamp 1644511149
transform 1 0 23092 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_247
timestamp 1644511149
transform 1 0 23828 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_250
timestamp 1644511149
transform 1 0 24104 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_261
timestamp 1644511149
transform 1 0 25116 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_19_269
timestamp 1644511149
transform 1 0 25852 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_277
timestamp 1644511149
transform 1 0 26588 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_19_281
timestamp 1644511149
transform 1 0 26956 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_19_289
timestamp 1644511149
transform 1 0 27692 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_300
timestamp 1644511149
transform 1 0 28704 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_314
timestamp 1644511149
transform 1 0 29992 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_322
timestamp 1644511149
transform 1 0 30728 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_334
timestamp 1644511149
transform 1 0 31832 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_340
timestamp 1644511149
transform 1 0 32384 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_352
timestamp 1644511149
transform 1 0 33488 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_19_364
timestamp 1644511149
transform 1 0 34592 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_19_376
timestamp 1644511149
transform 1 0 35696 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_19_388
timestamp 1644511149
transform 1 0 36800 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_393
timestamp 1644511149
transform 1 0 37260 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_397
timestamp 1644511149
transform 1 0 37628 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_404
timestamp 1644511149
transform 1 0 38272 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_19_412
timestamp 1644511149
transform 1 0 39008 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_424
timestamp 1644511149
transform 1 0 40112 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_19_432
timestamp 1644511149
transform 1 0 40848 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_19_442
timestamp 1644511149
transform 1 0 41768 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_19_455
timestamp 1644511149
transform 1 0 42964 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_467
timestamp 1644511149
transform 1 0 44068 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_475
timestamp 1644511149
transform 1 0 44804 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_19_480
timestamp 1644511149
transform 1 0 45264 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_19_492
timestamp 1644511149
transform 1 0 46368 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_19_497
timestamp 1644511149
transform 1 0 46828 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_503
timestamp 1644511149
transform 1 0 47380 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_512
timestamp 1644511149
transform 1 0 48208 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_19_524
timestamp 1644511149
transform 1 0 49312 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_19_532
timestamp 1644511149
transform 1 0 50048 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_19_536
timestamp 1644511149
transform 1 0 50416 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_545
timestamp 1644511149
transform 1 0 51244 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_555
timestamp 1644511149
transform 1 0 52164 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_19_559
timestamp 1644511149
transform 1 0 52532 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_19_561
timestamp 1644511149
transform 1 0 52716 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_19_573
timestamp 1644511149
transform 1 0 53820 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_582
timestamp 1644511149
transform 1 0 54648 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_594
timestamp 1644511149
transform 1 0 55752 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_19_609
timestamp 1644511149
transform 1 0 57132 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_615
timestamp 1644511149
transform 1 0 57684 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_617
timestamp 1644511149
transform 1 0 57868 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_3
timestamp 1644511149
transform 1 0 1380 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_24
timestamp 1644511149
transform 1 0 3312 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_29
timestamp 1644511149
transform 1 0 3772 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_20_41
timestamp 1644511149
transform 1 0 4876 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_75
timestamp 1644511149
transform 1 0 8004 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_83
timestamp 1644511149
transform 1 0 8740 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_20_85
timestamp 1644511149
transform 1 0 8924 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_94
timestamp 1644511149
transform 1 0 9752 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_100
timestamp 1644511149
transform 1 0 10304 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_106
timestamp 1644511149
transform 1 0 10856 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_114
timestamp 1644511149
transform 1 0 11592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_117
timestamp 1644511149
transform 1 0 11868 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_130
timestamp 1644511149
transform 1 0 13064 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_136
timestamp 1644511149
transform 1 0 13616 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_141
timestamp 1644511149
transform 1 0 14076 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_145
timestamp 1644511149
transform 1 0 14444 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_150
timestamp 1644511149
transform 1 0 14904 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_158
timestamp 1644511149
transform 1 0 15640 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_169
timestamp 1644511149
transform 1 0 16652 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_177
timestamp 1644511149
transform 1 0 17388 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_185
timestamp 1644511149
transform 1 0 18124 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_193
timestamp 1644511149
transform 1 0 18860 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_206
timestamp 1644511149
transform 1 0 20056 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_214
timestamp 1644511149
transform 1 0 20792 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_230
timestamp 1644511149
transform 1 0 22264 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_238
timestamp 1644511149
transform 1 0 23000 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_248
timestamp 1644511149
transform 1 0 23920 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_253
timestamp 1644511149
transform 1 0 24380 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_257
timestamp 1644511149
transform 1 0 24748 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_266
timestamp 1644511149
transform 1 0 25576 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_20_283
timestamp 1644511149
transform 1 0 27140 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_289
timestamp 1644511149
transform 1 0 27692 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_294
timestamp 1644511149
transform 1 0 28152 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_300
timestamp 1644511149
transform 1 0 28704 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_309
timestamp 1644511149
transform 1 0 29532 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_20_316
timestamp 1644511149
transform 1 0 30176 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_20_324
timestamp 1644511149
transform 1 0 30912 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_328
timestamp 1644511149
transform 1 0 31280 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_334
timestamp 1644511149
transform 1 0 31832 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_344
timestamp 1644511149
transform 1 0 32752 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_356
timestamp 1644511149
transform 1 0 33856 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_365
timestamp 1644511149
transform 1 0 34684 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_369
timestamp 1644511149
transform 1 0 35052 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_383
timestamp 1644511149
transform 1 0 36340 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_395
timestamp 1644511149
transform 1 0 37444 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_403
timestamp 1644511149
transform 1 0 38180 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_408
timestamp 1644511149
transform 1 0 38640 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_20_421
timestamp 1644511149
transform 1 0 39836 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_20_436
timestamp 1644511149
transform 1 0 41216 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_444
timestamp 1644511149
transform 1 0 41952 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_20_460
timestamp 1644511149
transform 1 0 43424 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_472
timestamp 1644511149
transform 1 0 44528 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_20_483
timestamp 1644511149
transform 1 0 45540 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_20_491
timestamp 1644511149
transform 1 0 46276 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_20_507
timestamp 1644511149
transform 1 0 47748 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_511
timestamp 1644511149
transform 1 0 48116 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_525
timestamp 1644511149
transform 1 0 49404 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_531
timestamp 1644511149
transform 1 0 49956 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_20_533
timestamp 1644511149
transform 1 0 50140 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_537
timestamp 1644511149
transform 1 0 50508 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_545
timestamp 1644511149
transform 1 0 51244 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_557
timestamp 1644511149
transform 1 0 52348 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_563
timestamp 1644511149
transform 1 0 52900 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_20_570
timestamp 1644511149
transform 1 0 53544 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_20_582
timestamp 1644511149
transform 1 0 54648 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_20_589
timestamp 1644511149
transform 1 0 55292 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_20_601
timestamp 1644511149
transform 1 0 56396 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_20_610
timestamp 1644511149
transform 1 0 57224 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_20_622
timestamp 1644511149
transform 1 0 58328 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_3
timestamp 1644511149
transform 1 0 1380 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_15
timestamp 1644511149
transform 1 0 2484 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_41
timestamp 1644511149
transform 1 0 4876 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_47
timestamp 1644511149
transform 1 0 5428 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_55
timestamp 1644511149
transform 1 0 6164 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_57
timestamp 1644511149
transform 1 0 6348 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_69
timestamp 1644511149
transform 1 0 7452 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_77
timestamp 1644511149
transform 1 0 8188 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_103
timestamp 1644511149
transform 1 0 10580 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_111
timestamp 1644511149
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_115
timestamp 1644511149
transform 1 0 11684 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_123
timestamp 1644511149
transform 1 0 12420 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_129
timestamp 1644511149
transform 1 0 12972 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_139
timestamp 1644511149
transform 1 0 13892 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_145
timestamp 1644511149
transform 1 0 14444 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_153
timestamp 1644511149
transform 1 0 15180 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_164
timestamp 1644511149
transform 1 0 16192 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_179
timestamp 1644511149
transform 1 0 17572 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_191
timestamp 1644511149
transform 1 0 18676 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_21_203
timestamp 1644511149
transform 1 0 19780 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_208
timestamp 1644511149
transform 1 0 20240 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_212
timestamp 1644511149
transform 1 0 20608 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_220
timestamp 1644511149
transform 1 0 21344 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_234
timestamp 1644511149
transform 1 0 22632 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_238
timestamp 1644511149
transform 1 0 23000 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_244
timestamp 1644511149
transform 1 0 23552 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_252
timestamp 1644511149
transform 1 0 24288 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_257
timestamp 1644511149
transform 1 0 24748 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_263
timestamp 1644511149
transform 1 0 25300 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_267
timestamp 1644511149
transform 1 0 25668 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_270
timestamp 1644511149
transform 1 0 25944 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_278
timestamp 1644511149
transform 1 0 26680 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_21_281
timestamp 1644511149
transform 1 0 26956 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_289
timestamp 1644511149
transform 1 0 27692 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_296
timestamp 1644511149
transform 1 0 28336 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_308
timestamp 1644511149
transform 1 0 29440 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_320
timestamp 1644511149
transform 1 0 30544 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_326
timestamp 1644511149
transform 1 0 31096 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_332
timestamp 1644511149
transform 1 0 31648 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_337
timestamp 1644511149
transform 1 0 32108 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_346
timestamp 1644511149
transform 1 0 32936 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_21_352
timestamp 1644511149
transform 1 0 33488 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_21_376
timestamp 1644511149
transform 1 0 35696 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_21_386
timestamp 1644511149
transform 1 0 36616 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_21_397
timestamp 1644511149
transform 1 0 37628 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_408
timestamp 1644511149
transform 1 0 38640 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_420
timestamp 1644511149
transform 1 0 39744 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_432
timestamp 1644511149
transform 1 0 40848 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_444
timestamp 1644511149
transform 1 0 41952 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_449
timestamp 1644511149
transform 1 0 42412 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_21_461
timestamp 1644511149
transform 1 0 43516 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_469
timestamp 1644511149
transform 1 0 44252 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_481
timestamp 1644511149
transform 1 0 45356 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_493
timestamp 1644511149
transform 1 0 46460 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_501
timestamp 1644511149
transform 1 0 47196 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_21_505
timestamp 1644511149
transform 1 0 47564 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_21_517
timestamp 1644511149
transform 1 0 48668 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_21_529
timestamp 1644511149
transform 1 0 49772 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_21_535
timestamp 1644511149
transform 1 0 50324 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_21_538
timestamp 1644511149
transform 1 0 50600 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_21_550
timestamp 1644511149
transform 1 0 51704 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_558
timestamp 1644511149
transform 1 0 52440 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_21_574
timestamp 1644511149
transform 1 0 53912 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_21_586
timestamp 1644511149
transform 1 0 55016 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_592
timestamp 1644511149
transform 1 0 55568 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_21_600
timestamp 1644511149
transform 1 0 56304 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_21_607
timestamp 1644511149
transform 1 0 56948 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_615
timestamp 1644511149
transform 1 0 57684 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_620
timestamp 1644511149
transform 1 0 58144 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_624
timestamp 1644511149
transform 1 0 58512 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_6
timestamp 1644511149
transform 1 0 1656 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_12
timestamp 1644511149
transform 1 0 2208 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_24
timestamp 1644511149
transform 1 0 3312 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_34
timestamp 1644511149
transform 1 0 4232 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_40
timestamp 1644511149
transform 1 0 4784 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_52
timestamp 1644511149
transform 1 0 5888 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_60
timestamp 1644511149
transform 1 0 6624 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_65
timestamp 1644511149
transform 1 0 7084 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_71
timestamp 1644511149
transform 1 0 7636 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_83
timestamp 1644511149
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_85
timestamp 1644511149
transform 1 0 8924 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_22_95
timestamp 1644511149
transform 1 0 9844 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_22_105
timestamp 1644511149
transform 1 0 10764 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_22_117
timestamp 1644511149
transform 1 0 11868 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_122
timestamp 1644511149
transform 1 0 12328 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_22_132
timestamp 1644511149
transform 1 0 13248 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_22_141
timestamp 1644511149
transform 1 0 14076 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_149
timestamp 1644511149
transform 1 0 14812 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_152
timestamp 1644511149
transform 1 0 15088 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_158
timestamp 1644511149
transform 1 0 15640 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_166
timestamp 1644511149
transform 1 0 16376 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_179
timestamp 1644511149
transform 1 0 17572 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_191
timestamp 1644511149
transform 1 0 18676 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_195
timestamp 1644511149
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_197
timestamp 1644511149
transform 1 0 19228 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_203
timestamp 1644511149
transform 1 0 19780 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_211
timestamp 1644511149
transform 1 0 20516 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_219
timestamp 1644511149
transform 1 0 21252 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_227
timestamp 1644511149
transform 1 0 21988 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_233
timestamp 1644511149
transform 1 0 22540 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_241
timestamp 1644511149
transform 1 0 23276 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_22_246
timestamp 1644511149
transform 1 0 23736 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_253
timestamp 1644511149
transform 1 0 24380 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_261
timestamp 1644511149
transform 1 0 25116 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_22_273
timestamp 1644511149
transform 1 0 26220 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_281
timestamp 1644511149
transform 1 0 26956 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_22_286
timestamp 1644511149
transform 1 0 27416 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_22_299
timestamp 1644511149
transform 1 0 28612 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_307
timestamp 1644511149
transform 1 0 29348 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_309
timestamp 1644511149
transform 1 0 29532 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_22_317
timestamp 1644511149
transform 1 0 30268 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_22_323
timestamp 1644511149
transform 1 0 30820 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_326
timestamp 1644511149
transform 1 0 31096 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_332
timestamp 1644511149
transform 1 0 31648 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_342
timestamp 1644511149
transform 1 0 32568 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_346
timestamp 1644511149
transform 1 0 32936 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_353
timestamp 1644511149
transform 1 0 33580 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_359
timestamp 1644511149
transform 1 0 34132 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_363
timestamp 1644511149
transform 1 0 34500 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_387
timestamp 1644511149
transform 1 0 36708 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_395
timestamp 1644511149
transform 1 0 37444 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_406
timestamp 1644511149
transform 1 0 38456 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_414
timestamp 1644511149
transform 1 0 39192 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_22_421
timestamp 1644511149
transform 1 0 39836 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_425
timestamp 1644511149
transform 1 0 40204 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_436
timestamp 1644511149
transform 1 0 41216 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_448
timestamp 1644511149
transform 1 0 42320 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_22_460
timestamp 1644511149
transform 1 0 43424 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_471
timestamp 1644511149
transform 1 0 44436 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_475
timestamp 1644511149
transform 1 0 44804 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_477
timestamp 1644511149
transform 1 0 44988 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_485
timestamp 1644511149
transform 1 0 45724 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_22_492
timestamp 1644511149
transform 1 0 46368 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_504
timestamp 1644511149
transform 1 0 47472 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_516
timestamp 1644511149
transform 1 0 48576 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_22_528
timestamp 1644511149
transform 1 0 49680 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_537
timestamp 1644511149
transform 1 0 50508 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_22_549
timestamp 1644511149
transform 1 0 51612 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_22_561
timestamp 1644511149
transform 1 0 52716 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_564
timestamp 1644511149
transform 1 0 52992 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_22_573
timestamp 1644511149
transform 1 0 53820 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_22_584
timestamp 1644511149
transform 1 0 54832 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_589
timestamp 1644511149
transform 1 0 55292 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_22_606
timestamp 1644511149
transform 1 0 56856 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_22_614
timestamp 1644511149
transform 1 0 57592 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_22_621
timestamp 1644511149
transform 1 0 58236 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_3
timestamp 1644511149
transform 1 0 1380 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_9
timestamp 1644511149
transform 1 0 1932 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_12
timestamp 1644511149
transform 1 0 2208 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_23
timestamp 1644511149
transform 1 0 3220 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_35
timestamp 1644511149
transform 1 0 4324 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_41
timestamp 1644511149
transform 1 0 4876 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_49
timestamp 1644511149
transform 1 0 5612 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_52
timestamp 1644511149
transform 1 0 5888 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_64
timestamp 1644511149
transform 1 0 6992 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_74
timestamp 1644511149
transform 1 0 7912 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_80
timestamp 1644511149
transform 1 0 8464 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_91
timestamp 1644511149
transform 1 0 9476 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_100
timestamp 1644511149
transform 1 0 10304 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_108
timestamp 1644511149
transform 1 0 11040 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_118
timestamp 1644511149
transform 1 0 11960 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_126
timestamp 1644511149
transform 1 0 12696 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_141
timestamp 1644511149
transform 1 0 14076 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_150
timestamp 1644511149
transform 1 0 14904 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_156
timestamp 1644511149
transform 1 0 15456 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_164
timestamp 1644511149
transform 1 0 16192 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_182
timestamp 1644511149
transform 1 0 17848 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_194
timestamp 1644511149
transform 1 0 18952 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_202
timestamp 1644511149
transform 1 0 19688 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_215
timestamp 1644511149
transform 1 0 20884 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_223
timestamp 1644511149
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_225
timestamp 1644511149
transform 1 0 21804 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_23_237
timestamp 1644511149
transform 1 0 22908 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_245
timestamp 1644511149
transform 1 0 23644 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_258
timestamp 1644511149
transform 1 0 24840 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_266
timestamp 1644511149
transform 1 0 25576 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_23_274
timestamp 1644511149
transform 1 0 26312 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_284
timestamp 1644511149
transform 1 0 27232 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_290
timestamp 1644511149
transform 1 0 27784 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_305
timestamp 1644511149
transform 1 0 29164 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_316
timestamp 1644511149
transform 1 0 30176 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_327
timestamp 1644511149
transform 1 0 31188 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_23_335
timestamp 1644511149
transform 1 0 31924 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_344
timestamp 1644511149
transform 1 0 32752 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_357
timestamp 1644511149
transform 1 0 33948 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_364
timestamp 1644511149
transform 1 0 34592 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_370
timestamp 1644511149
transform 1 0 35144 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_382
timestamp 1644511149
transform 1 0 36248 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_23_390
timestamp 1644511149
transform 1 0 36984 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_23_393
timestamp 1644511149
transform 1 0 37260 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_23_401
timestamp 1644511149
transform 1 0 37996 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_407
timestamp 1644511149
transform 1 0 38548 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_413
timestamp 1644511149
transform 1 0 39100 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_425
timestamp 1644511149
transform 1 0 40204 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_429
timestamp 1644511149
transform 1 0 40572 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_23_434
timestamp 1644511149
transform 1 0 41032 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_446
timestamp 1644511149
transform 1 0 42136 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_23_449
timestamp 1644511149
transform 1 0 42412 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_461
timestamp 1644511149
transform 1 0 43516 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_475
timestamp 1644511149
transform 1 0 44804 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_23_483
timestamp 1644511149
transform 1 0 45540 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_23_496
timestamp 1644511149
transform 1 0 46736 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_23_505
timestamp 1644511149
transform 1 0 47564 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_23_521
timestamp 1644511149
transform 1 0 49036 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_531
timestamp 1644511149
transform 1 0 49956 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_540
timestamp 1644511149
transform 1 0 50784 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_23_552
timestamp 1644511149
transform 1 0 51888 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_23_568
timestamp 1644511149
transform 1 0 53360 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_23_579
timestamp 1644511149
transform 1 0 54372 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_23_591
timestamp 1644511149
transform 1 0 55476 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_23_603
timestamp 1644511149
transform 1 0 56580 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_23_608
timestamp 1644511149
transform 1 0 57040 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_23_617
timestamp 1644511149
transform 1 0 57868 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_3
timestamp 1644511149
transform 1 0 1380 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_15
timestamp 1644511149
transform 1 0 2484 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_23
timestamp 1644511149
transform 1 0 3220 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_27
timestamp 1644511149
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_24_32
timestamp 1644511149
transform 1 0 4048 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_44
timestamp 1644511149
transform 1 0 5152 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_56
timestamp 1644511149
transform 1 0 6256 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_24_75
timestamp 1644511149
transform 1 0 8004 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_83
timestamp 1644511149
transform 1 0 8740 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_87
timestamp 1644511149
transform 1 0 9108 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_99
timestamp 1644511149
transform 1 0 10212 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_106
timestamp 1644511149
transform 1 0 10856 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_112
timestamp 1644511149
transform 1 0 11408 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_118
timestamp 1644511149
transform 1 0 11960 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_130
timestamp 1644511149
transform 1 0 13064 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_136
timestamp 1644511149
transform 1 0 13616 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_146
timestamp 1644511149
transform 1 0 14536 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_162
timestamp 1644511149
transform 1 0 16008 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_174
timestamp 1644511149
transform 1 0 17112 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_24_186
timestamp 1644511149
transform 1 0 18216 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_194
timestamp 1644511149
transform 1 0 18952 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_204
timestamp 1644511149
transform 1 0 19872 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_24_212
timestamp 1644511149
transform 1 0 20608 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_24_222
timestamp 1644511149
transform 1 0 21528 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_234
timestamp 1644511149
transform 1 0 22632 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_243
timestamp 1644511149
transform 1 0 23460 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_251
timestamp 1644511149
transform 1 0 24196 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_260
timestamp 1644511149
transform 1 0 25024 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_268
timestamp 1644511149
transform 1 0 25760 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_274
timestamp 1644511149
transform 1 0 26312 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_280
timestamp 1644511149
transform 1 0 26864 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_292
timestamp 1644511149
transform 1 0 27968 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_304
timestamp 1644511149
transform 1 0 29072 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_24_309
timestamp 1644511149
transform 1 0 29532 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_314
timestamp 1644511149
transform 1 0 29992 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_24_322
timestamp 1644511149
transform 1 0 30728 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_327
timestamp 1644511149
transform 1 0 31188 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_333
timestamp 1644511149
transform 1 0 31740 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_342
timestamp 1644511149
transform 1 0 32568 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_348
timestamp 1644511149
transform 1 0 33120 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_354
timestamp 1644511149
transform 1 0 33672 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_360
timestamp 1644511149
transform 1 0 34224 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_365
timestamp 1644511149
transform 1 0 34684 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_377
timestamp 1644511149
transform 1 0 35788 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_389
timestamp 1644511149
transform 1 0 36892 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_401
timestamp 1644511149
transform 1 0 37996 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_24_413
timestamp 1644511149
transform 1 0 39100 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_24_419
timestamp 1644511149
transform 1 0 39652 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_423
timestamp 1644511149
transform 1 0 40020 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_434
timestamp 1644511149
transform 1 0 41032 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_442
timestamp 1644511149
transform 1 0 41768 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_446
timestamp 1644511149
transform 1 0 42136 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_24_456
timestamp 1644511149
transform 1 0 43056 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_464
timestamp 1644511149
transform 1 0 43792 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_470
timestamp 1644511149
transform 1 0 44344 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_24_477
timestamp 1644511149
transform 1 0 44988 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_489
timestamp 1644511149
transform 1 0 46092 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_497
timestamp 1644511149
transform 1 0 46828 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_508
timestamp 1644511149
transform 1 0 47840 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_520
timestamp 1644511149
transform 1 0 48944 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_537
timestamp 1644511149
transform 1 0 50508 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_24_549
timestamp 1644511149
transform 1 0 51612 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_566
timestamp 1644511149
transform 1 0 53176 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_572
timestamp 1644511149
transform 1 0 53728 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_24_584
timestamp 1644511149
transform 1 0 54832 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_589
timestamp 1644511149
transform 1 0 55292 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_24_601
timestamp 1644511149
transform 1 0 56396 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_24_616
timestamp 1644511149
transform 1 0 57776 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_24_624
timestamp 1644511149
transform 1 0 58512 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_25_3
timestamp 1644511149
transform 1 0 1380 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_8
timestamp 1644511149
transform 1 0 1840 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_19
timestamp 1644511149
transform 1 0 2852 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_29
timestamp 1644511149
transform 1 0 3772 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_41
timestamp 1644511149
transform 1 0 4876 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_53
timestamp 1644511149
transform 1 0 5980 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_25_57
timestamp 1644511149
transform 1 0 6348 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_71
timestamp 1644511149
transform 1 0 7636 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_79
timestamp 1644511149
transform 1 0 8372 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_85
timestamp 1644511149
transform 1 0 8924 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_92
timestamp 1644511149
transform 1 0 9568 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_105
timestamp 1644511149
transform 1 0 10764 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_111
timestamp 1644511149
transform 1 0 11316 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_113
timestamp 1644511149
transform 1 0 11500 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_25_125
timestamp 1644511149
transform 1 0 12604 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_25_131
timestamp 1644511149
transform 1 0 13156 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_137
timestamp 1644511149
transform 1 0 13708 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_141
timestamp 1644511149
transform 1 0 14076 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_146
timestamp 1644511149
transform 1 0 14536 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_25_154
timestamp 1644511149
transform 1 0 15272 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_160
timestamp 1644511149
transform 1 0 15824 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_164
timestamp 1644511149
transform 1 0 16192 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_169
timestamp 1644511149
transform 1 0 16652 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_177
timestamp 1644511149
transform 1 0 17388 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_189
timestamp 1644511149
transform 1 0 18492 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_197
timestamp 1644511149
transform 1 0 19228 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_210
timestamp 1644511149
transform 1 0 20424 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_222
timestamp 1644511149
transform 1 0 21528 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_25_225
timestamp 1644511149
transform 1 0 21804 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_231
timestamp 1644511149
transform 1 0 22356 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_234
timestamp 1644511149
transform 1 0 22632 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_247
timestamp 1644511149
transform 1 0 23828 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_253
timestamp 1644511149
transform 1 0 24380 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_259
timestamp 1644511149
transform 1 0 24932 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_25_269
timestamp 1644511149
transform 1 0 25852 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_275
timestamp 1644511149
transform 1 0 26404 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_279
timestamp 1644511149
transform 1 0 26772 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_25_281
timestamp 1644511149
transform 1 0 26956 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_290
timestamp 1644511149
transform 1 0 27784 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_298
timestamp 1644511149
transform 1 0 28520 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_306
timestamp 1644511149
transform 1 0 29256 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_25_320
timestamp 1644511149
transform 1 0 30544 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_25_332
timestamp 1644511149
transform 1 0 31648 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_337
timestamp 1644511149
transform 1 0 32108 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_343
timestamp 1644511149
transform 1 0 32660 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_360
timestamp 1644511149
transform 1 0 34224 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_366
timestamp 1644511149
transform 1 0 34776 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_25_378
timestamp 1644511149
transform 1 0 35880 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_387
timestamp 1644511149
transform 1 0 36708 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_25_391
timestamp 1644511149
transform 1 0 37076 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_393
timestamp 1644511149
transform 1 0 37260 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_418
timestamp 1644511149
transform 1 0 39560 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_430
timestamp 1644511149
transform 1 0 40664 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_442
timestamp 1644511149
transform 1 0 41768 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_25_449
timestamp 1644511149
transform 1 0 42412 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_463
timestamp 1644511149
transform 1 0 43700 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_25_474
timestamp 1644511149
transform 1 0 44712 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_486
timestamp 1644511149
transform 1 0 45816 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_498
timestamp 1644511149
transform 1 0 46920 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_25_505
timestamp 1644511149
transform 1 0 47564 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_517
timestamp 1644511149
transform 1 0 48668 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_529
timestamp 1644511149
transform 1 0 49772 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_541
timestamp 1644511149
transform 1 0 50876 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_25_553
timestamp 1644511149
transform 1 0 51980 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_559
timestamp 1644511149
transform 1 0 52532 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_25_565
timestamp 1644511149
transform 1 0 53084 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_25_577
timestamp 1644511149
transform 1 0 54188 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_25_589
timestamp 1644511149
transform 1 0 55292 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_597
timestamp 1644511149
transform 1 0 56028 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_25_606
timestamp 1644511149
transform 1 0 56856 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_25_614
timestamp 1644511149
transform 1 0 57592 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_25_617
timestamp 1644511149
transform 1 0 57868 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_25_621
timestamp 1644511149
transform 1 0 58236 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_3
timestamp 1644511149
transform 1 0 1380 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_11
timestamp 1644511149
transform 1 0 2116 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_17
timestamp 1644511149
transform 1 0 2668 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_24
timestamp 1644511149
transform 1 0 3312 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_29
timestamp 1644511149
transform 1 0 3772 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_52
timestamp 1644511149
transform 1 0 5888 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_64
timestamp 1644511149
transform 1 0 6992 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_68
timestamp 1644511149
transform 1 0 7360 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_75
timestamp 1644511149
transform 1 0 8004 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_83
timestamp 1644511149
transform 1 0 8740 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_26_85
timestamp 1644511149
transform 1 0 8924 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_26_92
timestamp 1644511149
transform 1 0 9568 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_98
timestamp 1644511149
transform 1 0 10120 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_105
timestamp 1644511149
transform 1 0 10764 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_119
timestamp 1644511149
transform 1 0 12052 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_129
timestamp 1644511149
transform 1 0 12972 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_133
timestamp 1644511149
transform 1 0 13340 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_136
timestamp 1644511149
transform 1 0 13616 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_141
timestamp 1644511149
transform 1 0 14076 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_149
timestamp 1644511149
transform 1 0 14812 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_153
timestamp 1644511149
transform 1 0 15180 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_161
timestamp 1644511149
transform 1 0 15916 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_167
timestamp 1644511149
transform 1 0 16468 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_173
timestamp 1644511149
transform 1 0 17020 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_26_185
timestamp 1644511149
transform 1 0 18124 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_193
timestamp 1644511149
transform 1 0 18860 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_197
timestamp 1644511149
transform 1 0 19228 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_209
timestamp 1644511149
transform 1 0 20332 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_220
timestamp 1644511149
transform 1 0 21344 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_232
timestamp 1644511149
transform 1 0 22448 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_26_248
timestamp 1644511149
transform 1 0 23920 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_259
timestamp 1644511149
transform 1 0 24932 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_267
timestamp 1644511149
transform 1 0 25668 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_271
timestamp 1644511149
transform 1 0 26036 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_283
timestamp 1644511149
transform 1 0 27140 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_26_297
timestamp 1644511149
transform 1 0 28428 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_305
timestamp 1644511149
transform 1 0 29164 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_26_309
timestamp 1644511149
transform 1 0 29532 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_312
timestamp 1644511149
transform 1 0 29808 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_26_320
timestamp 1644511149
transform 1 0 30544 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_330
timestamp 1644511149
transform 1 0 31464 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_336
timestamp 1644511149
transform 1 0 32016 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_350
timestamp 1644511149
transform 1 0 33304 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_362
timestamp 1644511149
transform 1 0 34408 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_372
timestamp 1644511149
transform 1 0 35328 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_378
timestamp 1644511149
transform 1 0 35880 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_392
timestamp 1644511149
transform 1 0 37168 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_26_404
timestamp 1644511149
transform 1 0 38272 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_26_413
timestamp 1644511149
transform 1 0 39100 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_419
timestamp 1644511149
transform 1 0 39652 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_26_421
timestamp 1644511149
transform 1 0 39836 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_433
timestamp 1644511149
transform 1 0 40940 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_26_445
timestamp 1644511149
transform 1 0 42044 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_26_450
timestamp 1644511149
transform 1 0 42504 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_458
timestamp 1644511149
transform 1 0 43240 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_462
timestamp 1644511149
transform 1 0 43608 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_467
timestamp 1644511149
transform 1 0 44068 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_475
timestamp 1644511149
transform 1 0 44804 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_477
timestamp 1644511149
transform 1 0 44988 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_26_492
timestamp 1644511149
transform 1 0 46368 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_26_501
timestamp 1644511149
transform 1 0 47196 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_26_513
timestamp 1644511149
transform 1 0 48300 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_26_525
timestamp 1644511149
transform 1 0 49404 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_531
timestamp 1644511149
transform 1 0 49956 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_535
timestamp 1644511149
transform 1 0 50324 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_26_545
timestamp 1644511149
transform 1 0 51244 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_26_556
timestamp 1644511149
transform 1 0 52256 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_26_564
timestamp 1644511149
transform 1 0 52992 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_26_572
timestamp 1644511149
transform 1 0 53728 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_26_581
timestamp 1644511149
transform 1 0 54556 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_587
timestamp 1644511149
transform 1 0 55108 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_589
timestamp 1644511149
transform 1 0 55292 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_597
timestamp 1644511149
transform 1 0 56028 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_611
timestamp 1644511149
transform 1 0 57316 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_621
timestamp 1644511149
transform 1 0 58236 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_3
timestamp 1644511149
transform 1 0 1380 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_7
timestamp 1644511149
transform 1 0 1748 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_25
timestamp 1644511149
transform 1 0 3404 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_37
timestamp 1644511149
transform 1 0 4508 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_49
timestamp 1644511149
transform 1 0 5612 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_55
timestamp 1644511149
transform 1 0 6164 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_57
timestamp 1644511149
transform 1 0 6348 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_65
timestamp 1644511149
transform 1 0 7084 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_72
timestamp 1644511149
transform 1 0 7728 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_81
timestamp 1644511149
transform 1 0 8556 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_88
timestamp 1644511149
transform 1 0 9200 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_94
timestamp 1644511149
transform 1 0 9752 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_108
timestamp 1644511149
transform 1 0 11040 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_113
timestamp 1644511149
transform 1 0 11500 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_125
timestamp 1644511149
transform 1 0 12604 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_133
timestamp 1644511149
transform 1 0 13340 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_137
timestamp 1644511149
transform 1 0 13708 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_148
timestamp 1644511149
transform 1 0 14720 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_159
timestamp 1644511149
transform 1 0 15732 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_167
timestamp 1644511149
transform 1 0 16468 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_169
timestamp 1644511149
transform 1 0 16652 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_27_181
timestamp 1644511149
transform 1 0 17756 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_27_187
timestamp 1644511149
transform 1 0 18308 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_27_199
timestamp 1644511149
transform 1 0 19412 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_207
timestamp 1644511149
transform 1 0 20148 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_214
timestamp 1644511149
transform 1 0 20792 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_220
timestamp 1644511149
transform 1 0 21344 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_225
timestamp 1644511149
transform 1 0 21804 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_237
timestamp 1644511149
transform 1 0 22908 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_243
timestamp 1644511149
transform 1 0 23460 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_248
timestamp 1644511149
transform 1 0 23920 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_27_258
timestamp 1644511149
transform 1 0 24840 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_266
timestamp 1644511149
transform 1 0 25576 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_27_273
timestamp 1644511149
transform 1 0 26220 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_279
timestamp 1644511149
transform 1 0 26772 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_281
timestamp 1644511149
transform 1 0 26956 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_27_293
timestamp 1644511149
transform 1 0 28060 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_303
timestamp 1644511149
transform 1 0 28980 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_311
timestamp 1644511149
transform 1 0 29716 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_27_316
timestamp 1644511149
transform 1 0 30176 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_324
timestamp 1644511149
transform 1 0 30912 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_332
timestamp 1644511149
transform 1 0 31648 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_337
timestamp 1644511149
transform 1 0 32108 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_345
timestamp 1644511149
transform 1 0 32844 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_356
timestamp 1644511149
transform 1 0 33856 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_362
timestamp 1644511149
transform 1 0 34408 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_27_374
timestamp 1644511149
transform 1 0 35512 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_380
timestamp 1644511149
transform 1 0 36064 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_388
timestamp 1644511149
transform 1 0 36800 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_400
timestamp 1644511149
transform 1 0 37904 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_412
timestamp 1644511149
transform 1 0 39008 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_420
timestamp 1644511149
transform 1 0 39744 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_425
timestamp 1644511149
transform 1 0 40204 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_436
timestamp 1644511149
transform 1 0 41216 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_449
timestamp 1644511149
transform 1 0 42412 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_27_461
timestamp 1644511149
transform 1 0 43516 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_473
timestamp 1644511149
transform 1 0 44620 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_479
timestamp 1644511149
transform 1 0 45172 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_27_485
timestamp 1644511149
transform 1 0 45724 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_27_497
timestamp 1644511149
transform 1 0 46828 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_503
timestamp 1644511149
transform 1 0 47380 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_505
timestamp 1644511149
transform 1 0 47564 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_516
timestamp 1644511149
transform 1 0 48576 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_525
timestamp 1644511149
transform 1 0 49404 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_533
timestamp 1644511149
transform 1 0 50140 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_541
timestamp 1644511149
transform 1 0 50876 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_27_550
timestamp 1644511149
transform 1 0 51704 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_27_558
timestamp 1644511149
transform 1 0 52440 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_565
timestamp 1644511149
transform 1 0 53084 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_27_576
timestamp 1644511149
transform 1 0 54096 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_27_588
timestamp 1644511149
transform 1 0 55200 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_27_596
timestamp 1644511149
transform 1 0 55936 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_27_612
timestamp 1644511149
transform 1 0 57408 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_27_617
timestamp 1644511149
transform 1 0 57868 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_27_621
timestamp 1644511149
transform 1 0 58236 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_3
timestamp 1644511149
transform 1 0 1380 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_28_11
timestamp 1644511149
transform 1 0 2116 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_28_19
timestamp 1644511149
transform 1 0 2852 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_27
timestamp 1644511149
transform 1 0 3588 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_29
timestamp 1644511149
transform 1 0 3772 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_41
timestamp 1644511149
transform 1 0 4876 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_47
timestamp 1644511149
transform 1 0 5428 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_56
timestamp 1644511149
transform 1 0 6256 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_67
timestamp 1644511149
transform 1 0 7268 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_76
timestamp 1644511149
transform 1 0 8096 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_28_88
timestamp 1644511149
transform 1 0 9200 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_100
timestamp 1644511149
transform 1 0 10304 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_112
timestamp 1644511149
transform 1 0 11408 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_120
timestamp 1644511149
transform 1 0 12144 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_28_129
timestamp 1644511149
transform 1 0 12972 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_137
timestamp 1644511149
transform 1 0 13708 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_28_141
timestamp 1644511149
transform 1 0 14076 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_147
timestamp 1644511149
transform 1 0 14628 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_158
timestamp 1644511149
transform 1 0 15640 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_170
timestamp 1644511149
transform 1 0 16744 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_178
timestamp 1644511149
transform 1 0 17480 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_183
timestamp 1644511149
transform 1 0 17940 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_189
timestamp 1644511149
transform 1 0 18492 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_195
timestamp 1644511149
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_28_197
timestamp 1644511149
transform 1 0 19228 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_203
timestamp 1644511149
transform 1 0 19780 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_216
timestamp 1644511149
transform 1 0 20976 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_28_224
timestamp 1644511149
transform 1 0 21712 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_229
timestamp 1644511149
transform 1 0 22172 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_237
timestamp 1644511149
transform 1 0 22908 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_248
timestamp 1644511149
transform 1 0 23920 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_260
timestamp 1644511149
transform 1 0 25024 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_270
timestamp 1644511149
transform 1 0 25944 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_276
timestamp 1644511149
transform 1 0 26496 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_289
timestamp 1644511149
transform 1 0 27692 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_297
timestamp 1644511149
transform 1 0 28428 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_303
timestamp 1644511149
transform 1 0 28980 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_307
timestamp 1644511149
transform 1 0 29348 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_309
timestamp 1644511149
transform 1 0 29532 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_317
timestamp 1644511149
transform 1 0 30268 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_28_325
timestamp 1644511149
transform 1 0 31004 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_28_335
timestamp 1644511149
transform 1 0 31924 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_343
timestamp 1644511149
transform 1 0 32660 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_352
timestamp 1644511149
transform 1 0 33488 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_358
timestamp 1644511149
transform 1 0 34040 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_28_365
timestamp 1644511149
transform 1 0 34684 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_377
timestamp 1644511149
transform 1 0 35788 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_28_384
timestamp 1644511149
transform 1 0 36432 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_390
timestamp 1644511149
transform 1 0 36984 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_402
timestamp 1644511149
transform 1 0 38088 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_414
timestamp 1644511149
transform 1 0 39192 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_421
timestamp 1644511149
transform 1 0 39836 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_427
timestamp 1644511149
transform 1 0 40388 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_438
timestamp 1644511149
transform 1 0 41400 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_450
timestamp 1644511149
transform 1 0 42504 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_28_462
timestamp 1644511149
transform 1 0 43608 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_472
timestamp 1644511149
transform 1 0 44528 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_483
timestamp 1644511149
transform 1 0 45540 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_495
timestamp 1644511149
transform 1 0 46644 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_507
timestamp 1644511149
transform 1 0 47748 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_511
timestamp 1644511149
transform 1 0 48116 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_516
timestamp 1644511149
transform 1 0 48576 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_528
timestamp 1644511149
transform 1 0 49680 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_533
timestamp 1644511149
transform 1 0 50140 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_28_545
timestamp 1644511149
transform 1 0 51244 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_28_557
timestamp 1644511149
transform 1 0 52348 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_28_565
timestamp 1644511149
transform 1 0 53084 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_28_575
timestamp 1644511149
transform 1 0 54004 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_587
timestamp 1644511149
transform 1 0 55108 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_589
timestamp 1644511149
transform 1 0 55292 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_28_601
timestamp 1644511149
transform 1 0 56396 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_609
timestamp 1644511149
transform 1 0 57132 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_28_621
timestamp 1644511149
transform 1 0 58236 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_3
timestamp 1644511149
transform 1 0 1380 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_7
timestamp 1644511149
transform 1 0 1748 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_13
timestamp 1644511149
transform 1 0 2300 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_22
timestamp 1644511149
transform 1 0 3128 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_34
timestamp 1644511149
transform 1 0 4232 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_46
timestamp 1644511149
transform 1 0 5336 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_54
timestamp 1644511149
transform 1 0 6072 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_57
timestamp 1644511149
transform 1 0 6348 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_61
timestamp 1644511149
transform 1 0 6716 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_65
timestamp 1644511149
transform 1 0 7084 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_82
timestamp 1644511149
transform 1 0 8648 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_94
timestamp 1644511149
transform 1 0 9752 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_108
timestamp 1644511149
transform 1 0 11040 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_126
timestamp 1644511149
transform 1 0 12696 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_132
timestamp 1644511149
transform 1 0 13248 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_29_144
timestamp 1644511149
transform 1 0 14352 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_152
timestamp 1644511149
transform 1 0 15088 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_160
timestamp 1644511149
transform 1 0 15824 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_29_169
timestamp 1644511149
transform 1 0 16652 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_177
timestamp 1644511149
transform 1 0 17388 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_184
timestamp 1644511149
transform 1 0 18032 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_198
timestamp 1644511149
transform 1 0 19320 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_29_212
timestamp 1644511149
transform 1 0 20608 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_225
timestamp 1644511149
transform 1 0 21804 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_239
timestamp 1644511149
transform 1 0 23092 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_247
timestamp 1644511149
transform 1 0 23828 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_251
timestamp 1644511149
transform 1 0 24196 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_260
timestamp 1644511149
transform 1 0 25024 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_29_266
timestamp 1644511149
transform 1 0 25576 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_276
timestamp 1644511149
transform 1 0 26496 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_283
timestamp 1644511149
transform 1 0 27140 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_297
timestamp 1644511149
transform 1 0 28428 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_303
timestamp 1644511149
transform 1 0 28980 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_29_308
timestamp 1644511149
transform 1 0 29440 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_314
timestamp 1644511149
transform 1 0 29992 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_324
timestamp 1644511149
transform 1 0 30912 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_332
timestamp 1644511149
transform 1 0 31648 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_29_339
timestamp 1644511149
transform 1 0 32292 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_29_347
timestamp 1644511149
transform 1 0 33028 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_359
timestamp 1644511149
transform 1 0 34132 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_365
timestamp 1644511149
transform 1 0 34684 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_377
timestamp 1644511149
transform 1 0 35788 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_29_386
timestamp 1644511149
transform 1 0 36616 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_29_397
timestamp 1644511149
transform 1 0 37628 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_403
timestamp 1644511149
transform 1 0 38180 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_417
timestamp 1644511149
transform 1 0 39468 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_425
timestamp 1644511149
transform 1 0 40204 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_29_431
timestamp 1644511149
transform 1 0 40756 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_29_443
timestamp 1644511149
transform 1 0 41860 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_447
timestamp 1644511149
transform 1 0 42228 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_449
timestamp 1644511149
transform 1 0 42412 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_461
timestamp 1644511149
transform 1 0 43516 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_486
timestamp 1644511149
transform 1 0 45816 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_498
timestamp 1644511149
transform 1 0 46920 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_29_505
timestamp 1644511149
transform 1 0 47564 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_29_517
timestamp 1644511149
transform 1 0 48668 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_29_525
timestamp 1644511149
transform 1 0 49404 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_537
timestamp 1644511149
transform 1 0 50508 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_29_549
timestamp 1644511149
transform 1 0 51612 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_29_557
timestamp 1644511149
transform 1 0 52348 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_29_561
timestamp 1644511149
transform 1 0 52716 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_565
timestamp 1644511149
transform 1 0 53084 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_29_572
timestamp 1644511149
transform 1 0 53728 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_29_584
timestamp 1644511149
transform 1 0 54832 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_29_596
timestamp 1644511149
transform 1 0 55936 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_29_602
timestamp 1644511149
transform 1 0 56488 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_606
timestamp 1644511149
transform 1 0 56856 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_29_614
timestamp 1644511149
transform 1 0 57592 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_620
timestamp 1644511149
transform 1 0 58144 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_624
timestamp 1644511149
transform 1 0 58512 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_5
timestamp 1644511149
transform 1 0 1564 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_11
timestamp 1644511149
transform 1 0 2116 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_16
timestamp 1644511149
transform 1 0 2576 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_51
timestamp 1644511149
transform 1 0 5796 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_63
timestamp 1644511149
transform 1 0 6900 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_75
timestamp 1644511149
transform 1 0 8004 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_83
timestamp 1644511149
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_85
timestamp 1644511149
transform 1 0 8924 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_97
timestamp 1644511149
transform 1 0 10028 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_100
timestamp 1644511149
transform 1 0 10304 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_111
timestamp 1644511149
transform 1 0 11316 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_117
timestamp 1644511149
transform 1 0 11868 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_129
timestamp 1644511149
transform 1 0 12972 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_133
timestamp 1644511149
transform 1 0 13340 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_136
timestamp 1644511149
transform 1 0 13616 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_30_141
timestamp 1644511149
transform 1 0 14076 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_165
timestamp 1644511149
transform 1 0 16284 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_173
timestamp 1644511149
transform 1 0 17020 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_180
timestamp 1644511149
transform 1 0 17664 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_187
timestamp 1644511149
transform 1 0 18308 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_195
timestamp 1644511149
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_202
timestamp 1644511149
transform 1 0 19688 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_208
timestamp 1644511149
transform 1 0 20240 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_220
timestamp 1644511149
transform 1 0 21344 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_30_230
timestamp 1644511149
transform 1 0 22264 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_30_242
timestamp 1644511149
transform 1 0 23368 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_248
timestamp 1644511149
transform 1 0 23920 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_256
timestamp 1644511149
transform 1 0 24656 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_262
timestamp 1644511149
transform 1 0 25208 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_279
timestamp 1644511149
transform 1 0 26772 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_289
timestamp 1644511149
transform 1 0 27692 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_297
timestamp 1644511149
transform 1 0 28428 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_301
timestamp 1644511149
transform 1 0 28796 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_304
timestamp 1644511149
transform 1 0 29072 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_316
timestamp 1644511149
transform 1 0 30176 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_324
timestamp 1644511149
transform 1 0 30912 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_328
timestamp 1644511149
transform 1 0 31280 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_335
timestamp 1644511149
transform 1 0 31924 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_30_348
timestamp 1644511149
transform 1 0 33120 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_352
timestamp 1644511149
transform 1 0 33488 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_360
timestamp 1644511149
transform 1 0 34224 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_365
timestamp 1644511149
transform 1 0 34684 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_377
timestamp 1644511149
transform 1 0 35788 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_383
timestamp 1644511149
transform 1 0 36340 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_395
timestamp 1644511149
transform 1 0 37444 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_407
timestamp 1644511149
transform 1 0 38548 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_30_419
timestamp 1644511149
transform 1 0 39652 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_421
timestamp 1644511149
transform 1 0 39836 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_30_432
timestamp 1644511149
transform 1 0 40848 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_440
timestamp 1644511149
transform 1 0 41584 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_444
timestamp 1644511149
transform 1 0 41952 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_453
timestamp 1644511149
transform 1 0 42780 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_30_465
timestamp 1644511149
transform 1 0 43884 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_473
timestamp 1644511149
transform 1 0 44620 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_477
timestamp 1644511149
transform 1 0 44988 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_30_485
timestamp 1644511149
transform 1 0 45724 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_489
timestamp 1644511149
transform 1 0 46092 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_501
timestamp 1644511149
transform 1 0 47196 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_30_513
timestamp 1644511149
transform 1 0 48300 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_30_525
timestamp 1644511149
transform 1 0 49404 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_531
timestamp 1644511149
transform 1 0 49956 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_30_541
timestamp 1644511149
transform 1 0 50876 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_553
timestamp 1644511149
transform 1 0 51980 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_562
timestamp 1644511149
transform 1 0 52808 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_30_573
timestamp 1644511149
transform 1 0 53820 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_30_585
timestamp 1644511149
transform 1 0 54924 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_589
timestamp 1644511149
transform 1 0 55292 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_30_597
timestamp 1644511149
transform 1 0 56028 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_613
timestamp 1644511149
transform 1 0 57500 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_30_620
timestamp 1644511149
transform 1 0 58144 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_624
timestamp 1644511149
transform 1 0 58512 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_9
timestamp 1644511149
transform 1 0 1932 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_35
timestamp 1644511149
transform 1 0 4324 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_45
timestamp 1644511149
transform 1 0 5244 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_51
timestamp 1644511149
transform 1 0 5796 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_55
timestamp 1644511149
transform 1 0 6164 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_57
timestamp 1644511149
transform 1 0 6348 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_31_75
timestamp 1644511149
transform 1 0 8004 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_87
timestamp 1644511149
transform 1 0 9108 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_99
timestamp 1644511149
transform 1 0 10212 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_103
timestamp 1644511149
transform 1 0 10580 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_106
timestamp 1644511149
transform 1 0 10856 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_31_113
timestamp 1644511149
transform 1 0 11500 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_31_121
timestamp 1644511149
transform 1 0 12236 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_129
timestamp 1644511149
transform 1 0 12972 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_141
timestamp 1644511149
transform 1 0 14076 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_31_162
timestamp 1644511149
transform 1 0 16008 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_31_171
timestamp 1644511149
transform 1 0 16836 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_182
timestamp 1644511149
transform 1 0 17848 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_193
timestamp 1644511149
transform 1 0 18860 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_206
timestamp 1644511149
transform 1 0 20056 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_212
timestamp 1644511149
transform 1 0 20608 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_220
timestamp 1644511149
transform 1 0 21344 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_234
timestamp 1644511149
transform 1 0 22632 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_245
timestamp 1644511149
transform 1 0 23644 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_256
timestamp 1644511149
transform 1 0 24656 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_268
timestamp 1644511149
transform 1 0 25760 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_281
timestamp 1644511149
transform 1 0 26956 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_285
timestamp 1644511149
transform 1 0 27324 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_288
timestamp 1644511149
transform 1 0 27600 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_302
timestamp 1644511149
transform 1 0 28888 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_314
timestamp 1644511149
transform 1 0 29992 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_31_326
timestamp 1644511149
transform 1 0 31096 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_332
timestamp 1644511149
transform 1 0 31648 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_344
timestamp 1644511149
transform 1 0 32752 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_31_356
timestamp 1644511149
transform 1 0 33856 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_360
timestamp 1644511149
transform 1 0 34224 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_365
timestamp 1644511149
transform 1 0 34684 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_371
timestamp 1644511149
transform 1 0 35236 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_383
timestamp 1644511149
transform 1 0 36340 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_391
timestamp 1644511149
transform 1 0 37076 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_393
timestamp 1644511149
transform 1 0 37260 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_399
timestamp 1644511149
transform 1 0 37812 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_407
timestamp 1644511149
transform 1 0 38548 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_419
timestamp 1644511149
transform 1 0 39652 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_31_431
timestamp 1644511149
transform 1 0 40756 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_439
timestamp 1644511149
transform 1 0 41492 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_31_444
timestamp 1644511149
transform 1 0 41952 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_449
timestamp 1644511149
transform 1 0 42412 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_460
timestamp 1644511149
transform 1 0 43424 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_31_469
timestamp 1644511149
transform 1 0 44252 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_31_481
timestamp 1644511149
transform 1 0 45356 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_495
timestamp 1644511149
transform 1 0 46644 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_503
timestamp 1644511149
transform 1 0 47380 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_510
timestamp 1644511149
transform 1 0 48024 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_521
timestamp 1644511149
transform 1 0 49036 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_532
timestamp 1644511149
transform 1 0 50048 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_31_542
timestamp 1644511149
transform 1 0 50968 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_552
timestamp 1644511149
transform 1 0 51888 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_31_561
timestamp 1644511149
transform 1 0 52716 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_569
timestamp 1644511149
transform 1 0 53452 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_31_578
timestamp 1644511149
transform 1 0 54280 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_590
timestamp 1644511149
transform 1 0 55384 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_31_602
timestamp 1644511149
transform 1 0 56488 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_31_610
timestamp 1644511149
transform 1 0 57224 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_31_617
timestamp 1644511149
transform 1 0 57868 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_32_3
timestamp 1644511149
transform 1 0 1380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_15
timestamp 1644511149
transform 1 0 2484 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_24
timestamp 1644511149
transform 1 0 3312 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_29
timestamp 1644511149
transform 1 0 3772 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_32_35
timestamp 1644511149
transform 1 0 4324 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_42
timestamp 1644511149
transform 1 0 4968 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_51
timestamp 1644511149
transform 1 0 5796 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_57
timestamp 1644511149
transform 1 0 6348 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_71
timestamp 1644511149
transform 1 0 7636 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_80
timestamp 1644511149
transform 1 0 8464 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_85
timestamp 1644511149
transform 1 0 8924 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_32_98
timestamp 1644511149
transform 1 0 10120 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_32_113
timestamp 1644511149
transform 1 0 11500 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_119
timestamp 1644511149
transform 1 0 12052 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_131
timestamp 1644511149
transform 1 0 13156 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_136
timestamp 1644511149
transform 1 0 13616 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_144
timestamp 1644511149
transform 1 0 14352 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_150
timestamp 1644511149
transform 1 0 14904 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_32_156
timestamp 1644511149
transform 1 0 15456 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_32_168
timestamp 1644511149
transform 1 0 16560 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_176
timestamp 1644511149
transform 1 0 17296 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_188
timestamp 1644511149
transform 1 0 18400 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_197
timestamp 1644511149
transform 1 0 19228 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_208
timestamp 1644511149
transform 1 0 20240 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_220
timestamp 1644511149
transform 1 0 21344 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_225
timestamp 1644511149
transform 1 0 21804 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_237
timestamp 1644511149
transform 1 0 22908 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_32_243
timestamp 1644511149
transform 1 0 23460 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_251
timestamp 1644511149
transform 1 0 24196 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_253
timestamp 1644511149
transform 1 0 24380 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_265
timestamp 1644511149
transform 1 0 25484 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_279
timestamp 1644511149
transform 1 0 26772 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_287
timestamp 1644511149
transform 1 0 27508 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_298
timestamp 1644511149
transform 1 0 28520 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_304
timestamp 1644511149
transform 1 0 29072 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_309
timestamp 1644511149
transform 1 0 29532 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_321
timestamp 1644511149
transform 1 0 30636 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_324
timestamp 1644511149
transform 1 0 30912 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_336
timestamp 1644511149
transform 1 0 32016 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_341
timestamp 1644511149
transform 1 0 32476 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_32_353
timestamp 1644511149
transform 1 0 33580 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_360
timestamp 1644511149
transform 1 0 34224 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_369
timestamp 1644511149
transform 1 0 35052 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_32_377
timestamp 1644511149
transform 1 0 35788 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_391
timestamp 1644511149
transform 1 0 37076 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_403
timestamp 1644511149
transform 1 0 38180 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_409
timestamp 1644511149
transform 1 0 38732 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_32_417
timestamp 1644511149
transform 1 0 39468 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_32_421
timestamp 1644511149
transform 1 0 39836 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_433
timestamp 1644511149
transform 1 0 40940 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_445
timestamp 1644511149
transform 1 0 42044 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_451
timestamp 1644511149
transform 1 0 42596 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_460
timestamp 1644511149
transform 1 0 43424 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_472
timestamp 1644511149
transform 1 0 44528 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_477
timestamp 1644511149
transform 1 0 44988 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_489
timestamp 1644511149
transform 1 0 46092 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_506
timestamp 1644511149
transform 1 0 47656 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_518
timestamp 1644511149
transform 1 0 48760 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_32_530
timestamp 1644511149
transform 1 0 49864 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_32_540
timestamp 1644511149
transform 1 0 50784 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_32_552
timestamp 1644511149
transform 1 0 51888 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_564
timestamp 1644511149
transform 1 0 52992 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_568
timestamp 1644511149
transform 1 0 53360 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_575
timestamp 1644511149
transform 1 0 54004 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_583
timestamp 1644511149
transform 1 0 54740 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_587
timestamp 1644511149
transform 1 0 55108 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_589
timestamp 1644511149
transform 1 0 55292 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_32_601
timestamp 1644511149
transform 1 0 56396 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_32_609
timestamp 1644511149
transform 1 0 57132 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_32_621
timestamp 1644511149
transform 1 0 58236 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_3
timestamp 1644511149
transform 1 0 1380 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_33_16
timestamp 1644511149
transform 1 0 2576 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_22
timestamp 1644511149
transform 1 0 3128 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_33_37
timestamp 1644511149
transform 1 0 4508 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_43
timestamp 1644511149
transform 1 0 5060 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_46
timestamp 1644511149
transform 1 0 5336 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_54
timestamp 1644511149
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_57
timestamp 1644511149
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_69
timestamp 1644511149
transform 1 0 7452 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_77
timestamp 1644511149
transform 1 0 8188 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_89
timestamp 1644511149
transform 1 0 9292 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_102
timestamp 1644511149
transform 1 0 10488 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_110
timestamp 1644511149
transform 1 0 11224 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_113
timestamp 1644511149
transform 1 0 11500 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_125
timestamp 1644511149
transform 1 0 12604 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_129
timestamp 1644511149
transform 1 0 12972 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_138
timestamp 1644511149
transform 1 0 13800 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_146
timestamp 1644511149
transform 1 0 14536 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_149
timestamp 1644511149
transform 1 0 14812 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_157
timestamp 1644511149
transform 1 0 15548 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_160
timestamp 1644511149
transform 1 0 15824 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_169
timestamp 1644511149
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_33_181
timestamp 1644511149
transform 1 0 17756 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_185
timestamp 1644511149
transform 1 0 18124 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_192
timestamp 1644511149
transform 1 0 18768 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_196
timestamp 1644511149
transform 1 0 19136 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_201
timestamp 1644511149
transform 1 0 19596 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_209
timestamp 1644511149
transform 1 0 20332 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_221
timestamp 1644511149
transform 1 0 21436 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_227
timestamp 1644511149
transform 1 0 21988 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_239
timestamp 1644511149
transform 1 0 23092 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_33_247
timestamp 1644511149
transform 1 0 23828 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_33_251
timestamp 1644511149
transform 1 0 24196 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_33_265
timestamp 1644511149
transform 1 0 25484 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_273
timestamp 1644511149
transform 1 0 26220 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_279
timestamp 1644511149
transform 1 0 26772 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_283
timestamp 1644511149
transform 1 0 27140 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_287
timestamp 1644511149
transform 1 0 27508 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_292
timestamp 1644511149
transform 1 0 27968 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_300
timestamp 1644511149
transform 1 0 28704 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_306
timestamp 1644511149
transform 1 0 29256 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_314
timestamp 1644511149
transform 1 0 29992 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_320
timestamp 1644511149
transform 1 0 30544 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_33_328
timestamp 1644511149
transform 1 0 31280 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_33_337
timestamp 1644511149
transform 1 0 32108 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_345
timestamp 1644511149
transform 1 0 32844 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_348
timestamp 1644511149
transform 1 0 33120 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_358
timestamp 1644511149
transform 1 0 34040 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_369
timestamp 1644511149
transform 1 0 35052 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_33_381
timestamp 1644511149
transform 1 0 36156 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_33_389
timestamp 1644511149
transform 1 0 36892 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_33_393
timestamp 1644511149
transform 1 0 37260 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_401
timestamp 1644511149
transform 1 0 37996 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_415
timestamp 1644511149
transform 1 0 39284 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_419
timestamp 1644511149
transform 1 0 39652 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_422
timestamp 1644511149
transform 1 0 39928 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_33_433
timestamp 1644511149
transform 1 0 40940 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_445
timestamp 1644511149
transform 1 0 42044 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_455
timestamp 1644511149
transform 1 0 42964 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_464
timestamp 1644511149
transform 1 0 43792 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_33_470
timestamp 1644511149
transform 1 0 44344 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_33_480
timestamp 1644511149
transform 1 0 45264 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_492
timestamp 1644511149
transform 1 0 46368 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_505
timestamp 1644511149
transform 1 0 47564 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_517
timestamp 1644511149
transform 1 0 48668 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_529
timestamp 1644511149
transform 1 0 49772 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_33_541
timestamp 1644511149
transform 1 0 50876 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_33_552
timestamp 1644511149
transform 1 0 51888 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_33_561
timestamp 1644511149
transform 1 0 52716 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_573
timestamp 1644511149
transform 1 0 53820 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_585
timestamp 1644511149
transform 1 0 54924 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_33_597
timestamp 1644511149
transform 1 0 56028 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_603
timestamp 1644511149
transform 1 0 56580 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_611
timestamp 1644511149
transform 1 0 57316 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_615
timestamp 1644511149
transform 1 0 57684 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_33_617
timestamp 1644511149
transform 1 0 57868 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_33_621
timestamp 1644511149
transform 1 0 58236 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_5
timestamp 1644511149
transform 1 0 1564 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_34_13
timestamp 1644511149
transform 1 0 2300 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_34_20
timestamp 1644511149
transform 1 0 2944 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_34_29
timestamp 1644511149
transform 1 0 3772 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_41
timestamp 1644511149
transform 1 0 4876 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_53
timestamp 1644511149
transform 1 0 5980 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_57
timestamp 1644511149
transform 1 0 6348 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_66
timestamp 1644511149
transform 1 0 7176 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_78
timestamp 1644511149
transform 1 0 8280 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_85
timestamp 1644511149
transform 1 0 8924 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_89
timestamp 1644511149
transform 1 0 9292 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_92
timestamp 1644511149
transform 1 0 9568 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_100
timestamp 1644511149
transform 1 0 10304 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_108
timestamp 1644511149
transform 1 0 11040 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_34_120
timestamp 1644511149
transform 1 0 12144 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_128
timestamp 1644511149
transform 1 0 12880 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_133
timestamp 1644511149
transform 1 0 13340 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_139
timestamp 1644511149
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_143
timestamp 1644511149
transform 1 0 14260 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_156
timestamp 1644511149
transform 1 0 15456 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_169
timestamp 1644511149
transform 1 0 16652 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_175
timestamp 1644511149
transform 1 0 17204 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_183
timestamp 1644511149
transform 1 0 17940 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_192
timestamp 1644511149
transform 1 0 18768 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_206
timestamp 1644511149
transform 1 0 20056 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_210
timestamp 1644511149
transform 1 0 20424 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_218
timestamp 1644511149
transform 1 0 21160 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_230
timestamp 1644511149
transform 1 0 22264 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_242
timestamp 1644511149
transform 1 0 23368 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_248
timestamp 1644511149
transform 1 0 23920 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_263
timestamp 1644511149
transform 1 0 25300 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_271
timestamp 1644511149
transform 1 0 26036 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_275
timestamp 1644511149
transform 1 0 26404 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_280
timestamp 1644511149
transform 1 0 26864 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_291
timestamp 1644511149
transform 1 0 27876 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_297
timestamp 1644511149
transform 1 0 28428 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_301
timestamp 1644511149
transform 1 0 28796 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_304
timestamp 1644511149
transform 1 0 29072 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_34_316
timestamp 1644511149
transform 1 0 30176 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_327
timestamp 1644511149
transform 1 0 31188 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_338
timestamp 1644511149
transform 1 0 32200 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_348
timestamp 1644511149
transform 1 0 33120 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_34_360
timestamp 1644511149
transform 1 0 34224 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_369
timestamp 1644511149
transform 1 0 35052 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_381
timestamp 1644511149
transform 1 0 36156 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_387
timestamp 1644511149
transform 1 0 36708 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_395
timestamp 1644511149
transform 1 0 37444 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_407
timestamp 1644511149
transform 1 0 38548 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_34_419
timestamp 1644511149
transform 1 0 39652 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_421
timestamp 1644511149
transform 1 0 39836 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_34_429
timestamp 1644511149
transform 1 0 40572 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_34_441
timestamp 1644511149
transform 1 0 41676 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_456
timestamp 1644511149
transform 1 0 43056 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_467
timestamp 1644511149
transform 1 0 44068 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_475
timestamp 1644511149
transform 1 0 44804 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_483
timestamp 1644511149
transform 1 0 45540 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_495
timestamp 1644511149
transform 1 0 46644 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_34_507
timestamp 1644511149
transform 1 0 47748 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_34_519
timestamp 1644511149
transform 1 0 48852 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_528
timestamp 1644511149
transform 1 0 49680 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_533
timestamp 1644511149
transform 1 0 50140 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_541
timestamp 1644511149
transform 1 0 50876 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_34_558
timestamp 1644511149
transform 1 0 52440 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_34_570
timestamp 1644511149
transform 1 0 53544 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_34_579
timestamp 1644511149
transform 1 0 54372 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_587
timestamp 1644511149
transform 1 0 55108 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_34_589
timestamp 1644511149
transform 1 0 55292 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_34_595
timestamp 1644511149
transform 1 0 55844 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_607
timestamp 1644511149
transform 1 0 56948 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_621
timestamp 1644511149
transform 1 0 58236 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_6
timestamp 1644511149
transform 1 0 1656 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_14
timestamp 1644511149
transform 1 0 2392 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_23
timestamp 1644511149
transform 1 0 3220 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_29
timestamp 1644511149
transform 1 0 3772 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_52
timestamp 1644511149
transform 1 0 5888 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_57
timestamp 1644511149
transform 1 0 6348 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_63
timestamp 1644511149
transform 1 0 6900 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_86
timestamp 1644511149
transform 1 0 9016 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_90
timestamp 1644511149
transform 1 0 9384 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_95
timestamp 1644511149
transform 1 0 9844 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_103
timestamp 1644511149
transform 1 0 10580 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_111
timestamp 1644511149
transform 1 0 11316 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_115
timestamp 1644511149
transform 1 0 11684 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_127
timestamp 1644511149
transform 1 0 12788 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_136
timestamp 1644511149
transform 1 0 13616 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_140
timestamp 1644511149
transform 1 0 13984 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_145
timestamp 1644511149
transform 1 0 14444 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_157
timestamp 1644511149
transform 1 0 15548 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_163
timestamp 1644511149
transform 1 0 16100 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_167
timestamp 1644511149
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_169
timestamp 1644511149
transform 1 0 16652 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_177
timestamp 1644511149
transform 1 0 17388 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_191
timestamp 1644511149
transform 1 0 18676 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_204
timestamp 1644511149
transform 1 0 19872 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_212
timestamp 1644511149
transform 1 0 20608 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_218
timestamp 1644511149
transform 1 0 21160 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_225
timestamp 1644511149
transform 1 0 21804 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_237
timestamp 1644511149
transform 1 0 22908 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_35_241
timestamp 1644511149
transform 1 0 23276 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_247
timestamp 1644511149
transform 1 0 23828 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_256
timestamp 1644511149
transform 1 0 24656 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_267
timestamp 1644511149
transform 1 0 25668 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_275
timestamp 1644511149
transform 1 0 26404 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_279
timestamp 1644511149
transform 1 0 26772 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_281
timestamp 1644511149
transform 1 0 26956 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_285
timestamp 1644511149
transform 1 0 27324 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_289
timestamp 1644511149
transform 1 0 27692 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_301
timestamp 1644511149
transform 1 0 28796 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_35_315
timestamp 1644511149
transform 1 0 30084 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_332
timestamp 1644511149
transform 1 0 31648 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_337
timestamp 1644511149
transform 1 0 32108 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_345
timestamp 1644511149
transform 1 0 32844 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_35_352
timestamp 1644511149
transform 1 0 33488 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_360
timestamp 1644511149
transform 1 0 34224 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_363
timestamp 1644511149
transform 1 0 34500 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_35_371
timestamp 1644511149
transform 1 0 35236 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_35_377
timestamp 1644511149
transform 1 0 35788 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_35_389
timestamp 1644511149
transform 1 0 36892 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_35_393
timestamp 1644511149
transform 1 0 37260 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_405
timestamp 1644511149
transform 1 0 38364 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_417
timestamp 1644511149
transform 1 0 39468 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_429
timestamp 1644511149
transform 1 0 40572 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_441
timestamp 1644511149
transform 1 0 41676 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_447
timestamp 1644511149
transform 1 0 42228 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_35_449
timestamp 1644511149
transform 1 0 42412 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_457
timestamp 1644511149
transform 1 0 43148 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_35_460
timestamp 1644511149
transform 1 0 43424 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_35_472
timestamp 1644511149
transform 1 0 44528 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_35_484
timestamp 1644511149
transform 1 0 45632 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_35_495
timestamp 1644511149
transform 1 0 46644 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_35_503
timestamp 1644511149
transform 1 0 47380 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_505
timestamp 1644511149
transform 1 0 47564 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_522
timestamp 1644511149
transform 1 0 49128 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_35_531
timestamp 1644511149
transform 1 0 49956 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_543
timestamp 1644511149
transform 1 0 51060 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_35_549
timestamp 1644511149
transform 1 0 51612 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_35_556
timestamp 1644511149
transform 1 0 52256 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_35_569
timestamp 1644511149
transform 1 0 53452 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_35_580
timestamp 1644511149
transform 1 0 54464 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_35_592
timestamp 1644511149
transform 1 0 55568 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_603
timestamp 1644511149
transform 1 0 56580 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_35_610
timestamp 1644511149
transform 1 0 57224 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_35_620
timestamp 1644511149
transform 1 0 58144 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_35_624
timestamp 1644511149
transform 1 0 58512 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_3
timestamp 1644511149
transform 1 0 1380 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_9
timestamp 1644511149
transform 1 0 1932 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_16
timestamp 1644511149
transform 1 0 2576 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_20
timestamp 1644511149
transform 1 0 2944 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_24
timestamp 1644511149
transform 1 0 3312 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_29
timestamp 1644511149
transform 1 0 3772 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_39
timestamp 1644511149
transform 1 0 4692 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_48
timestamp 1644511149
transform 1 0 5520 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_60
timestamp 1644511149
transform 1 0 6624 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_66
timestamp 1644511149
transform 1 0 7176 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_74
timestamp 1644511149
transform 1 0 7912 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_80
timestamp 1644511149
transform 1 0 8464 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_36_85
timestamp 1644511149
transform 1 0 8924 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_92
timestamp 1644511149
transform 1 0 9568 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_104
timestamp 1644511149
transform 1 0 10672 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_112
timestamp 1644511149
transform 1 0 11408 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_36_124
timestamp 1644511149
transform 1 0 12512 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_36_128
timestamp 1644511149
transform 1 0 12880 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_136
timestamp 1644511149
transform 1 0 13616 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_148
timestamp 1644511149
transform 1 0 14720 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_156
timestamp 1644511149
transform 1 0 15456 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_36_161
timestamp 1644511149
transform 1 0 15916 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_169
timestamp 1644511149
transform 1 0 16652 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_181
timestamp 1644511149
transform 1 0 17756 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_193
timestamp 1644511149
transform 1 0 18860 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_36_199
timestamp 1644511149
transform 1 0 19412 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_207
timestamp 1644511149
transform 1 0 20148 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_214
timestamp 1644511149
transform 1 0 20792 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_225
timestamp 1644511149
transform 1 0 21804 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_239
timestamp 1644511149
transform 1 0 23092 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_248
timestamp 1644511149
transform 1 0 23920 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_260
timestamp 1644511149
transform 1 0 25024 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_268
timestamp 1644511149
transform 1 0 25760 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_274
timestamp 1644511149
transform 1 0 26312 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_280
timestamp 1644511149
transform 1 0 26864 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_292
timestamp 1644511149
transform 1 0 27968 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_304
timestamp 1644511149
transform 1 0 29072 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_36_309
timestamp 1644511149
transform 1 0 29532 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_36_317
timestamp 1644511149
transform 1 0 30268 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_322
timestamp 1644511149
transform 1 0 30728 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_334
timestamp 1644511149
transform 1 0 31832 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_346
timestamp 1644511149
transform 1 0 32936 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_36_352
timestamp 1644511149
transform 1 0 33488 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_36_360
timestamp 1644511149
transform 1 0 34224 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_369
timestamp 1644511149
transform 1 0 35052 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_375
timestamp 1644511149
transform 1 0 35604 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_394
timestamp 1644511149
transform 1 0 37352 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_36_402
timestamp 1644511149
transform 1 0 38088 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_405
timestamp 1644511149
transform 1 0 38364 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_416
timestamp 1644511149
transform 1 0 39376 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_36_421
timestamp 1644511149
transform 1 0 39836 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_425
timestamp 1644511149
transform 1 0 40204 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_432
timestamp 1644511149
transform 1 0 40848 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_444
timestamp 1644511149
transform 1 0 41952 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_36_456
timestamp 1644511149
transform 1 0 43056 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_468
timestamp 1644511149
transform 1 0 44160 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_36_477
timestamp 1644511149
transform 1 0 44988 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_483
timestamp 1644511149
transform 1 0 45540 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_36_490
timestamp 1644511149
transform 1 0 46184 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_36_498
timestamp 1644511149
transform 1 0 46920 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_510
timestamp 1644511149
transform 1 0 48024 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_36_522
timestamp 1644511149
transform 1 0 49128 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_36_530
timestamp 1644511149
transform 1 0 49864 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_36_533
timestamp 1644511149
transform 1 0 50140 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_545
timestamp 1644511149
transform 1 0 51244 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_557
timestamp 1644511149
transform 1 0 52348 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_36_569
timestamp 1644511149
transform 1 0 53452 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_36_581
timestamp 1644511149
transform 1 0 54556 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_36_587
timestamp 1644511149
transform 1 0 55108 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_36_589
timestamp 1644511149
transform 1 0 55292 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_36_601
timestamp 1644511149
transform 1 0 56396 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_36_608
timestamp 1644511149
transform 1 0 57040 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_36_620
timestamp 1644511149
transform 1 0 58144 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_36_624
timestamp 1644511149
transform 1 0 58512 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_37_3
timestamp 1644511149
transform 1 0 1380 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_7
timestamp 1644511149
transform 1 0 1748 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_15
timestamp 1644511149
transform 1 0 2484 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_39
timestamp 1644511149
transform 1 0 4692 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_45
timestamp 1644511149
transform 1 0 5244 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_53
timestamp 1644511149
transform 1 0 5980 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_37_57
timestamp 1644511149
transform 1 0 6348 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_61
timestamp 1644511149
transform 1 0 6716 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_69
timestamp 1644511149
transform 1 0 7452 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_74
timestamp 1644511149
transform 1 0 7912 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_86
timestamp 1644511149
transform 1 0 9016 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_92
timestamp 1644511149
transform 1 0 9568 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_98
timestamp 1644511149
transform 1 0 10120 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_101
timestamp 1644511149
transform 1 0 10396 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_109
timestamp 1644511149
transform 1 0 11132 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_37_117
timestamp 1644511149
transform 1 0 11868 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_123
timestamp 1644511149
transform 1 0 12420 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_134
timestamp 1644511149
transform 1 0 13432 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_147
timestamp 1644511149
transform 1 0 14628 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_37_155
timestamp 1644511149
transform 1 0 15364 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_161
timestamp 1644511149
transform 1 0 15916 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_164
timestamp 1644511149
transform 1 0 16192 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_177
timestamp 1644511149
transform 1 0 17388 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_37_189
timestamp 1644511149
transform 1 0 18492 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_192
timestamp 1644511149
transform 1 0 18768 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_204
timestamp 1644511149
transform 1 0 19872 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_212
timestamp 1644511149
transform 1 0 20608 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_37_220
timestamp 1644511149
transform 1 0 21344 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_232
timestamp 1644511149
transform 1 0 22448 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_240
timestamp 1644511149
transform 1 0 23184 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_243
timestamp 1644511149
transform 1 0 23460 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_251
timestamp 1644511149
transform 1 0 24196 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_257
timestamp 1644511149
transform 1 0 24748 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_263
timestamp 1644511149
transform 1 0 25300 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_275
timestamp 1644511149
transform 1 0 26404 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_279
timestamp 1644511149
transform 1 0 26772 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_281
timestamp 1644511149
transform 1 0 26956 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_289
timestamp 1644511149
transform 1 0 27692 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_37_298
timestamp 1644511149
transform 1 0 28520 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_310
timestamp 1644511149
transform 1 0 29624 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_37_319
timestamp 1644511149
transform 1 0 30452 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_37_331
timestamp 1644511149
transform 1 0 31556 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_37_335
timestamp 1644511149
transform 1 0 31924 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_37_337
timestamp 1644511149
transform 1 0 32108 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_345
timestamp 1644511149
transform 1 0 32844 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_348
timestamp 1644511149
transform 1 0 33120 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_359
timestamp 1644511149
transform 1 0 34132 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_369
timestamp 1644511149
transform 1 0 35052 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_377
timestamp 1644511149
transform 1 0 35788 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_37_385
timestamp 1644511149
transform 1 0 36524 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_37_388
timestamp 1644511149
transform 1 0 36800 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_37_400
timestamp 1644511149
transform 1 0 37904 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_412
timestamp 1644511149
transform 1 0 39008 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_420
timestamp 1644511149
transform 1 0 39744 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_37_430
timestamp 1644511149
transform 1 0 40664 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_442
timestamp 1644511149
transform 1 0 41768 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_37_449
timestamp 1644511149
transform 1 0 42412 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_37_457
timestamp 1644511149
transform 1 0 43148 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_469
timestamp 1644511149
transform 1 0 44252 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_481
timestamp 1644511149
transform 1 0 45356 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_37_489
timestamp 1644511149
transform 1 0 46092 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_37_496
timestamp 1644511149
transform 1 0 46736 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_37_505
timestamp 1644511149
transform 1 0 47564 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_37_517
timestamp 1644511149
transform 1 0 48668 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_37_536
timestamp 1644511149
transform 1 0 50416 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_37_548
timestamp 1644511149
transform 1 0 51520 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_37_569
timestamp 1644511149
transform 1 0 53452 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_37_577
timestamp 1644511149
transform 1 0 54188 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_37_590
timestamp 1644511149
transform 1 0 55384 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_37_603
timestamp 1644511149
transform 1 0 56580 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_37_612
timestamp 1644511149
transform 1 0 57408 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_37_617
timestamp 1644511149
transform 1 0 57868 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_38_3
timestamp 1644511149
transform 1 0 1380 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_11
timestamp 1644511149
transform 1 0 2116 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_23
timestamp 1644511149
transform 1 0 3220 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_27
timestamp 1644511149
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_29
timestamp 1644511149
transform 1 0 3772 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_37
timestamp 1644511149
transform 1 0 4508 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_45
timestamp 1644511149
transform 1 0 5244 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_48
timestamp 1644511149
transform 1 0 5520 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_59
timestamp 1644511149
transform 1 0 6532 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_63
timestamp 1644511149
transform 1 0 6900 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_70
timestamp 1644511149
transform 1 0 7544 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_78
timestamp 1644511149
transform 1 0 8280 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_38_85
timestamp 1644511149
transform 1 0 8924 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_93
timestamp 1644511149
transform 1 0 9660 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_38_105
timestamp 1644511149
transform 1 0 10764 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_117
timestamp 1644511149
transform 1 0 11868 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_125
timestamp 1644511149
transform 1 0 12604 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_130
timestamp 1644511149
transform 1 0 13064 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_136
timestamp 1644511149
transform 1 0 13616 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_146
timestamp 1644511149
transform 1 0 14536 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_154
timestamp 1644511149
transform 1 0 15272 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_38_166
timestamp 1644511149
transform 1 0 16376 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_172
timestamp 1644511149
transform 1 0 16928 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_183
timestamp 1644511149
transform 1 0 17940 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_195
timestamp 1644511149
transform 1 0 19044 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_197
timestamp 1644511149
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_209
timestamp 1644511149
transform 1 0 20332 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_212
timestamp 1644511149
transform 1 0 20608 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_224
timestamp 1644511149
transform 1 0 21712 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_38_236
timestamp 1644511149
transform 1 0 22816 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_241
timestamp 1644511149
transform 1 0 23276 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_248
timestamp 1644511149
transform 1 0 23920 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_253
timestamp 1644511149
transform 1 0 24380 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_261
timestamp 1644511149
transform 1 0 25116 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_273
timestamp 1644511149
transform 1 0 26220 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_284
timestamp 1644511149
transform 1 0 27232 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_292
timestamp 1644511149
transform 1 0 27968 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_38_300
timestamp 1644511149
transform 1 0 28704 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_304
timestamp 1644511149
transform 1 0 29072 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_314
timestamp 1644511149
transform 1 0 29992 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_324
timestamp 1644511149
transform 1 0 30912 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_38_341
timestamp 1644511149
transform 1 0 32476 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_349
timestamp 1644511149
transform 1 0 33212 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_38_354
timestamp 1644511149
transform 1 0 33672 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_360
timestamp 1644511149
transform 1 0 34224 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_365
timestamp 1644511149
transform 1 0 34684 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_371
timestamp 1644511149
transform 1 0 35236 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_38_377
timestamp 1644511149
transform 1 0 35788 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_389
timestamp 1644511149
transform 1 0 36892 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_401
timestamp 1644511149
transform 1 0 37996 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_38_413
timestamp 1644511149
transform 1 0 39100 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_419
timestamp 1644511149
transform 1 0 39652 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_38_421
timestamp 1644511149
transform 1 0 39836 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_433
timestamp 1644511149
transform 1 0 40940 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_445
timestamp 1644511149
transform 1 0 42044 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_38_457
timestamp 1644511149
transform 1 0 43148 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_38_469
timestamp 1644511149
transform 1 0 44252 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_38_475
timestamp 1644511149
transform 1 0 44804 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_38_477
timestamp 1644511149
transform 1 0 44988 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_38_485
timestamp 1644511149
transform 1 0 45724 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_38_494
timestamp 1644511149
transform 1 0 46552 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_38_508
timestamp 1644511149
transform 1 0 47840 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_38_520
timestamp 1644511149
transform 1 0 48944 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_38_546
timestamp 1644511149
transform 1 0 51336 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_38_570
timestamp 1644511149
transform 1 0 53544 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_38_578
timestamp 1644511149
transform 1 0 54280 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_38_584
timestamp 1644511149
transform 1 0 54832 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_38_594
timestamp 1644511149
transform 1 0 55752 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_38_598
timestamp 1644511149
transform 1 0 56120 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_38_621
timestamp 1644511149
transform 1 0 58236 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_3
timestamp 1644511149
transform 1 0 1380 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_39_31
timestamp 1644511149
transform 1 0 3956 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_39_41
timestamp 1644511149
transform 1 0 4876 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_52
timestamp 1644511149
transform 1 0 5888 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_57
timestamp 1644511149
transform 1 0 6348 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_61
timestamp 1644511149
transform 1 0 6716 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_66
timestamp 1644511149
transform 1 0 7176 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_75
timestamp 1644511149
transform 1 0 8004 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_81
timestamp 1644511149
transform 1 0 8556 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_84
timestamp 1644511149
transform 1 0 8832 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_92
timestamp 1644511149
transform 1 0 9568 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_101
timestamp 1644511149
transform 1 0 10396 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_107
timestamp 1644511149
transform 1 0 10948 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_111
timestamp 1644511149
transform 1 0 11316 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_39_113
timestamp 1644511149
transform 1 0 11500 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_39_121
timestamp 1644511149
transform 1 0 12236 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_130
timestamp 1644511149
transform 1 0 13064 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_139
timestamp 1644511149
transform 1 0 13892 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_145
timestamp 1644511149
transform 1 0 14444 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_157
timestamp 1644511149
transform 1 0 15548 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_165
timestamp 1644511149
transform 1 0 16284 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_39_176
timestamp 1644511149
transform 1 0 17296 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_39_186
timestamp 1644511149
transform 1 0 18216 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_192
timestamp 1644511149
transform 1 0 18768 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_39_197
timestamp 1644511149
transform 1 0 19228 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_204
timestamp 1644511149
transform 1 0 19872 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_39_217
timestamp 1644511149
transform 1 0 21068 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_223
timestamp 1644511149
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_225
timestamp 1644511149
transform 1 0 21804 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_239
timestamp 1644511149
transform 1 0 23092 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_251
timestamp 1644511149
transform 1 0 24196 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_263
timestamp 1644511149
transform 1 0 25300 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_271
timestamp 1644511149
transform 1 0 26036 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_279
timestamp 1644511149
transform 1 0 26772 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_281
timestamp 1644511149
transform 1 0 26956 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_293
timestamp 1644511149
transform 1 0 28060 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_298
timestamp 1644511149
transform 1 0 28520 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_312
timestamp 1644511149
transform 1 0 29808 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_318
timestamp 1644511149
transform 1 0 30360 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_39_329
timestamp 1644511149
transform 1 0 31372 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_335
timestamp 1644511149
transform 1 0 31924 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_337
timestamp 1644511149
transform 1 0 32108 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_349
timestamp 1644511149
transform 1 0 33212 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_361
timestamp 1644511149
transform 1 0 34316 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_39_368
timestamp 1644511149
transform 1 0 34960 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_380
timestamp 1644511149
transform 1 0 36064 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_39_388
timestamp 1644511149
transform 1 0 36800 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_401
timestamp 1644511149
transform 1 0 37996 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_39_413
timestamp 1644511149
transform 1 0 39100 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_418
timestamp 1644511149
transform 1 0 39560 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_429
timestamp 1644511149
transform 1 0 40572 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_39_441
timestamp 1644511149
transform 1 0 41676 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_39_447
timestamp 1644511149
transform 1 0 42228 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_449
timestamp 1644511149
transform 1 0 42412 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_39_461
timestamp 1644511149
transform 1 0 43516 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_39_468
timestamp 1644511149
transform 1 0 44160 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_39_480
timestamp 1644511149
transform 1 0 45264 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_39_488
timestamp 1644511149
transform 1 0 46000 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_39_493
timestamp 1644511149
transform 1 0 46460 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_500
timestamp 1644511149
transform 1 0 47104 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_39_511
timestamp 1644511149
transform 1 0 48116 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_523
timestamp 1644511149
transform 1 0 49220 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_538
timestamp 1644511149
transform 1 0 50600 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_39_545
timestamp 1644511149
transform 1 0 51244 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_39_551
timestamp 1644511149
transform 1 0 51796 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_39_559
timestamp 1644511149
transform 1 0 52532 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_567
timestamp 1644511149
transform 1 0 53268 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_39_579
timestamp 1644511149
transform 1 0 54372 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_591
timestamp 1644511149
transform 1 0 55476 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_595
timestamp 1644511149
transform 1 0 55844 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_39_599
timestamp 1644511149
transform 1 0 56212 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_39_611
timestamp 1644511149
transform 1 0 57316 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_39_615
timestamp 1644511149
transform 1 0 57684 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_39_617
timestamp 1644511149
transform 1 0 57868 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_39_621
timestamp 1644511149
transform 1 0 58236 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_3
timestamp 1644511149
transform 1 0 1380 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_15
timestamp 1644511149
transform 1 0 2484 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_27
timestamp 1644511149
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_31
timestamp 1644511149
transform 1 0 3956 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_43
timestamp 1644511149
transform 1 0 5060 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_55
timestamp 1644511149
transform 1 0 6164 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_67
timestamp 1644511149
transform 1 0 7268 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_73
timestamp 1644511149
transform 1 0 7820 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_79
timestamp 1644511149
transform 1 0 8372 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_83
timestamp 1644511149
transform 1 0 8740 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_85
timestamp 1644511149
transform 1 0 8924 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_89
timestamp 1644511149
transform 1 0 9292 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_94
timestamp 1644511149
transform 1 0 9752 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_106
timestamp 1644511149
transform 1 0 10856 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_114
timestamp 1644511149
transform 1 0 11592 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_40_126
timestamp 1644511149
transform 1 0 12696 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_136
timestamp 1644511149
transform 1 0 13616 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_150
timestamp 1644511149
transform 1 0 14904 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_162
timestamp 1644511149
transform 1 0 16008 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_172
timestamp 1644511149
transform 1 0 16928 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_185
timestamp 1644511149
transform 1 0 18124 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_191
timestamp 1644511149
transform 1 0 18676 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_195
timestamp 1644511149
transform 1 0 19044 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_40_197
timestamp 1644511149
transform 1 0 19228 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_40_210
timestamp 1644511149
transform 1 0 20424 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_223
timestamp 1644511149
transform 1 0 21620 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_229
timestamp 1644511149
transform 1 0 22172 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_40_241
timestamp 1644511149
transform 1 0 23276 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_248
timestamp 1644511149
transform 1 0 23920 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_253
timestamp 1644511149
transform 1 0 24380 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_262
timestamp 1644511149
transform 1 0 25208 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_274
timestamp 1644511149
transform 1 0 26312 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_40_282
timestamp 1644511149
transform 1 0 27048 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_40_285
timestamp 1644511149
transform 1 0 27324 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_294
timestamp 1644511149
transform 1 0 28152 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_40_302
timestamp 1644511149
transform 1 0 28888 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_40_309
timestamp 1644511149
transform 1 0 29532 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_314
timestamp 1644511149
transform 1 0 29992 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_320
timestamp 1644511149
transform 1 0 30544 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_330
timestamp 1644511149
transform 1 0 31464 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_342
timestamp 1644511149
transform 1 0 32568 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_352
timestamp 1644511149
transform 1 0 33488 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_359
timestamp 1644511149
transform 1 0 34132 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_40_363
timestamp 1644511149
transform 1 0 34500 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_40_371
timestamp 1644511149
transform 1 0 35236 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_383
timestamp 1644511149
transform 1 0 36340 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_398
timestamp 1644511149
transform 1 0 37720 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_408
timestamp 1644511149
transform 1 0 38640 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_40_416
timestamp 1644511149
transform 1 0 39376 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_421
timestamp 1644511149
transform 1 0 39836 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_40_429
timestamp 1644511149
transform 1 0 40572 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_40_439
timestamp 1644511149
transform 1 0 41492 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_40_448
timestamp 1644511149
transform 1 0 42320 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_40_460
timestamp 1644511149
transform 1 0 43424 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_40_466
timestamp 1644511149
transform 1 0 43976 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_474
timestamp 1644511149
transform 1 0 44712 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_485
timestamp 1644511149
transform 1 0 45724 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_497
timestamp 1644511149
transform 1 0 46828 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_505
timestamp 1644511149
transform 1 0 47564 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_40_520
timestamp 1644511149
transform 1 0 48944 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_533
timestamp 1644511149
transform 1 0 50140 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_40_545
timestamp 1644511149
transform 1 0 51244 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_40_557
timestamp 1644511149
transform 1 0 52348 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_40_568
timestamp 1644511149
transform 1 0 53360 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_40_580
timestamp 1644511149
transform 1 0 54464 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_40_596
timestamp 1644511149
transform 1 0 55936 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_40_605
timestamp 1644511149
transform 1 0 56764 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_40_613
timestamp 1644511149
transform 1 0 57500 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_40_621
timestamp 1644511149
transform 1 0 58236 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_41_3
timestamp 1644511149
transform 1 0 1380 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_7
timestamp 1644511149
transform 1 0 1748 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_18
timestamp 1644511149
transform 1 0 2760 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_28
timestamp 1644511149
transform 1 0 3680 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_34
timestamp 1644511149
transform 1 0 4232 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_46
timestamp 1644511149
transform 1 0 5336 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_54
timestamp 1644511149
transform 1 0 6072 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_41_57
timestamp 1644511149
transform 1 0 6348 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_41_71
timestamp 1644511149
transform 1 0 7636 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_79
timestamp 1644511149
transform 1 0 8372 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_95
timestamp 1644511149
transform 1 0 9844 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_103
timestamp 1644511149
transform 1 0 10580 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_111
timestamp 1644511149
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_113
timestamp 1644511149
transform 1 0 11500 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_41_125
timestamp 1644511149
transform 1 0 12604 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_131
timestamp 1644511149
transform 1 0 13156 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_137
timestamp 1644511149
transform 1 0 13708 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_143
timestamp 1644511149
transform 1 0 14260 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_155
timestamp 1644511149
transform 1 0 15364 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_167
timestamp 1644511149
transform 1 0 16468 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_169
timestamp 1644511149
transform 1 0 16652 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_177
timestamp 1644511149
transform 1 0 17388 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_185
timestamp 1644511149
transform 1 0 18124 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_197
timestamp 1644511149
transform 1 0 19228 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_209
timestamp 1644511149
transform 1 0 20332 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_216
timestamp 1644511149
transform 1 0 20976 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_41_225
timestamp 1644511149
transform 1 0 21804 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_237
timestamp 1644511149
transform 1 0 22908 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_241
timestamp 1644511149
transform 1 0 23276 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_41_244
timestamp 1644511149
transform 1 0 23552 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_41_250
timestamp 1644511149
transform 1 0 24104 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_255
timestamp 1644511149
transform 1 0 24564 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_276
timestamp 1644511149
transform 1 0 26496 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_41_281
timestamp 1644511149
transform 1 0 26956 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_41_289
timestamp 1644511149
transform 1 0 27692 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_294
timestamp 1644511149
transform 1 0 28152 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_300
timestamp 1644511149
transform 1 0 28704 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_312
timestamp 1644511149
transform 1 0 29808 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_41_328
timestamp 1644511149
transform 1 0 31280 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_41_337
timestamp 1644511149
transform 1 0 32108 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_351
timestamp 1644511149
transform 1 0 33396 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_362
timestamp 1644511149
transform 1 0 34408 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_372
timestamp 1644511149
transform 1 0 35328 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_384
timestamp 1644511149
transform 1 0 36432 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_393
timestamp 1644511149
transform 1 0 37260 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_397
timestamp 1644511149
transform 1 0 37628 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_403
timestamp 1644511149
transform 1 0 38180 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_415
timestamp 1644511149
transform 1 0 39284 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_41_426
timestamp 1644511149
transform 1 0 40296 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_41_438
timestamp 1644511149
transform 1 0 41400 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_41_443
timestamp 1644511149
transform 1 0 41860 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_447
timestamp 1644511149
transform 1 0 42228 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_449
timestamp 1644511149
transform 1 0 42412 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_461
timestamp 1644511149
transform 1 0 43516 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_41_479
timestamp 1644511149
transform 1 0 45172 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_41_491
timestamp 1644511149
transform 1 0 46276 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_41_503
timestamp 1644511149
transform 1 0 47380 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_41_505
timestamp 1644511149
transform 1 0 47564 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_41_517
timestamp 1644511149
transform 1 0 48668 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_41_525
timestamp 1644511149
transform 1 0 49404 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_41_528
timestamp 1644511149
transform 1 0 49680 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_41_545
timestamp 1644511149
transform 1 0 51244 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_41_557
timestamp 1644511149
transform 1 0 52348 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_41_561
timestamp 1644511149
transform 1 0 52716 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_41_573
timestamp 1644511149
transform 1 0 53820 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_41_585
timestamp 1644511149
transform 1 0 54924 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_41_589
timestamp 1644511149
transform 1 0 55292 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_41_598
timestamp 1644511149
transform 1 0 56120 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_41_612
timestamp 1644511149
transform 1 0 57408 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_41_621
timestamp 1644511149
transform 1 0 58236 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_3
timestamp 1644511149
transform 1 0 1380 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_11
timestamp 1644511149
transform 1 0 2116 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_24
timestamp 1644511149
transform 1 0 3312 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_36
timestamp 1644511149
transform 1 0 4416 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_43
timestamp 1644511149
transform 1 0 5060 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_55
timestamp 1644511149
transform 1 0 6164 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_62
timestamp 1644511149
transform 1 0 6808 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_42_76
timestamp 1644511149
transform 1 0 8096 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_42_85
timestamp 1644511149
transform 1 0 8924 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_93
timestamp 1644511149
transform 1 0 9660 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_101
timestamp 1644511149
transform 1 0 10396 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_113
timestamp 1644511149
transform 1 0 11500 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_125
timestamp 1644511149
transform 1 0 12604 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_136
timestamp 1644511149
transform 1 0 13616 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_150
timestamp 1644511149
transform 1 0 14904 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_162
timestamp 1644511149
transform 1 0 16008 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_168
timestamp 1644511149
transform 1 0 16560 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_176
timestamp 1644511149
transform 1 0 17296 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_42_191
timestamp 1644511149
transform 1 0 18676 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_195
timestamp 1644511149
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_197
timestamp 1644511149
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_209
timestamp 1644511149
transform 1 0 20332 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_42_213
timestamp 1644511149
transform 1 0 20700 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_221
timestamp 1644511149
transform 1 0 21436 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_226
timestamp 1644511149
transform 1 0 21896 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_234
timestamp 1644511149
transform 1 0 22632 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_239
timestamp 1644511149
transform 1 0 23092 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_243
timestamp 1644511149
transform 1 0 23460 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_247
timestamp 1644511149
transform 1 0 23828 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_251
timestamp 1644511149
transform 1 0 24196 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_261
timestamp 1644511149
transform 1 0 25116 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_273
timestamp 1644511149
transform 1 0 26220 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_42_285
timestamp 1644511149
transform 1 0 27324 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_42_291
timestamp 1644511149
transform 1 0 27876 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_304
timestamp 1644511149
transform 1 0 29072 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_309
timestamp 1644511149
transform 1 0 29532 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_323
timestamp 1644511149
transform 1 0 30820 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_334
timestamp 1644511149
transform 1 0 31832 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_346
timestamp 1644511149
transform 1 0 32936 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_360
timestamp 1644511149
transform 1 0 34224 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_372
timestamp 1644511149
transform 1 0 35328 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_42_378
timestamp 1644511149
transform 1 0 35880 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_42_390
timestamp 1644511149
transform 1 0 36984 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_396
timestamp 1644511149
transform 1 0 37536 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_403
timestamp 1644511149
transform 1 0 38180 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_42_415
timestamp 1644511149
transform 1 0 39284 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_419
timestamp 1644511149
transform 1 0 39652 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_42_421
timestamp 1644511149
transform 1 0 39836 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_42_429
timestamp 1644511149
transform 1 0 40572 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_438
timestamp 1644511149
transform 1 0 41400 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_42_447
timestamp 1644511149
transform 1 0 42228 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_42_456
timestamp 1644511149
transform 1 0 43056 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_462
timestamp 1644511149
transform 1 0 43608 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_42_469
timestamp 1644511149
transform 1 0 44252 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_42_475
timestamp 1644511149
transform 1 0 44804 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_42_477
timestamp 1644511149
transform 1 0 44988 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_42_485
timestamp 1644511149
transform 1 0 45724 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_494
timestamp 1644511149
transform 1 0 46552 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_506
timestamp 1644511149
transform 1 0 47656 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_42_518
timestamp 1644511149
transform 1 0 48760 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_530
timestamp 1644511149
transform 1 0 49864 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_42_538
timestamp 1644511149
transform 1 0 50600 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_550
timestamp 1644511149
transform 1 0 51704 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_42_558
timestamp 1644511149
transform 1 0 52440 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_42_567
timestamp 1644511149
transform 1 0 53268 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_42_579
timestamp 1644511149
transform 1 0 54372 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_42_584
timestamp 1644511149
transform 1 0 54832 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_42_589
timestamp 1644511149
transform 1 0 55292 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_42_597
timestamp 1644511149
transform 1 0 56028 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_42_609
timestamp 1644511149
transform 1 0 57132 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_42_621
timestamp 1644511149
transform 1 0 58236 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_3
timestamp 1644511149
transform 1 0 1380 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_15
timestamp 1644511149
transform 1 0 2484 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_25
timestamp 1644511149
transform 1 0 3404 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_35
timestamp 1644511149
transform 1 0 4324 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_47
timestamp 1644511149
transform 1 0 5428 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_52
timestamp 1644511149
transform 1 0 5888 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_57
timestamp 1644511149
transform 1 0 6348 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_61
timestamp 1644511149
transform 1 0 6716 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_43_77
timestamp 1644511149
transform 1 0 8188 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_85
timestamp 1644511149
transform 1 0 8924 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_92
timestamp 1644511149
transform 1 0 9568 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_103
timestamp 1644511149
transform 1 0 10580 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_111
timestamp 1644511149
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_117
timestamp 1644511149
transform 1 0 11868 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_43_129
timestamp 1644511149
transform 1 0 12972 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_43_139
timestamp 1644511149
transform 1 0 13892 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_147
timestamp 1644511149
transform 1 0 14628 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_159
timestamp 1644511149
transform 1 0 15732 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_167
timestamp 1644511149
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_43_169
timestamp 1644511149
transform 1 0 16652 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_182
timestamp 1644511149
transform 1 0 17848 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_188
timestamp 1644511149
transform 1 0 18400 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_192
timestamp 1644511149
transform 1 0 18768 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_197
timestamp 1644511149
transform 1 0 19228 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_209
timestamp 1644511149
transform 1 0 20332 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_215
timestamp 1644511149
transform 1 0 20884 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_220
timestamp 1644511149
transform 1 0 21344 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_43_225
timestamp 1644511149
transform 1 0 21804 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_43_232
timestamp 1644511149
transform 1 0 22448 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_43_240
timestamp 1644511149
transform 1 0 23184 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_248
timestamp 1644511149
transform 1 0 23920 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_257
timestamp 1644511149
transform 1 0 24748 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_269
timestamp 1644511149
transform 1 0 25852 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_277
timestamp 1644511149
transform 1 0 26588 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_43_281
timestamp 1644511149
transform 1 0 26956 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_43_289
timestamp 1644511149
transform 1 0 27692 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_43_296
timestamp 1644511149
transform 1 0 28336 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_43_308
timestamp 1644511149
transform 1 0 29440 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_43_316
timestamp 1644511149
transform 1 0 30176 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_324
timestamp 1644511149
transform 1 0 30912 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_337
timestamp 1644511149
transform 1 0 32108 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_349
timestamp 1644511149
transform 1 0 33212 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_361
timestamp 1644511149
transform 1 0 34316 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_373
timestamp 1644511149
transform 1 0 35420 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_385
timestamp 1644511149
transform 1 0 36524 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_43_391
timestamp 1644511149
transform 1 0 37076 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_43_400
timestamp 1644511149
transform 1 0 37904 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_410
timestamp 1644511149
transform 1 0 38824 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_422
timestamp 1644511149
transform 1 0 39928 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_434
timestamp 1644511149
transform 1 0 41032 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_446
timestamp 1644511149
transform 1 0 42136 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_43_449
timestamp 1644511149
transform 1 0 42412 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_43_457
timestamp 1644511149
transform 1 0 43148 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_43_467
timestamp 1644511149
transform 1 0 44068 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_479
timestamp 1644511149
transform 1 0 45172 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_43_491
timestamp 1644511149
transform 1 0 46276 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_43_500
timestamp 1644511149
transform 1 0 47104 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_510
timestamp 1644511149
transform 1 0 48024 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_43_527
timestamp 1644511149
transform 1 0 49588 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_534
timestamp 1644511149
transform 1 0 50232 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_43_546
timestamp 1644511149
transform 1 0 51336 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_43_558
timestamp 1644511149
transform 1 0 52440 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_43_567
timestamp 1644511149
transform 1 0 53268 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_43_576
timestamp 1644511149
transform 1 0 54096 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_588
timestamp 1644511149
transform 1 0 55200 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_43_592
timestamp 1644511149
transform 1 0 55568 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_43_600
timestamp 1644511149
transform 1 0 56304 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_43_612
timestamp 1644511149
transform 1 0 57408 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_43_617
timestamp 1644511149
transform 1 0 57868 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_3
timestamp 1644511149
transform 1 0 1380 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_44_7
timestamp 1644511149
transform 1 0 1748 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_19
timestamp 1644511149
transform 1 0 2852 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_27
timestamp 1644511149
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_31
timestamp 1644511149
transform 1 0 3956 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_43
timestamp 1644511149
transform 1 0 5060 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_59
timestamp 1644511149
transform 1 0 6532 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_73
timestamp 1644511149
transform 1 0 7820 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_44_81
timestamp 1644511149
transform 1 0 8556 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_44_85
timestamp 1644511149
transform 1 0 8924 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_97
timestamp 1644511149
transform 1 0 10028 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_106
timestamp 1644511149
transform 1 0 10856 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_114
timestamp 1644511149
transform 1 0 11592 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_126
timestamp 1644511149
transform 1 0 12696 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_138
timestamp 1644511149
transform 1 0 13800 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_143
timestamp 1644511149
transform 1 0 14260 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_147
timestamp 1644511149
transform 1 0 14628 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_152
timestamp 1644511149
transform 1 0 15088 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_164
timestamp 1644511149
transform 1 0 16192 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_172
timestamp 1644511149
transform 1 0 16928 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_180
timestamp 1644511149
transform 1 0 17664 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_192
timestamp 1644511149
transform 1 0 18768 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_206
timestamp 1644511149
transform 1 0 20056 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_214
timestamp 1644511149
transform 1 0 20792 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_44_222
timestamp 1644511149
transform 1 0 21528 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_44_232
timestamp 1644511149
transform 1 0 22448 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_44_248
timestamp 1644511149
transform 1 0 23920 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_256
timestamp 1644511149
transform 1 0 24656 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_262
timestamp 1644511149
transform 1 0 25208 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_274
timestamp 1644511149
transform 1 0 26312 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_286
timestamp 1644511149
transform 1 0 27416 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_44_290
timestamp 1644511149
transform 1 0 27784 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_294
timestamp 1644511149
transform 1 0 28152 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_306
timestamp 1644511149
transform 1 0 29256 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_44_309
timestamp 1644511149
transform 1 0 29532 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_317
timestamp 1644511149
transform 1 0 30268 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_44_332
timestamp 1644511149
transform 1 0 31648 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_344
timestamp 1644511149
transform 1 0 32752 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_352
timestamp 1644511149
transform 1 0 33488 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_360
timestamp 1644511149
transform 1 0 34224 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_371
timestamp 1644511149
transform 1 0 35236 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_383
timestamp 1644511149
transform 1 0 36340 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_44_391
timestamp 1644511149
transform 1 0 37076 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_44_399
timestamp 1644511149
transform 1 0 37812 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_44_408
timestamp 1644511149
transform 1 0 38640 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_44_421
timestamp 1644511149
transform 1 0 39836 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_44_429
timestamp 1644511149
transform 1 0 40572 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_44_439
timestamp 1644511149
transform 1 0 41492 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_451
timestamp 1644511149
transform 1 0 42596 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_463
timestamp 1644511149
transform 1 0 43700 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_44_475
timestamp 1644511149
transform 1 0 44804 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_477
timestamp 1644511149
transform 1 0 44988 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_489
timestamp 1644511149
transform 1 0 46092 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_501
timestamp 1644511149
transform 1 0 47196 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_513
timestamp 1644511149
transform 1 0 48300 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_44_525
timestamp 1644511149
transform 1 0 49404 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_531
timestamp 1644511149
transform 1 0 49956 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_540
timestamp 1644511149
transform 1 0 50784 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_549
timestamp 1644511149
transform 1 0 51612 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_555
timestamp 1644511149
transform 1 0 52164 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_44_558
timestamp 1644511149
transform 1 0 52440 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_44_566
timestamp 1644511149
transform 1 0 53176 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_44_572
timestamp 1644511149
transform 1 0 53728 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_44_584
timestamp 1644511149
transform 1 0 54832 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_44_589
timestamp 1644511149
transform 1 0 55292 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_44_595
timestamp 1644511149
transform 1 0 55844 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_44_599
timestamp 1644511149
transform 1 0 56212 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_44_611
timestamp 1644511149
transform 1 0 57316 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_44_623
timestamp 1644511149
transform 1 0 58420 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_3
timestamp 1644511149
transform 1 0 1380 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_11
timestamp 1644511149
transform 1 0 2116 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_23
timestamp 1644511149
transform 1 0 3220 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_35
timestamp 1644511149
transform 1 0 4324 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_45
timestamp 1644511149
transform 1 0 5244 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_52
timestamp 1644511149
transform 1 0 5888 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_57
timestamp 1644511149
transform 1 0 6348 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_61
timestamp 1644511149
transform 1 0 6716 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_69
timestamp 1644511149
transform 1 0 7452 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_78
timestamp 1644511149
transform 1 0 8280 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_90
timestamp 1644511149
transform 1 0 9384 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_96
timestamp 1644511149
transform 1 0 9936 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_102
timestamp 1644511149
transform 1 0 10488 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_110
timestamp 1644511149
transform 1 0 11224 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_113
timestamp 1644511149
transform 1 0 11500 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_121
timestamp 1644511149
transform 1 0 12236 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_131
timestamp 1644511149
transform 1 0 13156 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_141
timestamp 1644511149
transform 1 0 14076 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_154
timestamp 1644511149
transform 1 0 15272 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_45_162
timestamp 1644511149
transform 1 0 16008 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_45_169
timestamp 1644511149
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_181
timestamp 1644511149
transform 1 0 17756 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_184
timestamp 1644511149
transform 1 0 18032 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_192
timestamp 1644511149
transform 1 0 18768 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_45_197
timestamp 1644511149
transform 1 0 19228 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_45_205
timestamp 1644511149
transform 1 0 19964 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_213
timestamp 1644511149
transform 1 0 20700 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_219
timestamp 1644511149
transform 1 0 21252 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_223
timestamp 1644511149
transform 1 0 21620 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_45_225
timestamp 1644511149
transform 1 0 21804 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_233
timestamp 1644511149
transform 1 0 22540 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_45_238
timestamp 1644511149
transform 1 0 23000 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_250
timestamp 1644511149
transform 1 0 24104 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_262
timestamp 1644511149
transform 1 0 25208 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_274
timestamp 1644511149
transform 1 0 26312 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_45_281
timestamp 1644511149
transform 1 0 26956 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_45_289
timestamp 1644511149
transform 1 0 27692 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_45_300
timestamp 1644511149
transform 1 0 28704 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_311
timestamp 1644511149
transform 1 0 29716 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_323
timestamp 1644511149
transform 1 0 30820 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_335
timestamp 1644511149
transform 1 0 31924 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_337
timestamp 1644511149
transform 1 0 32108 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_349
timestamp 1644511149
transform 1 0 33212 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_45_361
timestamp 1644511149
transform 1 0 34316 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_45_365
timestamp 1644511149
transform 1 0 34684 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_373
timestamp 1644511149
transform 1 0 35420 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_385
timestamp 1644511149
transform 1 0 36524 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_391
timestamp 1644511149
transform 1 0 37076 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_393
timestamp 1644511149
transform 1 0 37260 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_45_405
timestamp 1644511149
transform 1 0 38364 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_45_412
timestamp 1644511149
transform 1 0 39008 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_45_424
timestamp 1644511149
transform 1 0 40112 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_45_429
timestamp 1644511149
transform 1 0 40572 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_45_438
timestamp 1644511149
transform 1 0 41400 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_446
timestamp 1644511149
transform 1 0 42136 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_45_449
timestamp 1644511149
transform 1 0 42412 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_461
timestamp 1644511149
transform 1 0 43516 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_45_474
timestamp 1644511149
transform 1 0 44712 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_45_481
timestamp 1644511149
transform 1 0 45356 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_493
timestamp 1644511149
transform 1 0 46460 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_45_501
timestamp 1644511149
transform 1 0 47196 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_45_505
timestamp 1644511149
transform 1 0 47564 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_45_517
timestamp 1644511149
transform 1 0 48668 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_529
timestamp 1644511149
transform 1 0 49772 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_45_537
timestamp 1644511149
transform 1 0 50508 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_45_542
timestamp 1644511149
transform 1 0 50968 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_45_554
timestamp 1644511149
transform 1 0 52072 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_45_561
timestamp 1644511149
transform 1 0 52716 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_45_567
timestamp 1644511149
transform 1 0 53268 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_45_573
timestamp 1644511149
transform 1 0 53820 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_45_585
timestamp 1644511149
transform 1 0 54924 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_45_597
timestamp 1644511149
transform 1 0 56028 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_45_612
timestamp 1644511149
transform 1 0 57408 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_45_617
timestamp 1644511149
transform 1 0 57868 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_45_621
timestamp 1644511149
transform 1 0 58236 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_3
timestamp 1644511149
transform 1 0 1380 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_9
timestamp 1644511149
transform 1 0 1932 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_17
timestamp 1644511149
transform 1 0 2668 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_21
timestamp 1644511149
transform 1 0 3036 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_24
timestamp 1644511149
transform 1 0 3312 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_29
timestamp 1644511149
transform 1 0 3772 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_41
timestamp 1644511149
transform 1 0 4876 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_46_53
timestamp 1644511149
transform 1 0 5980 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_65
timestamp 1644511149
transform 1 0 7084 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_73
timestamp 1644511149
transform 1 0 7820 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_80
timestamp 1644511149
transform 1 0 8464 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_87
timestamp 1644511149
transform 1 0 9108 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_46_99
timestamp 1644511149
transform 1 0 10212 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_106
timestamp 1644511149
transform 1 0 10856 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_118
timestamp 1644511149
transform 1 0 11960 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_133
timestamp 1644511149
transform 1 0 13340 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_139
timestamp 1644511149
transform 1 0 13892 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_149
timestamp 1644511149
transform 1 0 14812 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_155
timestamp 1644511149
transform 1 0 15364 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_46_167
timestamp 1644511149
transform 1 0 16468 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_174
timestamp 1644511149
transform 1 0 17112 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_180
timestamp 1644511149
transform 1 0 17664 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_186
timestamp 1644511149
transform 1 0 18216 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_194
timestamp 1644511149
transform 1 0 18952 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_197
timestamp 1644511149
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_46_209
timestamp 1644511149
transform 1 0 20332 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_46_217
timestamp 1644511149
transform 1 0 21068 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_229
timestamp 1644511149
transform 1 0 22172 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_237
timestamp 1644511149
transform 1 0 22908 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_246
timestamp 1644511149
transform 1 0 23736 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_46_253
timestamp 1644511149
transform 1 0 24380 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_46_266
timestamp 1644511149
transform 1 0 25576 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_275
timestamp 1644511149
transform 1 0 26404 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_284
timestamp 1644511149
transform 1 0 27232 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_290
timestamp 1644511149
transform 1 0 27784 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_299
timestamp 1644511149
transform 1 0 28612 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_307
timestamp 1644511149
transform 1 0 29348 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_46_309
timestamp 1644511149
transform 1 0 29532 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_46_316
timestamp 1644511149
transform 1 0 30176 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_320
timestamp 1644511149
transform 1 0 30544 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_327
timestamp 1644511149
transform 1 0 31188 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_339
timestamp 1644511149
transform 1 0 32292 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_46_348
timestamp 1644511149
transform 1 0 33120 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_354
timestamp 1644511149
transform 1 0 33672 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_46_362
timestamp 1644511149
transform 1 0 34408 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_365
timestamp 1644511149
transform 1 0 34684 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_377
timestamp 1644511149
transform 1 0 35788 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_381
timestamp 1644511149
transform 1 0 36156 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_46_385
timestamp 1644511149
transform 1 0 36524 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_397
timestamp 1644511149
transform 1 0 37628 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_46_408
timestamp 1644511149
transform 1 0 38640 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_421
timestamp 1644511149
transform 1 0 39836 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_46_433
timestamp 1644511149
transform 1 0 40940 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_46_441
timestamp 1644511149
transform 1 0 41676 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_46_453
timestamp 1644511149
transform 1 0 42780 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_46_465
timestamp 1644511149
transform 1 0 43884 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_46_473
timestamp 1644511149
transform 1 0 44620 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_46_484
timestamp 1644511149
transform 1 0 45632 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_46_496
timestamp 1644511149
transform 1 0 46736 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_46_500
timestamp 1644511149
transform 1 0 47104 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_508
timestamp 1644511149
transform 1 0 47840 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_518
timestamp 1644511149
transform 1 0 48760 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_46_525
timestamp 1644511149
transform 1 0 49404 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_46_531
timestamp 1644511149
transform 1 0 49956 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_46_533
timestamp 1644511149
transform 1 0 50140 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_541
timestamp 1644511149
transform 1 0 50876 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_46_548
timestamp 1644511149
transform 1 0 51520 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_46_558
timestamp 1644511149
transform 1 0 52440 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_584
timestamp 1644511149
transform 1 0 54832 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_46_597
timestamp 1644511149
transform 1 0 56028 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_46_608
timestamp 1644511149
transform 1 0 57040 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_46_616
timestamp 1644511149
transform 1 0 57776 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_46_621
timestamp 1644511149
transform 1 0 58236 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_3
timestamp 1644511149
transform 1 0 1380 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_11
timestamp 1644511149
transform 1 0 2116 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_22
timestamp 1644511149
transform 1 0 3128 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_33
timestamp 1644511149
transform 1 0 4140 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_39
timestamp 1644511149
transform 1 0 4692 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_51
timestamp 1644511149
transform 1 0 5796 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_55
timestamp 1644511149
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_47_57
timestamp 1644511149
transform 1 0 6348 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_64
timestamp 1644511149
transform 1 0 6992 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_72
timestamp 1644511149
transform 1 0 7728 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_76
timestamp 1644511149
transform 1 0 8096 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_81
timestamp 1644511149
transform 1 0 8556 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_89
timestamp 1644511149
transform 1 0 9292 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_95
timestamp 1644511149
transform 1 0 9844 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_107
timestamp 1644511149
transform 1 0 10948 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_111
timestamp 1644511149
transform 1 0 11316 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_113
timestamp 1644511149
transform 1 0 11500 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_125
timestamp 1644511149
transform 1 0 12604 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_129
timestamp 1644511149
transform 1 0 12972 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_140
timestamp 1644511149
transform 1 0 13984 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_152
timestamp 1644511149
transform 1 0 15088 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_158
timestamp 1644511149
transform 1 0 15640 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_166
timestamp 1644511149
transform 1 0 16376 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_47_191
timestamp 1644511149
transform 1 0 18676 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_203
timestamp 1644511149
transform 1 0 19780 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_211
timestamp 1644511149
transform 1 0 20516 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_47_214
timestamp 1644511149
transform 1 0 20792 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_222
timestamp 1644511149
transform 1 0 21528 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_47_225
timestamp 1644511149
transform 1 0 21804 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_228
timestamp 1644511149
transform 1 0 22080 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_242
timestamp 1644511149
transform 1 0 23368 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_47_252
timestamp 1644511149
transform 1 0 24288 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_259
timestamp 1644511149
transform 1 0 24932 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_47_266
timestamp 1644511149
transform 1 0 25576 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_272
timestamp 1644511149
transform 1 0 26128 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_281
timestamp 1644511149
transform 1 0 26956 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_293
timestamp 1644511149
transform 1 0 28060 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_305
timestamp 1644511149
transform 1 0 29164 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_309
timestamp 1644511149
transform 1 0 29532 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_312
timestamp 1644511149
transform 1 0 29808 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_47_316
timestamp 1644511149
transform 1 0 30176 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_47_319
timestamp 1644511149
transform 1 0 30452 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_47_330
timestamp 1644511149
transform 1 0 31464 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_47_337
timestamp 1644511149
transform 1 0 32108 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_349
timestamp 1644511149
transform 1 0 33212 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_361
timestamp 1644511149
transform 1 0 34316 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_373
timestamp 1644511149
transform 1 0 35420 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_381
timestamp 1644511149
transform 1 0 36156 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_388
timestamp 1644511149
transform 1 0 36800 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_47_393
timestamp 1644511149
transform 1 0 37260 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_47_405
timestamp 1644511149
transform 1 0 38364 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_47_416
timestamp 1644511149
transform 1 0 39376 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_428
timestamp 1644511149
transform 1 0 40480 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_47_441
timestamp 1644511149
transform 1 0 41676 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_447
timestamp 1644511149
transform 1 0 42228 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_455
timestamp 1644511149
transform 1 0 42964 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_47_467
timestamp 1644511149
transform 1 0 44068 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_47_473
timestamp 1644511149
transform 1 0 44620 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_478
timestamp 1644511149
transform 1 0 45080 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_490
timestamp 1644511149
transform 1 0 46184 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_502
timestamp 1644511149
transform 1 0 47288 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_47_505
timestamp 1644511149
transform 1 0 47564 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_517
timestamp 1644511149
transform 1 0 48668 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_529
timestamp 1644511149
transform 1 0 49772 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_47_541
timestamp 1644511149
transform 1 0 50876 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_47_551
timestamp 1644511149
transform 1 0 51796 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_47_559
timestamp 1644511149
transform 1 0 52532 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_47_561
timestamp 1644511149
transform 1 0 52716 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_47_573
timestamp 1644511149
transform 1 0 53820 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_47_585
timestamp 1644511149
transform 1 0 54924 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_597
timestamp 1644511149
transform 1 0 56028 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_47_605
timestamp 1644511149
transform 1 0 56764 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_47_612
timestamp 1644511149
transform 1 0 57408 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_47_617
timestamp 1644511149
transform 1 0 57868 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_3
timestamp 1644511149
transform 1 0 1380 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_15
timestamp 1644511149
transform 1 0 2484 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_27
timestamp 1644511149
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_29
timestamp 1644511149
transform 1 0 3772 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_41
timestamp 1644511149
transform 1 0 4876 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_53
timestamp 1644511149
transform 1 0 5980 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_48_61
timestamp 1644511149
transform 1 0 6716 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_48_66
timestamp 1644511149
transform 1 0 7176 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_72
timestamp 1644511149
transform 1 0 7728 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_88
timestamp 1644511149
transform 1 0 9200 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_97
timestamp 1644511149
transform 1 0 10028 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_105
timestamp 1644511149
transform 1 0 10764 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_48_111
timestamp 1644511149
transform 1 0 11316 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_117
timestamp 1644511149
transform 1 0 11868 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_128
timestamp 1644511149
transform 1 0 12880 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_141
timestamp 1644511149
transform 1 0 14076 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_149
timestamp 1644511149
transform 1 0 14812 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_161
timestamp 1644511149
transform 1 0 15916 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_173
timestamp 1644511149
transform 1 0 17020 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_185
timestamp 1644511149
transform 1 0 18124 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_192
timestamp 1644511149
transform 1 0 18768 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_210
timestamp 1644511149
transform 1 0 20424 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_218
timestamp 1644511149
transform 1 0 21160 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_226
timestamp 1644511149
transform 1 0 21896 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_237
timestamp 1644511149
transform 1 0 22908 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_48_248
timestamp 1644511149
transform 1 0 23920 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_257
timestamp 1644511149
transform 1 0 24748 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_263
timestamp 1644511149
transform 1 0 25300 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_275
timestamp 1644511149
transform 1 0 26404 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_48_290
timestamp 1644511149
transform 1 0 27784 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_48_299
timestamp 1644511149
transform 1 0 28612 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_307
timestamp 1644511149
transform 1 0 29348 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_309
timestamp 1644511149
transform 1 0 29532 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_48_323
timestamp 1644511149
transform 1 0 30820 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_332
timestamp 1644511149
transform 1 0 31648 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_344
timestamp 1644511149
transform 1 0 32752 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_356
timestamp 1644511149
transform 1 0 33856 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_48_372
timestamp 1644511149
transform 1 0 35328 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_384
timestamp 1644511149
transform 1 0 36432 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_48_401
timestamp 1644511149
transform 1 0 37996 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_48_407
timestamp 1644511149
transform 1 0 38548 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_415
timestamp 1644511149
transform 1 0 39284 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_419
timestamp 1644511149
transform 1 0 39652 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_421
timestamp 1644511149
transform 1 0 39836 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_48_433
timestamp 1644511149
transform 1 0 40940 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_48_441
timestamp 1644511149
transform 1 0 41676 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_48_451
timestamp 1644511149
transform 1 0 42596 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_463
timestamp 1644511149
transform 1 0 43700 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_475
timestamp 1644511149
transform 1 0 44804 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_477
timestamp 1644511149
transform 1 0 44988 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_48_481
timestamp 1644511149
transform 1 0 45356 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_48_485
timestamp 1644511149
transform 1 0 45724 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_497
timestamp 1644511149
transform 1 0 46828 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_48_509
timestamp 1644511149
transform 1 0 47932 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_516
timestamp 1644511149
transform 1 0 48576 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_524
timestamp 1644511149
transform 1 0 49312 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_528
timestamp 1644511149
transform 1 0 49680 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_48_533
timestamp 1644511149
transform 1 0 50140 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_549
timestamp 1644511149
transform 1 0 51612 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_561
timestamp 1644511149
transform 1 0 52716 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_48_573
timestamp 1644511149
transform 1 0 53820 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_48_585
timestamp 1644511149
transform 1 0 54924 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_48_589
timestamp 1644511149
transform 1 0 55292 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_597
timestamp 1644511149
transform 1 0 56028 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_48_600
timestamp 1644511149
transform 1 0 56304 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_48_608
timestamp 1644511149
transform 1 0 57040 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_48_615
timestamp 1644511149
transform 1 0 57684 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_48_621
timestamp 1644511149
transform 1 0 58236 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_3
timestamp 1644511149
transform 1 0 1380 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_15
timestamp 1644511149
transform 1 0 2484 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_27
timestamp 1644511149
transform 1 0 3588 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_49_39
timestamp 1644511149
transform 1 0 4692 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_50
timestamp 1644511149
transform 1 0 5704 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_49_57
timestamp 1644511149
transform 1 0 6348 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_49_69
timestamp 1644511149
transform 1 0 7452 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_81
timestamp 1644511149
transform 1 0 8556 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_87
timestamp 1644511149
transform 1 0 9108 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_49_92
timestamp 1644511149
transform 1 0 9568 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_49_100
timestamp 1644511149
transform 1 0 10304 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_108
timestamp 1644511149
transform 1 0 11040 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_113
timestamp 1644511149
transform 1 0 11500 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_49_129
timestamp 1644511149
transform 1 0 12972 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_141
timestamp 1644511149
transform 1 0 14076 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_152
timestamp 1644511149
transform 1 0 15088 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_49_158
timestamp 1644511149
transform 1 0 15640 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_166
timestamp 1644511149
transform 1 0 16376 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_191
timestamp 1644511149
transform 1 0 18676 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_199
timestamp 1644511149
transform 1 0 19412 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_207
timestamp 1644511149
transform 1 0 20148 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_213
timestamp 1644511149
transform 1 0 20700 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_219
timestamp 1644511149
transform 1 0 21252 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_223
timestamp 1644511149
transform 1 0 21620 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_49_225
timestamp 1644511149
transform 1 0 21804 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_230
timestamp 1644511149
transform 1 0 22264 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_236
timestamp 1644511149
transform 1 0 22816 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_242
timestamp 1644511149
transform 1 0 23368 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_246
timestamp 1644511149
transform 1 0 23736 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_260
timestamp 1644511149
transform 1 0 25024 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_49_272
timestamp 1644511149
transform 1 0 26128 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_276
timestamp 1644511149
transform 1 0 26496 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_284
timestamp 1644511149
transform 1 0 27232 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_295
timestamp 1644511149
transform 1 0 28244 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_49_304
timestamp 1644511149
transform 1 0 29072 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_49_310
timestamp 1644511149
transform 1 0 29624 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_49_323
timestamp 1644511149
transform 1 0 30820 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_49_335
timestamp 1644511149
transform 1 0 31924 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_49_337
timestamp 1644511149
transform 1 0 32108 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_341
timestamp 1644511149
transform 1 0 32476 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_353
timestamp 1644511149
transform 1 0 33580 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_49_363
timestamp 1644511149
transform 1 0 34500 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_369
timestamp 1644511149
transform 1 0 35052 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_381
timestamp 1644511149
transform 1 0 36156 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_389
timestamp 1644511149
transform 1 0 36892 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_393
timestamp 1644511149
transform 1 0 37260 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_405
timestamp 1644511149
transform 1 0 38364 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_417
timestamp 1644511149
transform 1 0 39468 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_429
timestamp 1644511149
transform 1 0 40572 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_441
timestamp 1644511149
transform 1 0 41676 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_447
timestamp 1644511149
transform 1 0 42228 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_449
timestamp 1644511149
transform 1 0 42412 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_453
timestamp 1644511149
transform 1 0 42780 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_459
timestamp 1644511149
transform 1 0 43332 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_49_471
timestamp 1644511149
transform 1 0 44436 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_49_481
timestamp 1644511149
transform 1 0 45356 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_493
timestamp 1644511149
transform 1 0 46460 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_49_501
timestamp 1644511149
transform 1 0 47196 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_49_505
timestamp 1644511149
transform 1 0 47564 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_511
timestamp 1644511149
transform 1 0 48116 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_519
timestamp 1644511149
transform 1 0 48852 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_49_528
timestamp 1644511149
transform 1 0 49680 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_49_540
timestamp 1644511149
transform 1 0 50784 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_49_548
timestamp 1644511149
transform 1 0 51520 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_49_555
timestamp 1644511149
transform 1 0 52164 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_559
timestamp 1644511149
transform 1 0 52532 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_49_561
timestamp 1644511149
transform 1 0 52716 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_49_573
timestamp 1644511149
transform 1 0 53820 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_49_598
timestamp 1644511149
transform 1 0 56120 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_49_604
timestamp 1644511149
transform 1 0 56672 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_612
timestamp 1644511149
transform 1 0 57408 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_49_617
timestamp 1644511149
transform 1 0 57868 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_49_621
timestamp 1644511149
transform 1 0 58236 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_7
timestamp 1644511149
transform 1 0 1748 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_13
timestamp 1644511149
transform 1 0 2300 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_25
timestamp 1644511149
transform 1 0 3404 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_50_36
timestamp 1644511149
transform 1 0 4416 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_42
timestamp 1644511149
transform 1 0 4968 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_46
timestamp 1644511149
transform 1 0 5336 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_50_54
timestamp 1644511149
transform 1 0 6072 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_50_72
timestamp 1644511149
transform 1 0 7728 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_85
timestamp 1644511149
transform 1 0 8924 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_96
timestamp 1644511149
transform 1 0 9936 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_107
timestamp 1644511149
transform 1 0 10948 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_119
timestamp 1644511149
transform 1 0 12052 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_50_130
timestamp 1644511149
transform 1 0 13064 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_50_138
timestamp 1644511149
transform 1 0 13800 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_141
timestamp 1644511149
transform 1 0 14076 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_147
timestamp 1644511149
transform 1 0 14628 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_156
timestamp 1644511149
transform 1 0 15456 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_165
timestamp 1644511149
transform 1 0 16284 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_177
timestamp 1644511149
transform 1 0 17388 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_189
timestamp 1644511149
transform 1 0 18492 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_192
timestamp 1644511149
transform 1 0 18768 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_200
timestamp 1644511149
transform 1 0 19504 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_206
timestamp 1644511149
transform 1 0 20056 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_218
timestamp 1644511149
transform 1 0 21160 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_50_224
timestamp 1644511149
transform 1 0 21712 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_50_230
timestamp 1644511149
transform 1 0 22264 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_238
timestamp 1644511149
transform 1 0 23000 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_248
timestamp 1644511149
transform 1 0 23920 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_261
timestamp 1644511149
transform 1 0 25116 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_273
timestamp 1644511149
transform 1 0 26220 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_50_285
timestamp 1644511149
transform 1 0 27324 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_50_295
timestamp 1644511149
transform 1 0 28244 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_307
timestamp 1644511149
transform 1 0 29348 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_50_309
timestamp 1644511149
transform 1 0 29532 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_315
timestamp 1644511149
transform 1 0 30084 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_318
timestamp 1644511149
transform 1 0 30360 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_335
timestamp 1644511149
transform 1 0 31924 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_347
timestamp 1644511149
transform 1 0 33028 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_359
timestamp 1644511149
transform 1 0 34132 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_363
timestamp 1644511149
transform 1 0 34500 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_365
timestamp 1644511149
transform 1 0 34684 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_377
timestamp 1644511149
transform 1 0 35788 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_50_383
timestamp 1644511149
transform 1 0 36340 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_50_389
timestamp 1644511149
transform 1 0 36892 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_396
timestamp 1644511149
transform 1 0 37536 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_408
timestamp 1644511149
transform 1 0 38640 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_421
timestamp 1644511149
transform 1 0 39836 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_50_433
timestamp 1644511149
transform 1 0 40940 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_445
timestamp 1644511149
transform 1 0 42044 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_50_456
timestamp 1644511149
transform 1 0 43056 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_50_468
timestamp 1644511149
transform 1 0 44160 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_50_482
timestamp 1644511149
transform 1 0 45448 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_50_494
timestamp 1644511149
transform 1 0 46552 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_50_509
timestamp 1644511149
transform 1 0 47932 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_50_519
timestamp 1644511149
transform 1 0 48852 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_50_531
timestamp 1644511149
transform 1 0 49956 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_50_533
timestamp 1644511149
transform 1 0 50140 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_50_545
timestamp 1644511149
transform 1 0 51244 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_50_570
timestamp 1644511149
transform 1 0 53544 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_50_582
timestamp 1644511149
transform 1 0 54648 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_50_606
timestamp 1644511149
transform 1 0 56856 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_50_620
timestamp 1644511149
transform 1 0 58144 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_50_624
timestamp 1644511149
transform 1 0 58512 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_3
timestamp 1644511149
transform 1 0 1380 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_15
timestamp 1644511149
transform 1 0 2484 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_27
timestamp 1644511149
transform 1 0 3588 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_39
timestamp 1644511149
transform 1 0 4692 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_51
timestamp 1644511149
transform 1 0 5796 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_55
timestamp 1644511149
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_57
timestamp 1644511149
transform 1 0 6348 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_65
timestamp 1644511149
transform 1 0 7084 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_72
timestamp 1644511149
transform 1 0 7728 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_84
timestamp 1644511149
transform 1 0 8832 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_51_98
timestamp 1644511149
transform 1 0 10120 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_104
timestamp 1644511149
transform 1 0 10672 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_51_113
timestamp 1644511149
transform 1 0 11500 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_125
timestamp 1644511149
transform 1 0 12604 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_51_132
timestamp 1644511149
transform 1 0 13248 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_144
timestamp 1644511149
transform 1 0 14352 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_51_152
timestamp 1644511149
transform 1 0 15088 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_164
timestamp 1644511149
transform 1 0 16192 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_175
timestamp 1644511149
transform 1 0 17204 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_193
timestamp 1644511149
transform 1 0 18860 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_201
timestamp 1644511149
transform 1 0 19596 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_209
timestamp 1644511149
transform 1 0 20332 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_217
timestamp 1644511149
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_223
timestamp 1644511149
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_225
timestamp 1644511149
transform 1 0 21804 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_231
timestamp 1644511149
transform 1 0 22356 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_234
timestamp 1644511149
transform 1 0 22632 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_241
timestamp 1644511149
transform 1 0 23276 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_249
timestamp 1644511149
transform 1 0 24012 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_255
timestamp 1644511149
transform 1 0 24564 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_261
timestamp 1644511149
transform 1 0 25116 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_273
timestamp 1644511149
transform 1 0 26220 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_279
timestamp 1644511149
transform 1 0 26772 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_281
timestamp 1644511149
transform 1 0 26956 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_285
timestamp 1644511149
transform 1 0 27324 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_288
timestamp 1644511149
transform 1 0 27600 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_300
timestamp 1644511149
transform 1 0 28704 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_312
timestamp 1644511149
transform 1 0 29808 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_51_320
timestamp 1644511149
transform 1 0 30544 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_51_332
timestamp 1644511149
transform 1 0 31648 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_51_337
timestamp 1644511149
transform 1 0 32108 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_51_341
timestamp 1644511149
transform 1 0 32476 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_355
timestamp 1644511149
transform 1 0 33764 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_367
timestamp 1644511149
transform 1 0 34868 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_375
timestamp 1644511149
transform 1 0 35604 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_385
timestamp 1644511149
transform 1 0 36524 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_391
timestamp 1644511149
transform 1 0 37076 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_51_403
timestamp 1644511149
transform 1 0 38180 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_51_415
timestamp 1644511149
transform 1 0 39284 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_51_425
timestamp 1644511149
transform 1 0 40204 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_435
timestamp 1644511149
transform 1 0 41124 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_51_447
timestamp 1644511149
transform 1 0 42228 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_453
timestamp 1644511149
transform 1 0 42780 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_51_462
timestamp 1644511149
transform 1 0 43608 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_468
timestamp 1644511149
transform 1 0 44160 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_472
timestamp 1644511149
transform 1 0 44528 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_483
timestamp 1644511149
transform 1 0 45540 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_51_495
timestamp 1644511149
transform 1 0 46644 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_503
timestamp 1644511149
transform 1 0 47380 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_505
timestamp 1644511149
transform 1 0 47564 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_51_517
timestamp 1644511149
transform 1 0 48668 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_51_529
timestamp 1644511149
transform 1 0 49772 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_51_541
timestamp 1644511149
transform 1 0 50876 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_51_556
timestamp 1644511149
transform 1 0 52256 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_51_568
timestamp 1644511149
transform 1 0 53360 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_51_580
timestamp 1644511149
transform 1 0 54464 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_51_586
timestamp 1644511149
transform 1 0 55016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_51_592
timestamp 1644511149
transform 1 0 55568 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_51_599
timestamp 1644511149
transform 1 0 56212 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_51_607
timestamp 1644511149
transform 1 0 56948 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_51_610
timestamp 1644511149
transform 1 0 57224 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_51_617
timestamp 1644511149
transform 1 0 57868 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_52_3
timestamp 1644511149
transform 1 0 1380 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_15
timestamp 1644511149
transform 1 0 2484 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_27
timestamp 1644511149
transform 1 0 3588 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_29
timestamp 1644511149
transform 1 0 3772 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_41
timestamp 1644511149
transform 1 0 4876 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_53
timestamp 1644511149
transform 1 0 5980 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_65
timestamp 1644511149
transform 1 0 7084 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_70
timestamp 1644511149
transform 1 0 7544 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_52_82
timestamp 1644511149
transform 1 0 8648 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_52_85
timestamp 1644511149
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_104
timestamp 1644511149
transform 1 0 10672 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_116
timestamp 1644511149
transform 1 0 11776 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_128
timestamp 1644511149
transform 1 0 12880 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_52_134
timestamp 1644511149
transform 1 0 13432 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_52_163
timestamp 1644511149
transform 1 0 16100 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_175
timestamp 1644511149
transform 1 0 17204 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_180
timestamp 1644511149
transform 1 0 17664 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_191
timestamp 1644511149
transform 1 0 18676 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_52_195
timestamp 1644511149
transform 1 0 19044 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_199
timestamp 1644511149
transform 1 0 19412 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_205
timestamp 1644511149
transform 1 0 19964 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_217
timestamp 1644511149
transform 1 0 21068 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_225
timestamp 1644511149
transform 1 0 21804 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_52_230
timestamp 1644511149
transform 1 0 22264 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_240
timestamp 1644511149
transform 1 0 23184 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_255
timestamp 1644511149
transform 1 0 24564 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_267
timestamp 1644511149
transform 1 0 25668 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_286
timestamp 1644511149
transform 1 0 27416 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_295
timestamp 1644511149
transform 1 0 28244 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_52_301
timestamp 1644511149
transform 1 0 28796 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_307
timestamp 1644511149
transform 1 0 29348 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_52_309
timestamp 1644511149
transform 1 0 29532 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_317
timestamp 1644511149
transform 1 0 30268 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_52_325
timestamp 1644511149
transform 1 0 31004 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_331
timestamp 1644511149
transform 1 0 31556 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_343
timestamp 1644511149
transform 1 0 32660 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_52_355
timestamp 1644511149
transform 1 0 33764 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_52_363
timestamp 1644511149
transform 1 0 34500 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_365
timestamp 1644511149
transform 1 0 34684 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_377
timestamp 1644511149
transform 1 0 35788 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_52_389
timestamp 1644511149
transform 1 0 36892 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_52_395
timestamp 1644511149
transform 1 0 37444 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_407
timestamp 1644511149
transform 1 0 38548 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_52_419
timestamp 1644511149
transform 1 0 39652 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_421
timestamp 1644511149
transform 1 0 39836 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_433
timestamp 1644511149
transform 1 0 40940 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_445
timestamp 1644511149
transform 1 0 42044 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_457
timestamp 1644511149
transform 1 0 43148 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_52_469
timestamp 1644511149
transform 1 0 44252 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_52_475
timestamp 1644511149
transform 1 0 44804 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_52_485
timestamp 1644511149
transform 1 0 45724 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_497
timestamp 1644511149
transform 1 0 46828 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_509
timestamp 1644511149
transform 1 0 47932 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_52_521
timestamp 1644511149
transform 1 0 49036 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_52_529
timestamp 1644511149
transform 1 0 49772 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_52_533
timestamp 1644511149
transform 1 0 50140 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_52_546
timestamp 1644511149
transform 1 0 51336 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_572
timestamp 1644511149
transform 1 0 53728 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_52_584
timestamp 1644511149
transform 1 0 54832 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_52_595
timestamp 1644511149
transform 1 0 55844 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_52_601
timestamp 1644511149
transform 1 0 56396 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_52_613
timestamp 1644511149
transform 1 0 57500 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_3
timestamp 1644511149
transform 1 0 1380 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_53_7
timestamp 1644511149
transform 1 0 1748 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_19
timestamp 1644511149
transform 1 0 2852 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_31
timestamp 1644511149
transform 1 0 3956 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_43
timestamp 1644511149
transform 1 0 5060 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_55
timestamp 1644511149
transform 1 0 6164 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_53_57
timestamp 1644511149
transform 1 0 6348 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_53_77
timestamp 1644511149
transform 1 0 8188 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_89
timestamp 1644511149
transform 1 0 9292 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_93
timestamp 1644511149
transform 1 0 9660 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_99
timestamp 1644511149
transform 1 0 10212 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_111
timestamp 1644511149
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_113
timestamp 1644511149
transform 1 0 11500 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_125
timestamp 1644511149
transform 1 0 12604 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_138
timestamp 1644511149
transform 1 0 13800 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_150
timestamp 1644511149
transform 1 0 14904 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_162
timestamp 1644511149
transform 1 0 16008 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_53_169
timestamp 1644511149
transform 1 0 16652 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_53_181
timestamp 1644511149
transform 1 0 17756 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_53_192
timestamp 1644511149
transform 1 0 18768 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_204
timestamp 1644511149
transform 1 0 19872 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_53_216
timestamp 1644511149
transform 1 0 20976 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_220
timestamp 1644511149
transform 1 0 21344 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_232
timestamp 1644511149
transform 1 0 22448 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_238
timestamp 1644511149
transform 1 0 23000 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_250
timestamp 1644511149
transform 1 0 24104 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_262
timestamp 1644511149
transform 1 0 25208 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_274
timestamp 1644511149
transform 1 0 26312 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_53_289
timestamp 1644511149
transform 1 0 27692 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_300
timestamp 1644511149
transform 1 0 28704 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_53_306
timestamp 1644511149
transform 1 0 29256 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_316
timestamp 1644511149
transform 1 0 30176 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_328
timestamp 1644511149
transform 1 0 31280 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_53_343
timestamp 1644511149
transform 1 0 32660 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_355
timestamp 1644511149
transform 1 0 33764 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_367
timestamp 1644511149
transform 1 0 34868 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_379
timestamp 1644511149
transform 1 0 35972 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_53_391
timestamp 1644511149
transform 1 0 37076 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_400
timestamp 1644511149
transform 1 0 37904 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_412
timestamp 1644511149
transform 1 0 39008 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_424
timestamp 1644511149
transform 1 0 40112 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_53_428
timestamp 1644511149
transform 1 0 40480 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_53_436
timestamp 1644511149
transform 1 0 41216 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_449
timestamp 1644511149
transform 1 0 42412 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_461
timestamp 1644511149
transform 1 0 43516 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_53_469
timestamp 1644511149
transform 1 0 44252 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_53_477
timestamp 1644511149
transform 1 0 44988 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_488
timestamp 1644511149
transform 1 0 46000 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_53_500
timestamp 1644511149
transform 1 0 47104 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_53_505
timestamp 1644511149
transform 1 0 47564 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_53_520
timestamp 1644511149
transform 1 0 48944 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_530
timestamp 1644511149
transform 1 0 49864 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_53_542
timestamp 1644511149
transform 1 0 50968 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_53_548
timestamp 1644511149
transform 1 0 51520 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_53_556
timestamp 1644511149
transform 1 0 52256 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_53_561
timestamp 1644511149
transform 1 0 52716 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_573
timestamp 1644511149
transform 1 0 53820 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_592
timestamp 1644511149
transform 1 0 55568 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_53_604
timestamp 1644511149
transform 1 0 56672 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_53_617
timestamp 1644511149
transform 1 0 57868 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_54_3
timestamp 1644511149
transform 1 0 1380 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_11
timestamp 1644511149
transform 1 0 2116 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_18
timestamp 1644511149
transform 1 0 2760 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_24
timestamp 1644511149
transform 1 0 3312 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_29
timestamp 1644511149
transform 1 0 3772 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_41
timestamp 1644511149
transform 1 0 4876 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_53
timestamp 1644511149
transform 1 0 5980 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_57
timestamp 1644511149
transform 1 0 6348 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_80
timestamp 1644511149
transform 1 0 8464 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_91
timestamp 1644511149
transform 1 0 9476 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_99
timestamp 1644511149
transform 1 0 10212 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_108
timestamp 1644511149
transform 1 0 11040 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_120
timestamp 1644511149
transform 1 0 12144 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_136
timestamp 1644511149
transform 1 0 13616 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_141
timestamp 1644511149
transform 1 0 14076 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_54_159
timestamp 1644511149
transform 1 0 15732 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_168
timestamp 1644511149
transform 1 0 16560 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_54_172
timestamp 1644511149
transform 1 0 16928 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_175
timestamp 1644511149
transform 1 0 17204 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_54_189
timestamp 1644511149
transform 1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_195
timestamp 1644511149
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_54_197
timestamp 1644511149
transform 1 0 19228 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_205
timestamp 1644511149
transform 1 0 19964 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_209
timestamp 1644511149
transform 1 0 20332 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_226
timestamp 1644511149
transform 1 0 21896 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_237
timestamp 1644511149
transform 1 0 22908 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_243
timestamp 1644511149
transform 1 0 23460 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_251
timestamp 1644511149
transform 1 0 24196 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_260
timestamp 1644511149
transform 1 0 25024 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_272
timestamp 1644511149
transform 1 0 26128 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_54_278
timestamp 1644511149
transform 1 0 26680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_287
timestamp 1644511149
transform 1 0 27508 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_299
timestamp 1644511149
transform 1 0 28612 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_304
timestamp 1644511149
transform 1 0 29072 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_322
timestamp 1644511149
transform 1 0 30728 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_334
timestamp 1644511149
transform 1 0 31832 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_54_343
timestamp 1644511149
transform 1 0 32660 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_54_355
timestamp 1644511149
transform 1 0 33764 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_54_360
timestamp 1644511149
transform 1 0 34224 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_378
timestamp 1644511149
transform 1 0 35880 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_390
timestamp 1644511149
transform 1 0 36984 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_54_398
timestamp 1644511149
transform 1 0 37720 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_54_404
timestamp 1644511149
transform 1 0 38272 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_416
timestamp 1644511149
transform 1 0 39376 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_54_421
timestamp 1644511149
transform 1 0 39836 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_433
timestamp 1644511149
transform 1 0 40940 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_54_444
timestamp 1644511149
transform 1 0 41952 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_54_456
timestamp 1644511149
transform 1 0 43056 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_468
timestamp 1644511149
transform 1 0 44160 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_477
timestamp 1644511149
transform 1 0 44988 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_54_487
timestamp 1644511149
transform 1 0 45908 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_54_499
timestamp 1644511149
transform 1 0 47012 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_507
timestamp 1644511149
transform 1 0 47748 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_511
timestamp 1644511149
transform 1 0 48116 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_54_522
timestamp 1644511149
transform 1 0 49128 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_54_530
timestamp 1644511149
transform 1 0 49864 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_54_533
timestamp 1644511149
transform 1 0 50140 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_54_545
timestamp 1644511149
transform 1 0 51244 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_54_573
timestamp 1644511149
transform 1 0 53820 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_54_585
timestamp 1644511149
transform 1 0 54924 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_54_602
timestamp 1644511149
transform 1 0 56488 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_54_610
timestamp 1644511149
transform 1 0 57224 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_54_613
timestamp 1644511149
transform 1 0 57500 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_54_621
timestamp 1644511149
transform 1 0 58236 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_3
timestamp 1644511149
transform 1 0 1380 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_15
timestamp 1644511149
transform 1 0 2484 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_27
timestamp 1644511149
transform 1 0 3588 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_39
timestamp 1644511149
transform 1 0 4692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_51
timestamp 1644511149
transform 1 0 5796 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_55
timestamp 1644511149
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_57
timestamp 1644511149
transform 1 0 6348 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_55_87
timestamp 1644511149
transform 1 0 9108 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_55_93
timestamp 1644511149
transform 1 0 9660 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_55_105
timestamp 1644511149
transform 1 0 10764 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_111
timestamp 1644511149
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_113
timestamp 1644511149
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_125
timestamp 1644511149
transform 1 0 12604 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_55_149
timestamp 1644511149
transform 1 0 14812 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_55_156
timestamp 1644511149
transform 1 0 15456 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_175
timestamp 1644511149
transform 1 0 17204 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_181
timestamp 1644511149
transform 1 0 17756 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_185
timestamp 1644511149
transform 1 0 18124 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_192
timestamp 1644511149
transform 1 0 18768 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_204
timestamp 1644511149
transform 1 0 19872 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_216
timestamp 1644511149
transform 1 0 20976 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_55_225
timestamp 1644511149
transform 1 0 21804 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_55_233
timestamp 1644511149
transform 1 0 22540 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_245
timestamp 1644511149
transform 1 0 23644 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_55_256
timestamp 1644511149
transform 1 0 24656 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_268
timestamp 1644511149
transform 1 0 25760 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_283
timestamp 1644511149
transform 1 0 27140 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_287
timestamp 1644511149
transform 1 0 27508 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_290
timestamp 1644511149
transform 1 0 27784 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_302
timestamp 1644511149
transform 1 0 28888 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_55_314
timestamp 1644511149
transform 1 0 29992 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_318
timestamp 1644511149
transform 1 0 30360 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_322
timestamp 1644511149
transform 1 0 30728 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_334
timestamp 1644511149
transform 1 0 31832 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_55_337
timestamp 1644511149
transform 1 0 32108 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_349
timestamp 1644511149
transform 1 0 33212 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_55_358
timestamp 1644511149
transform 1 0 34040 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_362
timestamp 1644511149
transform 1 0 34408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_369
timestamp 1644511149
transform 1 0 35052 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_381
timestamp 1644511149
transform 1 0 36156 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_389
timestamp 1644511149
transform 1 0 36892 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_55_399
timestamp 1644511149
transform 1 0 37812 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_55_406
timestamp 1644511149
transform 1 0 38456 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_55_410
timestamp 1644511149
transform 1 0 38824 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_424
timestamp 1644511149
transform 1 0 40112 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_55_432
timestamp 1644511149
transform 1 0 40848 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_55_442
timestamp 1644511149
transform 1 0 41768 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_55_449
timestamp 1644511149
transform 1 0 42412 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_55_464
timestamp 1644511149
transform 1 0 43792 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_476
timestamp 1644511149
transform 1 0 44896 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_55_485
timestamp 1644511149
transform 1 0 45724 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_55_497
timestamp 1644511149
transform 1 0 46828 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_55_503
timestamp 1644511149
transform 1 0 47380 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_55_505
timestamp 1644511149
transform 1 0 47564 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_513
timestamp 1644511149
transform 1 0 48300 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_527
timestamp 1644511149
transform 1 0 49588 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_539
timestamp 1644511149
transform 1 0 50692 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_55_551
timestamp 1644511149
transform 1 0 51796 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_55_559
timestamp 1644511149
transform 1 0 52532 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_55_566
timestamp 1644511149
transform 1 0 53176 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_578
timestamp 1644511149
transform 1 0 54280 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_590
timestamp 1644511149
transform 1 0 55384 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_55_602
timestamp 1644511149
transform 1 0 56488 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_55_614
timestamp 1644511149
transform 1 0 57592 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_55_617
timestamp 1644511149
transform 1 0 57868 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_56_3
timestamp 1644511149
transform 1 0 1380 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_56_7
timestamp 1644511149
transform 1 0 1748 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_19
timestamp 1644511149
transform 1 0 2852 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_27
timestamp 1644511149
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_29
timestamp 1644511149
transform 1 0 3772 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_41
timestamp 1644511149
transform 1 0 4876 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_53
timestamp 1644511149
transform 1 0 5980 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_56_72
timestamp 1644511149
transform 1 0 7728 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_80
timestamp 1644511149
transform 1 0 8464 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_87
timestamp 1644511149
transform 1 0 9108 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_99
timestamp 1644511149
transform 1 0 10212 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_111
timestamp 1644511149
transform 1 0 11316 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_56_126
timestamp 1644511149
transform 1 0 12696 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_138
timestamp 1644511149
transform 1 0 13800 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_56_141
timestamp 1644511149
transform 1 0 14076 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_153
timestamp 1644511149
transform 1 0 15180 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_161
timestamp 1644511149
transform 1 0 15916 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_171
timestamp 1644511149
transform 1 0 16836 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_56_177
timestamp 1644511149
transform 1 0 17388 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_185
timestamp 1644511149
transform 1 0 18124 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_56_190
timestamp 1644511149
transform 1 0 18584 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_204
timestamp 1644511149
transform 1 0 19872 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_210
timestamp 1644511149
transform 1 0 20424 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_56_222
timestamp 1644511149
transform 1 0 21528 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_56_237
timestamp 1644511149
transform 1 0 22908 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_56_249
timestamp 1644511149
transform 1 0 24012 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_253
timestamp 1644511149
transform 1 0 24380 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_265
timestamp 1644511149
transform 1 0 25484 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_56_280
timestamp 1644511149
transform 1 0 26864 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_288
timestamp 1644511149
transform 1 0 27600 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_56_296
timestamp 1644511149
transform 1 0 28336 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_309
timestamp 1644511149
transform 1 0 29532 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_315
timestamp 1644511149
transform 1 0 30084 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_329
timestamp 1644511149
transform 1 0 31372 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_341
timestamp 1644511149
transform 1 0 32476 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_353
timestamp 1644511149
transform 1 0 33580 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_361
timestamp 1644511149
transform 1 0 34316 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_56_378
timestamp 1644511149
transform 1 0 35880 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_56_390
timestamp 1644511149
transform 1 0 36984 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_56_398
timestamp 1644511149
transform 1 0 37720 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_401
timestamp 1644511149
transform 1 0 37996 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_405
timestamp 1644511149
transform 1 0 38364 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_412
timestamp 1644511149
transform 1 0 39008 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_56_421
timestamp 1644511149
transform 1 0 39836 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_433
timestamp 1644511149
transform 1 0 40940 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_445
timestamp 1644511149
transform 1 0 42044 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_457
timestamp 1644511149
transform 1 0 43148 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_469
timestamp 1644511149
transform 1 0 44252 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_475
timestamp 1644511149
transform 1 0 44804 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_56_480
timestamp 1644511149
transform 1 0 45264 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_484
timestamp 1644511149
transform 1 0 45632 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_56_507
timestamp 1644511149
transform 1 0 47748 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_56_515
timestamp 1644511149
transform 1 0 48484 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_56_521
timestamp 1644511149
transform 1 0 49036 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_56_527
timestamp 1644511149
transform 1 0 49588 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_56_531
timestamp 1644511149
transform 1 0 49956 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_533
timestamp 1644511149
transform 1 0 50140 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_545
timestamp 1644511149
transform 1 0 51244 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_557
timestamp 1644511149
transform 1 0 52348 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_569
timestamp 1644511149
transform 1 0 53452 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_581
timestamp 1644511149
transform 1 0 54556 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_56_587
timestamp 1644511149
transform 1 0 55108 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_56_589
timestamp 1644511149
transform 1 0 55292 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_56_601
timestamp 1644511149
transform 1 0 56396 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_56_613
timestamp 1644511149
transform 1 0 57500 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_56_621
timestamp 1644511149
transform 1 0 58236 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_3
timestamp 1644511149
transform 1 0 1380 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_11
timestamp 1644511149
transform 1 0 2116 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_23
timestamp 1644511149
transform 1 0 3220 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_35
timestamp 1644511149
transform 1 0 4324 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_47
timestamp 1644511149
transform 1 0 5428 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_55
timestamp 1644511149
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_57_57
timestamp 1644511149
transform 1 0 6348 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_64
timestamp 1644511149
transform 1 0 6992 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_75
timestamp 1644511149
transform 1 0 8004 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_82
timestamp 1644511149
transform 1 0 8648 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_88
timestamp 1644511149
transform 1 0 9200 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_94
timestamp 1644511149
transform 1 0 9752 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_106
timestamp 1644511149
transform 1 0 10856 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_57_113
timestamp 1644511149
transform 1 0 11500 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_57_121
timestamp 1644511149
transform 1 0 12236 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_133
timestamp 1644511149
transform 1 0 13340 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_145
timestamp 1644511149
transform 1 0 14444 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_157
timestamp 1644511149
transform 1 0 15548 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_57_165
timestamp 1644511149
transform 1 0 16284 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_169
timestamp 1644511149
transform 1 0 16652 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_57_179
timestamp 1644511149
transform 1 0 17572 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_185
timestamp 1644511149
transform 1 0 18124 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_197
timestamp 1644511149
transform 1 0 19228 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_209
timestamp 1644511149
transform 1 0 20332 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_221
timestamp 1644511149
transform 1 0 21436 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_57_225
timestamp 1644511149
transform 1 0 21804 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_233
timestamp 1644511149
transform 1 0 22540 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_57_242
timestamp 1644511149
transform 1 0 23368 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_254
timestamp 1644511149
transform 1 0 24472 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_57_263
timestamp 1644511149
transform 1 0 25300 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_57_275
timestamp 1644511149
transform 1 0 26404 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_57_279
timestamp 1644511149
transform 1 0 26772 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_57_283
timestamp 1644511149
transform 1 0 27140 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_57_291
timestamp 1644511149
transform 1 0 27876 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_297
timestamp 1644511149
transform 1 0 28428 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_305
timestamp 1644511149
transform 1 0 29164 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_317
timestamp 1644511149
transform 1 0 30268 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_323
timestamp 1644511149
transform 1 0 30820 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_57_330
timestamp 1644511149
transform 1 0 31464 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_57_337
timestamp 1644511149
transform 1 0 32108 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_349
timestamp 1644511149
transform 1 0 33212 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_361
timestamp 1644511149
transform 1 0 34316 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_57_373
timestamp 1644511149
transform 1 0 35420 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_57_382
timestamp 1644511149
transform 1 0 36248 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_57_390
timestamp 1644511149
transform 1 0 36984 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_57_393
timestamp 1644511149
transform 1 0 37260 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_405
timestamp 1644511149
transform 1 0 38364 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_417
timestamp 1644511149
transform 1 0 39468 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_429
timestamp 1644511149
transform 1 0 40572 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_441
timestamp 1644511149
transform 1 0 41676 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_447
timestamp 1644511149
transform 1 0 42228 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_452
timestamp 1644511149
transform 1 0 42688 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_57_464
timestamp 1644511149
transform 1 0 43792 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_57_472
timestamp 1644511149
transform 1 0 44528 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_57_485
timestamp 1644511149
transform 1 0 45724 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_497
timestamp 1644511149
transform 1 0 46828 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_57_503
timestamp 1644511149
transform 1 0 47380 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_57_505
timestamp 1644511149
transform 1 0 47564 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_57_510
timestamp 1644511149
transform 1 0 48024 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_536
timestamp 1644511149
transform 1 0 50416 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_57_548
timestamp 1644511149
transform 1 0 51520 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_57_556
timestamp 1644511149
transform 1 0 52256 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_57_566
timestamp 1644511149
transform 1 0 53176 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_578
timestamp 1644511149
transform 1 0 54280 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_590
timestamp 1644511149
transform 1 0 55384 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_57_602
timestamp 1644511149
transform 1 0 56488 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_57_614
timestamp 1644511149
transform 1 0 57592 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_57_621
timestamp 1644511149
transform 1 0 58236 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_3
timestamp 1644511149
transform 1 0 1380 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_15
timestamp 1644511149
transform 1 0 2484 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_27
timestamp 1644511149
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_29
timestamp 1644511149
transform 1 0 3772 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_41
timestamp 1644511149
transform 1 0 4876 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_53
timestamp 1644511149
transform 1 0 5980 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_65
timestamp 1644511149
transform 1 0 7084 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_69
timestamp 1644511149
transform 1 0 7452 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_80
timestamp 1644511149
transform 1 0 8464 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_85
timestamp 1644511149
transform 1 0 8924 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_93
timestamp 1644511149
transform 1 0 9660 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_105
timestamp 1644511149
transform 1 0 10764 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_109
timestamp 1644511149
transform 1 0 11132 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_129
timestamp 1644511149
transform 1 0 12972 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_58_137
timestamp 1644511149
transform 1 0 13708 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_58_141
timestamp 1644511149
transform 1 0 14076 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_149
timestamp 1644511149
transform 1 0 14812 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_154
timestamp 1644511149
transform 1 0 15272 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_163
timestamp 1644511149
transform 1 0 16100 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_175
timestamp 1644511149
transform 1 0 17204 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_58_187
timestamp 1644511149
transform 1 0 18308 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_192
timestamp 1644511149
transform 1 0 18768 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_203
timestamp 1644511149
transform 1 0 19780 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_215
timestamp 1644511149
transform 1 0 20884 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_58_227
timestamp 1644511149
transform 1 0 21988 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_58_246
timestamp 1644511149
transform 1 0 23736 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_58_253
timestamp 1644511149
transform 1 0 24380 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_58_262
timestamp 1644511149
transform 1 0 25208 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_274
timestamp 1644511149
transform 1 0 26312 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_58_286
timestamp 1644511149
transform 1 0 27416 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_294
timestamp 1644511149
transform 1 0 28152 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_303
timestamp 1644511149
transform 1 0 28980 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_307
timestamp 1644511149
transform 1 0 29348 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_309
timestamp 1644511149
transform 1 0 29532 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_321
timestamp 1644511149
transform 1 0 30636 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_325
timestamp 1644511149
transform 1 0 31004 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_58_339
timestamp 1644511149
transform 1 0 32292 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_349
timestamp 1644511149
transform 1 0 33212 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_58_361
timestamp 1644511149
transform 1 0 34316 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_58_365
timestamp 1644511149
transform 1 0 34684 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_58_382
timestamp 1644511149
transform 1 0 36248 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_390
timestamp 1644511149
transform 1 0 36984 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_395
timestamp 1644511149
transform 1 0 37444 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_58_399
timestamp 1644511149
transform 1 0 37812 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_406
timestamp 1644511149
transform 1 0 38456 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_58_418
timestamp 1644511149
transform 1 0 39560 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_58_421
timestamp 1644511149
transform 1 0 39836 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_425
timestamp 1644511149
transform 1 0 40204 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_58_434
timestamp 1644511149
transform 1 0 41032 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_440
timestamp 1644511149
transform 1 0 41584 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_58_448
timestamp 1644511149
transform 1 0 42320 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_58_460
timestamp 1644511149
transform 1 0 43424 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_469
timestamp 1644511149
transform 1 0 44252 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_58_475
timestamp 1644511149
transform 1 0 44804 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_58_483
timestamp 1644511149
transform 1 0 45540 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_495
timestamp 1644511149
transform 1 0 46644 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_58_507
timestamp 1644511149
transform 1 0 47748 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_58_515
timestamp 1644511149
transform 1 0 48484 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_58_519
timestamp 1644511149
transform 1 0 48852 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_528
timestamp 1644511149
transform 1 0 49680 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_58_533
timestamp 1644511149
transform 1 0 50140 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_58_541
timestamp 1644511149
transform 1 0 50876 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_58_551
timestamp 1644511149
transform 1 0 51796 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_572
timestamp 1644511149
transform 1 0 53728 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_58_584
timestamp 1644511149
transform 1 0 54832 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_58_589
timestamp 1644511149
transform 1 0 55292 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_601
timestamp 1644511149
transform 1 0 56396 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_58_613
timestamp 1644511149
transform 1 0 57500 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_3
timestamp 1644511149
transform 1 0 1380 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_15
timestamp 1644511149
transform 1 0 2484 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_27
timestamp 1644511149
transform 1 0 3588 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_39
timestamp 1644511149
transform 1 0 4692 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_51
timestamp 1644511149
transform 1 0 5796 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_55
timestamp 1644511149
transform 1 0 6164 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_57
timestamp 1644511149
transform 1 0 6348 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_59_67
timestamp 1644511149
transform 1 0 7268 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_76
timestamp 1644511149
transform 1 0 8096 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_82
timestamp 1644511149
transform 1 0 8648 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_88
timestamp 1644511149
transform 1 0 9200 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_59_100
timestamp 1644511149
transform 1 0 10304 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_59_108
timestamp 1644511149
transform 1 0 11040 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_117
timestamp 1644511149
transform 1 0 11868 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_59_143
timestamp 1644511149
transform 1 0 14260 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_59_164
timestamp 1644511149
transform 1 0 16192 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_172
timestamp 1644511149
transform 1 0 16928 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_184
timestamp 1644511149
transform 1 0 18032 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_59_189
timestamp 1644511149
transform 1 0 18492 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_201
timestamp 1644511149
transform 1 0 19596 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_59_205
timestamp 1644511149
transform 1 0 19964 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_209
timestamp 1644511149
transform 1 0 20332 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_59_218
timestamp 1644511149
transform 1 0 21160 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_59_225
timestamp 1644511149
transform 1 0 21804 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_237
timestamp 1644511149
transform 1 0 22908 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_249
timestamp 1644511149
transform 1 0 24012 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_257
timestamp 1644511149
transform 1 0 24748 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_59_265
timestamp 1644511149
transform 1 0 25484 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_59_277
timestamp 1644511149
transform 1 0 26588 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_59_281
timestamp 1644511149
transform 1 0 26956 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_285
timestamp 1644511149
transform 1 0 27324 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_293
timestamp 1644511149
transform 1 0 28060 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_299
timestamp 1644511149
transform 1 0 28612 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_311
timestamp 1644511149
transform 1 0 29716 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_323
timestamp 1644511149
transform 1 0 30820 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_335
timestamp 1644511149
transform 1 0 31924 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_59_359
timestamp 1644511149
transform 1 0 34132 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_59_367
timestamp 1644511149
transform 1 0 34868 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_373
timestamp 1644511149
transform 1 0 35420 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_380
timestamp 1644511149
transform 1 0 36064 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_59_393
timestamp 1644511149
transform 1 0 37260 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_404
timestamp 1644511149
transform 1 0 38272 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_415
timestamp 1644511149
transform 1 0 39284 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_426
timestamp 1644511149
transform 1 0 40296 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_438
timestamp 1644511149
transform 1 0 41400 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_446
timestamp 1644511149
transform 1 0 42136 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_59_449
timestamp 1644511149
transform 1 0 42412 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_59_458
timestamp 1644511149
transform 1 0 43240 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_470
timestamp 1644511149
transform 1 0 44344 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_482
timestamp 1644511149
transform 1 0 45448 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_59_494
timestamp 1644511149
transform 1 0 46552 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_502
timestamp 1644511149
transform 1 0 47288 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_59_505
timestamp 1644511149
transform 1 0 47564 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_59_513
timestamp 1644511149
transform 1 0 48300 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_519
timestamp 1644511149
transform 1 0 48852 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_540
timestamp 1644511149
transform 1 0 50784 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_59_552
timestamp 1644511149
transform 1 0 51888 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_59_556
timestamp 1644511149
transform 1 0 52256 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_565
timestamp 1644511149
transform 1 0 53084 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_59_572
timestamp 1644511149
transform 1 0 53728 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_59_578
timestamp 1644511149
transform 1 0 54280 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_590
timestamp 1644511149
transform 1 0 55384 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_59_602
timestamp 1644511149
transform 1 0 56488 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_59_614
timestamp 1644511149
transform 1 0 57592 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_59_617
timestamp 1644511149
transform 1 0 57868 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_59_621
timestamp 1644511149
transform 1 0 58236 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_3
timestamp 1644511149
transform 1 0 1380 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_15
timestamp 1644511149
transform 1 0 2484 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_60_27
timestamp 1644511149
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_29
timestamp 1644511149
transform 1 0 3772 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_41
timestamp 1644511149
transform 1 0 4876 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_53
timestamp 1644511149
transform 1 0 5980 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_60_68
timestamp 1644511149
transform 1 0 7360 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_78
timestamp 1644511149
transform 1 0 8280 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_60_87
timestamp 1644511149
transform 1 0 9108 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_93
timestamp 1644511149
transform 1 0 9660 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_107
timestamp 1644511149
transform 1 0 10948 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_116
timestamp 1644511149
transform 1 0 11776 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_127
timestamp 1644511149
transform 1 0 12788 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_133
timestamp 1644511149
transform 1 0 13340 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_139
timestamp 1644511149
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_141
timestamp 1644511149
transform 1 0 14076 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_153
timestamp 1644511149
transform 1 0 15180 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_157
timestamp 1644511149
transform 1 0 15548 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_163
timestamp 1644511149
transform 1 0 16100 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_169
timestamp 1644511149
transform 1 0 16652 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_175
timestamp 1644511149
transform 1 0 17204 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_192
timestamp 1644511149
transform 1 0 18768 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_60_197
timestamp 1644511149
transform 1 0 19228 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_209
timestamp 1644511149
transform 1 0 20332 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_226
timestamp 1644511149
transform 1 0 21896 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_236
timestamp 1644511149
transform 1 0 22816 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_242
timestamp 1644511149
transform 1 0 23368 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_60_248
timestamp 1644511149
transform 1 0 23920 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_60_253
timestamp 1644511149
transform 1 0 24380 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_269
timestamp 1644511149
transform 1 0 25852 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_281
timestamp 1644511149
transform 1 0 26956 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_60_293
timestamp 1644511149
transform 1 0 28060 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_60_300
timestamp 1644511149
transform 1 0 28704 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_309
timestamp 1644511149
transform 1 0 29532 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_321
timestamp 1644511149
transform 1 0 30636 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_333
timestamp 1644511149
transform 1 0 31740 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_345
timestamp 1644511149
transform 1 0 32844 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_60_357
timestamp 1644511149
transform 1 0 33948 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_363
timestamp 1644511149
transform 1 0 34500 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_372
timestamp 1644511149
transform 1 0 35328 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_384
timestamp 1644511149
transform 1 0 36432 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_60_392
timestamp 1644511149
transform 1 0 37168 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_60_400
timestamp 1644511149
transform 1 0 37904 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_60_412
timestamp 1644511149
transform 1 0 39008 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_60_421
timestamp 1644511149
transform 1 0 39836 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_433
timestamp 1644511149
transform 1 0 40940 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_445
timestamp 1644511149
transform 1 0 42044 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_464
timestamp 1644511149
transform 1 0 43792 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_477
timestamp 1644511149
transform 1 0 44988 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_489
timestamp 1644511149
transform 1 0 46092 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_501
timestamp 1644511149
transform 1 0 47196 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_60_518
timestamp 1644511149
transform 1 0 48760 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_60_525
timestamp 1644511149
transform 1 0 49404 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_60_531
timestamp 1644511149
transform 1 0 49956 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_535
timestamp 1644511149
transform 1 0 50324 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_547
timestamp 1644511149
transform 1 0 51428 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_559
timestamp 1644511149
transform 1 0 52532 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_563
timestamp 1644511149
transform 1 0 52900 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_571
timestamp 1644511149
transform 1 0 53636 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_60_583
timestamp 1644511149
transform 1 0 54740 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_60_587
timestamp 1644511149
transform 1 0 55108 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_60_589
timestamp 1644511149
transform 1 0 55292 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_60_601
timestamp 1644511149
transform 1 0 56396 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_60_613
timestamp 1644511149
transform 1 0 57500 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_60_621
timestamp 1644511149
transform 1 0 58236 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_3
timestamp 1644511149
transform 1 0 1380 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_15
timestamp 1644511149
transform 1 0 2484 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_27
timestamp 1644511149
transform 1 0 3588 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_39
timestamp 1644511149
transform 1 0 4692 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_51
timestamp 1644511149
transform 1 0 5796 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_55
timestamp 1644511149
transform 1 0 6164 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_61_64
timestamp 1644511149
transform 1 0 6992 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_61_79
timestamp 1644511149
transform 1 0 8372 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_86
timestamp 1644511149
transform 1 0 9016 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_92
timestamp 1644511149
transform 1 0 9568 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_98
timestamp 1644511149
transform 1 0 10120 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_110
timestamp 1644511149
transform 1 0 11224 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_61_113
timestamp 1644511149
transform 1 0 11500 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_120
timestamp 1644511149
transform 1 0 12144 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_126
timestamp 1644511149
transform 1 0 12696 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_138
timestamp 1644511149
transform 1 0 13800 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_150
timestamp 1644511149
transform 1 0 14904 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_162
timestamp 1644511149
transform 1 0 16008 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_61_169
timestamp 1644511149
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_181
timestamp 1644511149
transform 1 0 17756 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_61_189
timestamp 1644511149
transform 1 0 18492 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_61_197
timestamp 1644511149
transform 1 0 19228 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_207
timestamp 1644511149
transform 1 0 20148 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_219
timestamp 1644511149
transform 1 0 21252 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_61_223
timestamp 1644511149
transform 1 0 21620 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_225
timestamp 1644511149
transform 1 0 21804 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_237
timestamp 1644511149
transform 1 0 22908 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_243
timestamp 1644511149
transform 1 0 23460 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_255
timestamp 1644511149
transform 1 0 24564 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_267
timestamp 1644511149
transform 1 0 25668 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_279
timestamp 1644511149
transform 1 0 26772 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_281
timestamp 1644511149
transform 1 0 26956 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_293
timestamp 1644511149
transform 1 0 28060 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_300
timestamp 1644511149
transform 1 0 28704 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_61_311
timestamp 1644511149
transform 1 0 29716 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_317
timestamp 1644511149
transform 1 0 30268 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_329
timestamp 1644511149
transform 1 0 31372 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_335
timestamp 1644511149
transform 1 0 31924 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_337
timestamp 1644511149
transform 1 0 32108 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_61_346
timestamp 1644511149
transform 1 0 32936 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_358
timestamp 1644511149
transform 1 0 34040 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_370
timestamp 1644511149
transform 1 0 35144 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_382
timestamp 1644511149
transform 1 0 36248 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_390
timestamp 1644511149
transform 1 0 36984 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_61_393
timestamp 1644511149
transform 1 0 37260 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_405
timestamp 1644511149
transform 1 0 38364 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_417
timestamp 1644511149
transform 1 0 39468 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_423
timestamp 1644511149
transform 1 0 40020 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_61_426
timestamp 1644511149
transform 1 0 40296 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_432
timestamp 1644511149
transform 1 0 40848 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_435
timestamp 1644511149
transform 1 0 41124 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_61_447
timestamp 1644511149
transform 1 0 42228 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_61_449
timestamp 1644511149
transform 1 0 42412 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_461
timestamp 1644511149
transform 1 0 43516 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_61_473
timestamp 1644511149
transform 1 0 44620 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_61_490
timestamp 1644511149
transform 1 0 46184 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_61_502
timestamp 1644511149
transform 1 0 47288 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_61_505
timestamp 1644511149
transform 1 0 47564 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_517
timestamp 1644511149
transform 1 0 48668 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_61_526
timestamp 1644511149
transform 1 0 49496 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_538
timestamp 1644511149
transform 1 0 50600 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_61_550
timestamp 1644511149
transform 1 0 51704 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_61_558
timestamp 1644511149
transform 1 0 52440 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_61_561
timestamp 1644511149
transform 1 0 52716 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_573
timestamp 1644511149
transform 1 0 53820 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_585
timestamp 1644511149
transform 1 0 54924 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_61_597
timestamp 1644511149
transform 1 0 56028 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_61_609
timestamp 1644511149
transform 1 0 57132 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_61_615
timestamp 1644511149
transform 1 0 57684 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_61_617
timestamp 1644511149
transform 1 0 57868 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_61_621
timestamp 1644511149
transform 1 0 58236 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_7
timestamp 1644511149
transform 1 0 1748 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_19
timestamp 1644511149
transform 1 0 2852 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_27
timestamp 1644511149
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_29
timestamp 1644511149
transform 1 0 3772 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_41
timestamp 1644511149
transform 1 0 4876 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_53
timestamp 1644511149
transform 1 0 5980 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_62_61
timestamp 1644511149
transform 1 0 6716 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_66
timestamp 1644511149
transform 1 0 7176 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_70
timestamp 1644511149
transform 1 0 7544 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_73
timestamp 1644511149
transform 1 0 7820 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_80
timestamp 1644511149
transform 1 0 8464 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_90
timestamp 1644511149
transform 1 0 9384 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_96
timestamp 1644511149
transform 1 0 9936 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_108
timestamp 1644511149
transform 1 0 11040 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_120
timestamp 1644511149
transform 1 0 12144 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_132
timestamp 1644511149
transform 1 0 13248 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_62_141
timestamp 1644511149
transform 1 0 14076 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_153
timestamp 1644511149
transform 1 0 15180 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_165
timestamp 1644511149
transform 1 0 16284 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_177
timestamp 1644511149
transform 1 0 17388 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_189
timestamp 1644511149
transform 1 0 18492 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_195
timestamp 1644511149
transform 1 0 19044 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_203
timestamp 1644511149
transform 1 0 19780 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_62_215
timestamp 1644511149
transform 1 0 20884 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_225
timestamp 1644511149
transform 1 0 21804 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_234
timestamp 1644511149
transform 1 0 22632 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_62_242
timestamp 1644511149
transform 1 0 23368 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_62_248
timestamp 1644511149
transform 1 0 23920 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_62_258
timestamp 1644511149
transform 1 0 24840 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_62_270
timestamp 1644511149
transform 1 0 25944 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_62_276
timestamp 1644511149
transform 1 0 26496 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_62_288
timestamp 1644511149
transform 1 0 27600 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_296
timestamp 1644511149
transform 1 0 28336 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_300
timestamp 1644511149
transform 1 0 28704 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_62_316
timestamp 1644511149
transform 1 0 30176 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_320
timestamp 1644511149
transform 1 0 30544 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_324
timestamp 1644511149
transform 1 0 30912 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_334
timestamp 1644511149
transform 1 0 31832 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_62_345
timestamp 1644511149
transform 1 0 32844 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_354
timestamp 1644511149
transform 1 0 33672 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_62_362
timestamp 1644511149
transform 1 0 34408 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_62_365
timestamp 1644511149
transform 1 0 34684 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_373
timestamp 1644511149
transform 1 0 35420 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_396
timestamp 1644511149
transform 1 0 37536 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_62_400
timestamp 1644511149
transform 1 0 37904 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_408
timestamp 1644511149
transform 1 0 38640 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_62_414
timestamp 1644511149
transform 1 0 39192 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_62_443
timestamp 1644511149
transform 1 0 41860 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_449
timestamp 1644511149
transform 1 0 42412 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_62_472
timestamp 1644511149
transform 1 0 44528 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_62_477
timestamp 1644511149
transform 1 0 44988 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_485
timestamp 1644511149
transform 1 0 45724 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_62_508
timestamp 1644511149
transform 1 0 47840 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_62_523
timestamp 1644511149
transform 1 0 49220 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_62_531
timestamp 1644511149
transform 1 0 49956 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_533
timestamp 1644511149
transform 1 0 50140 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_545
timestamp 1644511149
transform 1 0 51244 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_557
timestamp 1644511149
transform 1 0 52348 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_569
timestamp 1644511149
transform 1 0 53452 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_62_581
timestamp 1644511149
transform 1 0 54556 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_62_587
timestamp 1644511149
transform 1 0 55108 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_62_589
timestamp 1644511149
transform 1 0 55292 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_62_601
timestamp 1644511149
transform 1 0 56396 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_62_613
timestamp 1644511149
transform 1 0 57500 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_62_621
timestamp 1644511149
transform 1 0 58236 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_7
timestamp 1644511149
transform 1 0 1748 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_19
timestamp 1644511149
transform 1 0 2852 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_33
timestamp 1644511149
transform 1 0 4140 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_52
timestamp 1644511149
transform 1 0 5888 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_59
timestamp 1644511149
transform 1 0 6532 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_63_72
timestamp 1644511149
transform 1 0 7728 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_82
timestamp 1644511149
transform 1 0 8648 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_88
timestamp 1644511149
transform 1 0 9200 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_100
timestamp 1644511149
transform 1 0 10304 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_113
timestamp 1644511149
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_125
timestamp 1644511149
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_137
timestamp 1644511149
transform 1 0 13708 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_143
timestamp 1644511149
transform 1 0 14260 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_155
timestamp 1644511149
transform 1 0 15364 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_167
timestamp 1644511149
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_169
timestamp 1644511149
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_181
timestamp 1644511149
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_193
timestamp 1644511149
transform 1 0 18860 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_201
timestamp 1644511149
transform 1 0 19596 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_215
timestamp 1644511149
transform 1 0 20884 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_223
timestamp 1644511149
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_225
timestamp 1644511149
transform 1 0 21804 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_229
timestamp 1644511149
transform 1 0 22172 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_63_237
timestamp 1644511149
transform 1 0 22908 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_63_245
timestamp 1644511149
transform 1 0 23644 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_63_260
timestamp 1644511149
transform 1 0 25024 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_266
timestamp 1644511149
transform 1 0 25576 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_275
timestamp 1644511149
transform 1 0 26404 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_279
timestamp 1644511149
transform 1 0 26772 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_294
timestamp 1644511149
transform 1 0 28152 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_305
timestamp 1644511149
transform 1 0 29164 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_313
timestamp 1644511149
transform 1 0 29900 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_318
timestamp 1644511149
transform 1 0 30360 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_330
timestamp 1644511149
transform 1 0 31464 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_63_344
timestamp 1644511149
transform 1 0 32752 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_356
timestamp 1644511149
transform 1 0 33856 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_63_364
timestamp 1644511149
transform 1 0 34592 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_370
timestamp 1644511149
transform 1 0 35144 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_63_381
timestamp 1644511149
transform 1 0 36156 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_389
timestamp 1644511149
transform 1 0 36892 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_63_393
timestamp 1644511149
transform 1 0 37260 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_63_397
timestamp 1644511149
transform 1 0 37628 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_403
timestamp 1644511149
transform 1 0 38180 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_411
timestamp 1644511149
transform 1 0 38916 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_422
timestamp 1644511149
transform 1 0 39928 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_63_431
timestamp 1644511149
transform 1 0 40756 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_63_444
timestamp 1644511149
transform 1 0 41952 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_63_449
timestamp 1644511149
transform 1 0 42412 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_457
timestamp 1644511149
transform 1 0 43148 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_466
timestamp 1644511149
transform 1 0 43976 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_63_500
timestamp 1644511149
transform 1 0 47104 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_510
timestamp 1644511149
transform 1 0 48024 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_516
timestamp 1644511149
transform 1 0 48576 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_63_522
timestamp 1644511149
transform 1 0 49128 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_63_534
timestamp 1644511149
transform 1 0 50232 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_63_537
timestamp 1644511149
transform 1 0 50508 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_63_549
timestamp 1644511149
transform 1 0 51612 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_63_557
timestamp 1644511149
transform 1 0 52348 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_63_561
timestamp 1644511149
transform 1 0 52716 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_573
timestamp 1644511149
transform 1 0 53820 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_63_585
timestamp 1644511149
transform 1 0 54924 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_63_597
timestamp 1644511149
transform 1 0 56028 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_63_603
timestamp 1644511149
transform 1 0 56580 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_63_606
timestamp 1644511149
transform 1 0 56856 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_612
timestamp 1644511149
transform 1 0 57408 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_63_621
timestamp 1644511149
transform 1 0 58236 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_7
timestamp 1644511149
transform 1 0 1748 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_15
timestamp 1644511149
transform 1 0 2484 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_21
timestamp 1644511149
transform 1 0 3036 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_27
timestamp 1644511149
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_29
timestamp 1644511149
transform 1 0 3772 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_37
timestamp 1644511149
transform 1 0 4508 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_49
timestamp 1644511149
transform 1 0 5612 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_55
timestamp 1644511149
transform 1 0 6164 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_61
timestamp 1644511149
transform 1 0 6716 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_69
timestamp 1644511149
transform 1 0 7452 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_76
timestamp 1644511149
transform 1 0 8096 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_85
timestamp 1644511149
transform 1 0 8924 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_90
timestamp 1644511149
transform 1 0 9384 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_98
timestamp 1644511149
transform 1 0 10120 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_110
timestamp 1644511149
transform 1 0 11224 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_64_113
timestamp 1644511149
transform 1 0 11500 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_118
timestamp 1644511149
transform 1 0 11960 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_126
timestamp 1644511149
transform 1 0 12696 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_138
timestamp 1644511149
transform 1 0 13800 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_141
timestamp 1644511149
transform 1 0 14076 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_153
timestamp 1644511149
transform 1 0 15180 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_161
timestamp 1644511149
transform 1 0 15916 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_164
timestamp 1644511149
transform 1 0 16192 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_173
timestamp 1644511149
transform 1 0 17020 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_189
timestamp 1644511149
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_195
timestamp 1644511149
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_64_197
timestamp 1644511149
transform 1 0 19228 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_202
timestamp 1644511149
transform 1 0 19688 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_215
timestamp 1644511149
transform 1 0 20884 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_223
timestamp 1644511149
transform 1 0 21620 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_225
timestamp 1644511149
transform 1 0 21804 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_233
timestamp 1644511149
transform 1 0 22540 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_239
timestamp 1644511149
transform 1 0 23092 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_245
timestamp 1644511149
transform 1 0 23644 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_248
timestamp 1644511149
transform 1 0 23920 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_257
timestamp 1644511149
transform 1 0 24748 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_64_265
timestamp 1644511149
transform 1 0 25484 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_272
timestamp 1644511149
transform 1 0 26128 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_64_281
timestamp 1644511149
transform 1 0 26956 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_289
timestamp 1644511149
transform 1 0 27692 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_293
timestamp 1644511149
transform 1 0 28060 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_301
timestamp 1644511149
transform 1 0 28796 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_307
timestamp 1644511149
transform 1 0 29348 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_64_309
timestamp 1644511149
transform 1 0 29532 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_314
timestamp 1644511149
transform 1 0 29992 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_322
timestamp 1644511149
transform 1 0 30728 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_64_334
timestamp 1644511149
transform 1 0 31832 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_64_337
timestamp 1644511149
transform 1 0 32108 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_64_343
timestamp 1644511149
transform 1 0 32660 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_64_353
timestamp 1644511149
transform 1 0 33580 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_360
timestamp 1644511149
transform 1 0 34224 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_365
timestamp 1644511149
transform 1 0 34684 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_371
timestamp 1644511149
transform 1 0 35236 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_382
timestamp 1644511149
transform 1 0 36248 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_64_390
timestamp 1644511149
transform 1 0 36984 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_64_393
timestamp 1644511149
transform 1 0 37260 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_403
timestamp 1644511149
transform 1 0 38180 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_409
timestamp 1644511149
transform 1 0 38732 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_415
timestamp 1644511149
transform 1 0 39284 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_64_419
timestamp 1644511149
transform 1 0 39652 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_425
timestamp 1644511149
transform 1 0 40204 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_433
timestamp 1644511149
transform 1 0 40940 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_64_444
timestamp 1644511149
transform 1 0 41952 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_454
timestamp 1644511149
transform 1 0 42872 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_460
timestamp 1644511149
transform 1 0 43424 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_64_472
timestamp 1644511149
transform 1 0 44528 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_477
timestamp 1644511149
transform 1 0 44988 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_64_489
timestamp 1644511149
transform 1 0 46092 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_64_497
timestamp 1644511149
transform 1 0 46828 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_503
timestamp 1644511149
transform 1 0 47380 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_505
timestamp 1644511149
transform 1 0 47564 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_64_515
timestamp 1644511149
transform 1 0 48484 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_64_525
timestamp 1644511149
transform 1 0 49404 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_531
timestamp 1644511149
transform 1 0 49956 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_533
timestamp 1644511149
transform 1 0 50140 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_543
timestamp 1644511149
transform 1 0 51060 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_64_551
timestamp 1644511149
transform 1 0 51796 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_556
timestamp 1644511149
transform 1 0 52256 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_64_565
timestamp 1644511149
transform 1 0 53084 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_64_581
timestamp 1644511149
transform 1 0 54556 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_64_587
timestamp 1644511149
transform 1 0 55108 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_64_589
timestamp 1644511149
transform 1 0 55292 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_64_594
timestamp 1644511149
transform 1 0 55752 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_64_607
timestamp 1644511149
transform 1 0 56948 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_64_615
timestamp 1644511149
transform 1 0 57684 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_64_621
timestamp 1644511149
transform 1 0 58236 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1644511149
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1644511149
transform -1 0 58880 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1644511149
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1644511149
transform -1 0 58880 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1644511149
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1644511149
transform -1 0 58880 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1644511149
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1644511149
transform -1 0 58880 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1644511149
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1644511149
transform -1 0 58880 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1644511149
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1644511149
transform -1 0 58880 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1644511149
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1644511149
transform -1 0 58880 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1644511149
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1644511149
transform -1 0 58880 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1644511149
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1644511149
transform -1 0 58880 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1644511149
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1644511149
transform -1 0 58880 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1644511149
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1644511149
transform -1 0 58880 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1644511149
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1644511149
transform -1 0 58880 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1644511149
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1644511149
transform -1 0 58880 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1644511149
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1644511149
transform -1 0 58880 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1644511149
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1644511149
transform -1 0 58880 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1644511149
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1644511149
transform -1 0 58880 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1644511149
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1644511149
transform -1 0 58880 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1644511149
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1644511149
transform -1 0 58880 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1644511149
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1644511149
transform -1 0 58880 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1644511149
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1644511149
transform -1 0 58880 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1644511149
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1644511149
transform -1 0 58880 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1644511149
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1644511149
transform -1 0 58880 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1644511149
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1644511149
transform -1 0 58880 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1644511149
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1644511149
transform -1 0 58880 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1644511149
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1644511149
transform -1 0 58880 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1644511149
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1644511149
transform -1 0 58880 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1644511149
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1644511149
transform -1 0 58880 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1644511149
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1644511149
transform -1 0 58880 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1644511149
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1644511149
transform -1 0 58880 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1644511149
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1644511149
transform -1 0 58880 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1644511149
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1644511149
transform -1 0 58880 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1644511149
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1644511149
transform -1 0 58880 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1644511149
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1644511149
transform -1 0 58880 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1644511149
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1644511149
transform -1 0 58880 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1644511149
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1644511149
transform -1 0 58880 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1644511149
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1644511149
transform -1 0 58880 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1644511149
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1644511149
transform -1 0 58880 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1644511149
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1644511149
transform -1 0 58880 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1644511149
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1644511149
transform -1 0 58880 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1644511149
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1644511149
transform -1 0 58880 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1644511149
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1644511149
transform -1 0 58880 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1644511149
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1644511149
transform -1 0 58880 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1644511149
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1644511149
transform -1 0 58880 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1644511149
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1644511149
transform -1 0 58880 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1644511149
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1644511149
transform -1 0 58880 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1644511149
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1644511149
transform -1 0 58880 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1644511149
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1644511149
transform -1 0 58880 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1644511149
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1644511149
transform -1 0 58880 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1644511149
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1644511149
transform -1 0 58880 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1644511149
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1644511149
transform -1 0 58880 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1644511149
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1644511149
transform -1 0 58880 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1644511149
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1644511149
transform -1 0 58880 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1644511149
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1644511149
transform -1 0 58880 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1644511149
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1644511149
transform -1 0 58880 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1644511149
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1644511149
transform -1 0 58880 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1644511149
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1644511149
transform -1 0 58880 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1644511149
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1644511149
transform -1 0 58880 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1644511149
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1644511149
transform -1 0 58880 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1644511149
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1644511149
transform -1 0 58880 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1644511149
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1644511149
transform -1 0 58880 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1644511149
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1644511149
transform -1 0 58880 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1644511149
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1644511149
transform -1 0 58880 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1644511149
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1644511149
transform -1 0 58880 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1644511149
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1644511149
transform -1 0 58880 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1644511149
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1644511149
transform -1 0 58880 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130 pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1644511149
transform 1 0 6256 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1644511149
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1644511149
transform 1 0 11408 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1644511149
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1644511149
transform 1 0 16560 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1644511149
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1644511149
transform 1 0 21712 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1644511149
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1644511149
transform 1 0 26864 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1644511149
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1644511149
transform 1 0 32016 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1644511149
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1644511149
transform 1 0 37168 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1644511149
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1644511149
transform 1 0 42320 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1644511149
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1644511149
transform 1 0 47472 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1644511149
transform 1 0 50048 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1644511149
transform 1 0 52624 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1644511149
transform 1 0 55200 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1644511149
transform 1 0 57776 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1644511149
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1644511149
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1644511149
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1644511149
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1644511149
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1644511149
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1644511149
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1644511149
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1644511149
transform 1 0 47472 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1644511149
transform 1 0 52624 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1644511149
transform 1 0 57776 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1644511149
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1644511149
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1644511149
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1644511149
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1644511149
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1644511149
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1644511149
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1644511149
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1644511149
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1644511149
transform 1 0 50048 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1644511149
transform 1 0 55200 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1644511149
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1644511149
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1644511149
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1644511149
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1644511149
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1644511149
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1644511149
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1644511149
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1644511149
transform 1 0 47472 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1644511149
transform 1 0 52624 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1644511149
transform 1 0 57776 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1644511149
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1644511149
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1644511149
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1644511149
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1644511149
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1644511149
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1644511149
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1644511149
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1644511149
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1644511149
transform 1 0 50048 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1644511149
transform 1 0 55200 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1644511149
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1644511149
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1644511149
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1644511149
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1644511149
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1644511149
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1644511149
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1644511149
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1644511149
transform 1 0 47472 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1644511149
transform 1 0 52624 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1644511149
transform 1 0 57776 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1644511149
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1644511149
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1644511149
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1644511149
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1644511149
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1644511149
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1644511149
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1644511149
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1644511149
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1644511149
transform 1 0 50048 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1644511149
transform 1 0 55200 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1644511149
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1644511149
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1644511149
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1644511149
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1644511149
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1644511149
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1644511149
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1644511149
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1644511149
transform 1 0 47472 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1644511149
transform 1 0 52624 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1644511149
transform 1 0 57776 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1644511149
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1644511149
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1644511149
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1644511149
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1644511149
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1644511149
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1644511149
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1644511149
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1644511149
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1644511149
transform 1 0 50048 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1644511149
transform 1 0 55200 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1644511149
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1644511149
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1644511149
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1644511149
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1644511149
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1644511149
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1644511149
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1644511149
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1644511149
transform 1 0 47472 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1644511149
transform 1 0 52624 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1644511149
transform 1 0 57776 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1644511149
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1644511149
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1644511149
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1644511149
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1644511149
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1644511149
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1644511149
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1644511149
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1644511149
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1644511149
transform 1 0 50048 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1644511149
transform 1 0 55200 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1644511149
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1644511149
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1644511149
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1644511149
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1644511149
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1644511149
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1644511149
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1644511149
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1644511149
transform 1 0 47472 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1644511149
transform 1 0 52624 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1644511149
transform 1 0 57776 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1644511149
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1644511149
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1644511149
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1644511149
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1644511149
transform 1 0 24288 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1644511149
transform 1 0 29440 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1644511149
transform 1 0 34592 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1644511149
transform 1 0 39744 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1644511149
transform 1 0 44896 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1644511149
transform 1 0 50048 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1644511149
transform 1 0 55200 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1644511149
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1644511149
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1644511149
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1644511149
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1644511149
transform 1 0 26864 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1644511149
transform 1 0 32016 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1644511149
transform 1 0 37168 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1644511149
transform 1 0 42320 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1644511149
transform 1 0 47472 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1644511149
transform 1 0 52624 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1644511149
transform 1 0 57776 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1644511149
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1644511149
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1644511149
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1644511149
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1644511149
transform 1 0 24288 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1644511149
transform 1 0 29440 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1644511149
transform 1 0 34592 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1644511149
transform 1 0 39744 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1644511149
transform 1 0 44896 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1644511149
transform 1 0 50048 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1644511149
transform 1 0 55200 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1644511149
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1644511149
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1644511149
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1644511149
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1644511149
transform 1 0 26864 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1644511149
transform 1 0 32016 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1644511149
transform 1 0 37168 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1644511149
transform 1 0 42320 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1644511149
transform 1 0 47472 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1644511149
transform 1 0 52624 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1644511149
transform 1 0 57776 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1644511149
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1644511149
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1644511149
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1644511149
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1644511149
transform 1 0 24288 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1644511149
transform 1 0 29440 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1644511149
transform 1 0 34592 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1644511149
transform 1 0 39744 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1644511149
transform 1 0 44896 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1644511149
transform 1 0 50048 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1644511149
transform 1 0 55200 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1644511149
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1644511149
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1644511149
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1644511149
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1644511149
transform 1 0 26864 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1644511149
transform 1 0 32016 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1644511149
transform 1 0 37168 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1644511149
transform 1 0 42320 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1644511149
transform 1 0 47472 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1644511149
transform 1 0 52624 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1644511149
transform 1 0 57776 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1644511149
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1644511149
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1644511149
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1644511149
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1644511149
transform 1 0 24288 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1644511149
transform 1 0 29440 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1644511149
transform 1 0 34592 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1644511149
transform 1 0 39744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1644511149
transform 1 0 44896 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1644511149
transform 1 0 50048 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1644511149
transform 1 0 55200 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1644511149
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1644511149
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1644511149
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1644511149
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1644511149
transform 1 0 26864 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1644511149
transform 1 0 32016 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1644511149
transform 1 0 37168 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1644511149
transform 1 0 42320 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1644511149
transform 1 0 47472 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1644511149
transform 1 0 52624 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1644511149
transform 1 0 57776 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1644511149
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1644511149
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1644511149
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1644511149
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1644511149
transform 1 0 24288 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1644511149
transform 1 0 29440 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1644511149
transform 1 0 34592 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1644511149
transform 1 0 39744 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1644511149
transform 1 0 44896 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1644511149
transform 1 0 50048 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1644511149
transform 1 0 55200 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1644511149
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1644511149
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1644511149
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1644511149
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1644511149
transform 1 0 26864 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1644511149
transform 1 0 32016 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1644511149
transform 1 0 37168 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1644511149
transform 1 0 42320 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1644511149
transform 1 0 47472 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1644511149
transform 1 0 52624 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1644511149
transform 1 0 57776 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1644511149
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1644511149
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1644511149
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1644511149
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1644511149
transform 1 0 24288 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1644511149
transform 1 0 29440 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1644511149
transform 1 0 34592 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1644511149
transform 1 0 39744 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1644511149
transform 1 0 44896 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1644511149
transform 1 0 50048 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1644511149
transform 1 0 55200 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1644511149
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1644511149
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1644511149
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1644511149
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1644511149
transform 1 0 26864 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1644511149
transform 1 0 32016 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1644511149
transform 1 0 37168 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1644511149
transform 1 0 42320 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1644511149
transform 1 0 47472 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1644511149
transform 1 0 52624 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1644511149
transform 1 0 57776 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1644511149
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1644511149
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1644511149
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1644511149
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1644511149
transform 1 0 24288 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1644511149
transform 1 0 29440 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1644511149
transform 1 0 34592 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1644511149
transform 1 0 39744 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1644511149
transform 1 0 44896 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1644511149
transform 1 0 50048 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1644511149
transform 1 0 55200 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1644511149
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1644511149
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1644511149
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1644511149
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1644511149
transform 1 0 26864 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1644511149
transform 1 0 32016 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1644511149
transform 1 0 37168 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1644511149
transform 1 0 42320 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1644511149
transform 1 0 47472 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1644511149
transform 1 0 52624 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1644511149
transform 1 0 57776 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1644511149
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1644511149
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1644511149
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1644511149
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1644511149
transform 1 0 24288 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1644511149
transform 1 0 29440 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1644511149
transform 1 0 34592 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1644511149
transform 1 0 39744 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1644511149
transform 1 0 44896 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1644511149
transform 1 0 50048 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1644511149
transform 1 0 55200 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1644511149
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1644511149
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1644511149
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1644511149
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1644511149
transform 1 0 26864 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1644511149
transform 1 0 32016 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1644511149
transform 1 0 37168 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1644511149
transform 1 0 42320 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1644511149
transform 1 0 47472 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1644511149
transform 1 0 52624 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1644511149
transform 1 0 57776 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1644511149
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1644511149
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1644511149
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1644511149
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1644511149
transform 1 0 24288 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1644511149
transform 1 0 29440 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1644511149
transform 1 0 34592 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1644511149
transform 1 0 39744 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1644511149
transform 1 0 44896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1644511149
transform 1 0 50048 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1644511149
transform 1 0 55200 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1644511149
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1644511149
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1644511149
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1644511149
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1644511149
transform 1 0 26864 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1644511149
transform 1 0 32016 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1644511149
transform 1 0 37168 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1644511149
transform 1 0 42320 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1644511149
transform 1 0 47472 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1644511149
transform 1 0 52624 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1644511149
transform 1 0 57776 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1644511149
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1644511149
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1644511149
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1644511149
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1644511149
transform 1 0 24288 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_476
timestamp 1644511149
transform 1 0 29440 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_477
timestamp 1644511149
transform 1 0 34592 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_478
timestamp 1644511149
transform 1 0 39744 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_479
timestamp 1644511149
transform 1 0 44896 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_480
timestamp 1644511149
transform 1 0 50048 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_481
timestamp 1644511149
transform 1 0 55200 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_482
timestamp 1644511149
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_483
timestamp 1644511149
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_484
timestamp 1644511149
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_485
timestamp 1644511149
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_486
timestamp 1644511149
transform 1 0 26864 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_487
timestamp 1644511149
transform 1 0 32016 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_488
timestamp 1644511149
transform 1 0 37168 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_489
timestamp 1644511149
transform 1 0 42320 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_490
timestamp 1644511149
transform 1 0 47472 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_491
timestamp 1644511149
transform 1 0 52624 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_492
timestamp 1644511149
transform 1 0 57776 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_493
timestamp 1644511149
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_494
timestamp 1644511149
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_495
timestamp 1644511149
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_496
timestamp 1644511149
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_497
timestamp 1644511149
transform 1 0 24288 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_498
timestamp 1644511149
transform 1 0 29440 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_499
timestamp 1644511149
transform 1 0 34592 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_500
timestamp 1644511149
transform 1 0 39744 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_501
timestamp 1644511149
transform 1 0 44896 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_502
timestamp 1644511149
transform 1 0 50048 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_503
timestamp 1644511149
transform 1 0 55200 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_504
timestamp 1644511149
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_505
timestamp 1644511149
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_506
timestamp 1644511149
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_507
timestamp 1644511149
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_508
timestamp 1644511149
transform 1 0 26864 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_509
timestamp 1644511149
transform 1 0 32016 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_510
timestamp 1644511149
transform 1 0 37168 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_511
timestamp 1644511149
transform 1 0 42320 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_512
timestamp 1644511149
transform 1 0 47472 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_513
timestamp 1644511149
transform 1 0 52624 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_514
timestamp 1644511149
transform 1 0 57776 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_515
timestamp 1644511149
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_516
timestamp 1644511149
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_517
timestamp 1644511149
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_518
timestamp 1644511149
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_519
timestamp 1644511149
transform 1 0 24288 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_520
timestamp 1644511149
transform 1 0 29440 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_521
timestamp 1644511149
transform 1 0 34592 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_522
timestamp 1644511149
transform 1 0 39744 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_523
timestamp 1644511149
transform 1 0 44896 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_524
timestamp 1644511149
transform 1 0 50048 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_525
timestamp 1644511149
transform 1 0 55200 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_526
timestamp 1644511149
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_527
timestamp 1644511149
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_528
timestamp 1644511149
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_529
timestamp 1644511149
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_530
timestamp 1644511149
transform 1 0 26864 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_531
timestamp 1644511149
transform 1 0 32016 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_532
timestamp 1644511149
transform 1 0 37168 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_533
timestamp 1644511149
transform 1 0 42320 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_534
timestamp 1644511149
transform 1 0 47472 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_535
timestamp 1644511149
transform 1 0 52624 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_536
timestamp 1644511149
transform 1 0 57776 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_537
timestamp 1644511149
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_538
timestamp 1644511149
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_539
timestamp 1644511149
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_540
timestamp 1644511149
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_541
timestamp 1644511149
transform 1 0 24288 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_542
timestamp 1644511149
transform 1 0 29440 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_543
timestamp 1644511149
transform 1 0 34592 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_544
timestamp 1644511149
transform 1 0 39744 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_545
timestamp 1644511149
transform 1 0 44896 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_546
timestamp 1644511149
transform 1 0 50048 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_547
timestamp 1644511149
transform 1 0 55200 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_548
timestamp 1644511149
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_549
timestamp 1644511149
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_550
timestamp 1644511149
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_551
timestamp 1644511149
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_552
timestamp 1644511149
transform 1 0 26864 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_553
timestamp 1644511149
transform 1 0 32016 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_554
timestamp 1644511149
transform 1 0 37168 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_555
timestamp 1644511149
transform 1 0 42320 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_556
timestamp 1644511149
transform 1 0 47472 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_557
timestamp 1644511149
transform 1 0 52624 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_558
timestamp 1644511149
transform 1 0 57776 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_559
timestamp 1644511149
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_560
timestamp 1644511149
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_561
timestamp 1644511149
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_562
timestamp 1644511149
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_563
timestamp 1644511149
transform 1 0 24288 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_564
timestamp 1644511149
transform 1 0 29440 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_565
timestamp 1644511149
transform 1 0 34592 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_566
timestamp 1644511149
transform 1 0 39744 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_567
timestamp 1644511149
transform 1 0 44896 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_568
timestamp 1644511149
transform 1 0 50048 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_569
timestamp 1644511149
transform 1 0 55200 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_570
timestamp 1644511149
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_571
timestamp 1644511149
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_572
timestamp 1644511149
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_573
timestamp 1644511149
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_574
timestamp 1644511149
transform 1 0 26864 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_575
timestamp 1644511149
transform 1 0 32016 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_576
timestamp 1644511149
transform 1 0 37168 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_577
timestamp 1644511149
transform 1 0 42320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_578
timestamp 1644511149
transform 1 0 47472 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_579
timestamp 1644511149
transform 1 0 52624 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_580
timestamp 1644511149
transform 1 0 57776 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_581
timestamp 1644511149
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_582
timestamp 1644511149
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_583
timestamp 1644511149
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_584
timestamp 1644511149
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_585
timestamp 1644511149
transform 1 0 24288 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_586
timestamp 1644511149
transform 1 0 29440 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_587
timestamp 1644511149
transform 1 0 34592 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_588
timestamp 1644511149
transform 1 0 39744 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_589
timestamp 1644511149
transform 1 0 44896 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_590
timestamp 1644511149
transform 1 0 50048 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_591
timestamp 1644511149
transform 1 0 55200 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_592
timestamp 1644511149
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_593
timestamp 1644511149
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_594
timestamp 1644511149
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_595
timestamp 1644511149
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_596
timestamp 1644511149
transform 1 0 26864 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_597
timestamp 1644511149
transform 1 0 32016 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_598
timestamp 1644511149
transform 1 0 37168 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_599
timestamp 1644511149
transform 1 0 42320 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_600
timestamp 1644511149
transform 1 0 47472 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_601
timestamp 1644511149
transform 1 0 52624 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_602
timestamp 1644511149
transform 1 0 57776 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_603
timestamp 1644511149
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_604
timestamp 1644511149
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_605
timestamp 1644511149
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_606
timestamp 1644511149
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_607
timestamp 1644511149
transform 1 0 24288 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_608
timestamp 1644511149
transform 1 0 29440 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_609
timestamp 1644511149
transform 1 0 34592 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_610
timestamp 1644511149
transform 1 0 39744 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_611
timestamp 1644511149
transform 1 0 44896 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_612
timestamp 1644511149
transform 1 0 50048 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_613
timestamp 1644511149
transform 1 0 55200 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_614
timestamp 1644511149
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_615
timestamp 1644511149
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_616
timestamp 1644511149
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_617
timestamp 1644511149
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_618
timestamp 1644511149
transform 1 0 26864 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_619
timestamp 1644511149
transform 1 0 32016 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_620
timestamp 1644511149
transform 1 0 37168 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_621
timestamp 1644511149
transform 1 0 42320 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_622
timestamp 1644511149
transform 1 0 47472 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_623
timestamp 1644511149
transform 1 0 52624 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_624
timestamp 1644511149
transform 1 0 57776 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_625
timestamp 1644511149
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_626
timestamp 1644511149
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_627
timestamp 1644511149
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_628
timestamp 1644511149
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_629
timestamp 1644511149
transform 1 0 24288 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_630
timestamp 1644511149
transform 1 0 29440 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_631
timestamp 1644511149
transform 1 0 34592 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_632
timestamp 1644511149
transform 1 0 39744 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_633
timestamp 1644511149
transform 1 0 44896 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_634
timestamp 1644511149
transform 1 0 50048 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_635
timestamp 1644511149
transform 1 0 55200 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_636
timestamp 1644511149
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_637
timestamp 1644511149
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_638
timestamp 1644511149
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_639
timestamp 1644511149
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_640
timestamp 1644511149
transform 1 0 26864 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_641
timestamp 1644511149
transform 1 0 32016 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_642
timestamp 1644511149
transform 1 0 37168 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_643
timestamp 1644511149
transform 1 0 42320 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_644
timestamp 1644511149
transform 1 0 47472 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_645
timestamp 1644511149
transform 1 0 52624 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_646
timestamp 1644511149
transform 1 0 57776 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_647
timestamp 1644511149
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_648
timestamp 1644511149
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_649
timestamp 1644511149
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_650
timestamp 1644511149
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_651
timestamp 1644511149
transform 1 0 24288 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_652
timestamp 1644511149
transform 1 0 29440 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_653
timestamp 1644511149
transform 1 0 34592 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_654
timestamp 1644511149
transform 1 0 39744 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_655
timestamp 1644511149
transform 1 0 44896 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_656
timestamp 1644511149
transform 1 0 50048 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_657
timestamp 1644511149
transform 1 0 55200 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_658
timestamp 1644511149
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_659
timestamp 1644511149
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_660
timestamp 1644511149
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_661
timestamp 1644511149
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_662
timestamp 1644511149
transform 1 0 26864 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_663
timestamp 1644511149
transform 1 0 32016 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_664
timestamp 1644511149
transform 1 0 37168 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_665
timestamp 1644511149
transform 1 0 42320 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_666
timestamp 1644511149
transform 1 0 47472 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_667
timestamp 1644511149
transform 1 0 52624 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_668
timestamp 1644511149
transform 1 0 57776 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_669
timestamp 1644511149
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_670
timestamp 1644511149
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_671
timestamp 1644511149
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_672
timestamp 1644511149
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_673
timestamp 1644511149
transform 1 0 24288 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_674
timestamp 1644511149
transform 1 0 29440 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_675
timestamp 1644511149
transform 1 0 34592 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_676
timestamp 1644511149
transform 1 0 39744 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_677
timestamp 1644511149
transform 1 0 44896 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_678
timestamp 1644511149
transform 1 0 50048 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_679
timestamp 1644511149
transform 1 0 55200 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_680
timestamp 1644511149
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_681
timestamp 1644511149
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_682
timestamp 1644511149
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_683
timestamp 1644511149
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_684
timestamp 1644511149
transform 1 0 26864 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_685
timestamp 1644511149
transform 1 0 32016 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_686
timestamp 1644511149
transform 1 0 37168 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_687
timestamp 1644511149
transform 1 0 42320 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_688
timestamp 1644511149
transform 1 0 47472 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_689
timestamp 1644511149
transform 1 0 52624 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_690
timestamp 1644511149
transform 1 0 57776 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_691
timestamp 1644511149
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_692
timestamp 1644511149
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_693
timestamp 1644511149
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_694
timestamp 1644511149
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_695
timestamp 1644511149
transform 1 0 24288 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_696
timestamp 1644511149
transform 1 0 29440 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_697
timestamp 1644511149
transform 1 0 34592 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_698
timestamp 1644511149
transform 1 0 39744 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_699
timestamp 1644511149
transform 1 0 44896 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_700
timestamp 1644511149
transform 1 0 50048 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_701
timestamp 1644511149
transform 1 0 55200 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_702
timestamp 1644511149
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_703
timestamp 1644511149
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_704
timestamp 1644511149
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_705
timestamp 1644511149
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_706
timestamp 1644511149
transform 1 0 26864 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_707
timestamp 1644511149
transform 1 0 32016 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_708
timestamp 1644511149
transform 1 0 37168 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_709
timestamp 1644511149
transform 1 0 42320 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_710
timestamp 1644511149
transform 1 0 47472 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_711
timestamp 1644511149
transform 1 0 52624 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_712
timestamp 1644511149
transform 1 0 57776 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_713
timestamp 1644511149
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_714
timestamp 1644511149
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_715
timestamp 1644511149
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_716
timestamp 1644511149
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_717
timestamp 1644511149
transform 1 0 24288 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_718
timestamp 1644511149
transform 1 0 29440 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_719
timestamp 1644511149
transform 1 0 34592 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_720
timestamp 1644511149
transform 1 0 39744 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_721
timestamp 1644511149
transform 1 0 44896 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_722
timestamp 1644511149
transform 1 0 50048 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_723
timestamp 1644511149
transform 1 0 55200 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_724
timestamp 1644511149
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_725
timestamp 1644511149
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_726
timestamp 1644511149
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_727
timestamp 1644511149
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_728
timestamp 1644511149
transform 1 0 26864 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_729
timestamp 1644511149
transform 1 0 32016 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_730
timestamp 1644511149
transform 1 0 37168 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_731
timestamp 1644511149
transform 1 0 42320 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_732
timestamp 1644511149
transform 1 0 47472 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_733
timestamp 1644511149
transform 1 0 52624 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_734
timestamp 1644511149
transform 1 0 57776 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_735
timestamp 1644511149
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_736
timestamp 1644511149
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_737
timestamp 1644511149
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_738
timestamp 1644511149
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_739
timestamp 1644511149
transform 1 0 24288 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_740
timestamp 1644511149
transform 1 0 29440 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_741
timestamp 1644511149
transform 1 0 34592 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_742
timestamp 1644511149
transform 1 0 39744 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_743
timestamp 1644511149
transform 1 0 44896 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_744
timestamp 1644511149
transform 1 0 50048 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_745
timestamp 1644511149
transform 1 0 55200 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_746
timestamp 1644511149
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_747
timestamp 1644511149
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_748
timestamp 1644511149
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_749
timestamp 1644511149
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_750
timestamp 1644511149
transform 1 0 26864 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_751
timestamp 1644511149
transform 1 0 32016 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_752
timestamp 1644511149
transform 1 0 37168 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_753
timestamp 1644511149
transform 1 0 42320 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_754
timestamp 1644511149
transform 1 0 47472 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_755
timestamp 1644511149
transform 1 0 52624 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_756
timestamp 1644511149
transform 1 0 57776 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_757
timestamp 1644511149
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_758
timestamp 1644511149
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_759
timestamp 1644511149
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_760
timestamp 1644511149
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_761
timestamp 1644511149
transform 1 0 24288 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_762
timestamp 1644511149
transform 1 0 29440 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_763
timestamp 1644511149
transform 1 0 34592 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_764
timestamp 1644511149
transform 1 0 39744 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_765
timestamp 1644511149
transform 1 0 44896 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_766
timestamp 1644511149
transform 1 0 50048 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_767
timestamp 1644511149
transform 1 0 55200 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_768
timestamp 1644511149
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_769
timestamp 1644511149
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_770
timestamp 1644511149
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_771
timestamp 1644511149
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_772
timestamp 1644511149
transform 1 0 26864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_773
timestamp 1644511149
transform 1 0 32016 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_774
timestamp 1644511149
transform 1 0 37168 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_775
timestamp 1644511149
transform 1 0 42320 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_776
timestamp 1644511149
transform 1 0 47472 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_777
timestamp 1644511149
transform 1 0 52624 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_778
timestamp 1644511149
transform 1 0 57776 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_779
timestamp 1644511149
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_780
timestamp 1644511149
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_781
timestamp 1644511149
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_782
timestamp 1644511149
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_783
timestamp 1644511149
transform 1 0 24288 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_784
timestamp 1644511149
transform 1 0 29440 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_785
timestamp 1644511149
transform 1 0 34592 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_786
timestamp 1644511149
transform 1 0 39744 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_787
timestamp 1644511149
transform 1 0 44896 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_788
timestamp 1644511149
transform 1 0 50048 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_789
timestamp 1644511149
transform 1 0 55200 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_790
timestamp 1644511149
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_791
timestamp 1644511149
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_792
timestamp 1644511149
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_793
timestamp 1644511149
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_794
timestamp 1644511149
transform 1 0 26864 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_795
timestamp 1644511149
transform 1 0 32016 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_796
timestamp 1644511149
transform 1 0 37168 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_797
timestamp 1644511149
transform 1 0 42320 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_798
timestamp 1644511149
transform 1 0 47472 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_799
timestamp 1644511149
transform 1 0 52624 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_800
timestamp 1644511149
transform 1 0 57776 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_801
timestamp 1644511149
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_802
timestamp 1644511149
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_803
timestamp 1644511149
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_804
timestamp 1644511149
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_805
timestamp 1644511149
transform 1 0 24288 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_806
timestamp 1644511149
transform 1 0 29440 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_807
timestamp 1644511149
transform 1 0 34592 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_808
timestamp 1644511149
transform 1 0 39744 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_809
timestamp 1644511149
transform 1 0 44896 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_810
timestamp 1644511149
transform 1 0 50048 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_811
timestamp 1644511149
transform 1 0 55200 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_812
timestamp 1644511149
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_813
timestamp 1644511149
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_814
timestamp 1644511149
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_815
timestamp 1644511149
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_816
timestamp 1644511149
transform 1 0 26864 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_817
timestamp 1644511149
transform 1 0 32016 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_818
timestamp 1644511149
transform 1 0 37168 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_819
timestamp 1644511149
transform 1 0 42320 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_820
timestamp 1644511149
transform 1 0 47472 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_821
timestamp 1644511149
transform 1 0 52624 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_822
timestamp 1644511149
transform 1 0 57776 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_823
timestamp 1644511149
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_824
timestamp 1644511149
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_825
timestamp 1644511149
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_826
timestamp 1644511149
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_827
timestamp 1644511149
transform 1 0 24288 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_828
timestamp 1644511149
transform 1 0 29440 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_829
timestamp 1644511149
transform 1 0 34592 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_830
timestamp 1644511149
transform 1 0 39744 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_831
timestamp 1644511149
transform 1 0 44896 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_832
timestamp 1644511149
transform 1 0 50048 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_833
timestamp 1644511149
transform 1 0 55200 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_834
timestamp 1644511149
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_835
timestamp 1644511149
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_836
timestamp 1644511149
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_837
timestamp 1644511149
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_838
timestamp 1644511149
transform 1 0 26864 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_839
timestamp 1644511149
transform 1 0 32016 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_840
timestamp 1644511149
transform 1 0 37168 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_841
timestamp 1644511149
transform 1 0 42320 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_842
timestamp 1644511149
transform 1 0 47472 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_843
timestamp 1644511149
transform 1 0 52624 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_844
timestamp 1644511149
transform 1 0 57776 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_845
timestamp 1644511149
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_846
timestamp 1644511149
transform 1 0 6256 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_847
timestamp 1644511149
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_848
timestamp 1644511149
transform 1 0 11408 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_849
timestamp 1644511149
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_850
timestamp 1644511149
transform 1 0 16560 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_851
timestamp 1644511149
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_852
timestamp 1644511149
transform 1 0 21712 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_853
timestamp 1644511149
transform 1 0 24288 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_854
timestamp 1644511149
transform 1 0 26864 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_855
timestamp 1644511149
transform 1 0 29440 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_856
timestamp 1644511149
transform 1 0 32016 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_857
timestamp 1644511149
transform 1 0 34592 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_858
timestamp 1644511149
transform 1 0 37168 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_859
timestamp 1644511149
transform 1 0 39744 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_860
timestamp 1644511149
transform 1 0 42320 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_861
timestamp 1644511149
transform 1 0 44896 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_862
timestamp 1644511149
transform 1 0 47472 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_863
timestamp 1644511149
transform 1 0 50048 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_864
timestamp 1644511149
transform 1 0 52624 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_865
timestamp 1644511149
transform 1 0 55200 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_866
timestamp 1644511149
transform 1 0 57776 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__or2_1  _1475_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 53728 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1476_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 52716 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o211ai_4  _1477_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 54280 0 1 10880
box -38 -48 1602 592
use sky130_fd_sc_hd__xnor2_4  _1478_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 5980 0 1 13056
box -38 -48 2062 592
use sky130_fd_sc_hd__xor2_1  _1479_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 7360 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1480_
timestamp 1644511149
transform 1 0 8096 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1481_
timestamp 1644511149
transform -1 0 7728 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1482_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 8372 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1483_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 7728 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_2  _1484_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6348 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1485_
timestamp 1644511149
transform 1 0 9108 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o31ai_4  _1486_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 9936 0 -1 13056
box -38 -48 1602 592
use sky130_fd_sc_hd__nor2_1  _1487_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 8188 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1488_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 9108 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1489_
timestamp 1644511149
transform 1 0 10580 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o2bb2a_1  _1490_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 10304 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1491_
timestamp 1644511149
transform -1 0 17112 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1492_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 14352 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1493_
timestamp 1644511149
transform -1 0 17296 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1494_
timestamp 1644511149
transform 1 0 15640 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1495_
timestamp 1644511149
transform 1 0 14444 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1496_
timestamp 1644511149
transform 1 0 12880 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _1497_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 14076 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _1498_
timestamp 1644511149
transform -1 0 13524 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1499_
timestamp 1644511149
transform 1 0 27508 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _1500_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 27324 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1501_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17204 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1502_
timestamp 1644511149
transform 1 0 18492 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1503_
timestamp 1644511149
transform -1 0 20424 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1504_
timestamp 1644511149
transform -1 0 25944 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1505_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20148 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1506_
timestamp 1644511149
transform -1 0 20516 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1507_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19780 0 -1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _1508_
timestamp 1644511149
transform -1 0 10672 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1509_
timestamp 1644511149
transform -1 0 10212 0 1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1510_
timestamp 1644511149
transform -1 0 7268 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1511_
timestamp 1644511149
transform -1 0 8188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _1512_
timestamp 1644511149
transform -1 0 6624 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1513_
timestamp 1644511149
transform -1 0 6992 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1514_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 6072 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1515_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6440 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1516_
timestamp 1644511149
transform -1 0 6808 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1517_
timestamp 1644511149
transform 1 0 6348 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1518_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 5888 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _1519_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 4324 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _1520_
timestamp 1644511149
transform -1 0 3312 0 1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _1521_
timestamp 1644511149
transform -1 0 3404 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1522_
timestamp 1644511149
transform -1 0 2668 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _1523_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6348 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1524_
timestamp 1644511149
transform -1 0 17940 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1525_
timestamp 1644511149
transform -1 0 20332 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1526_
timestamp 1644511149
transform 1 0 16560 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1527_
timestamp 1644511149
transform 1 0 16560 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1528_
timestamp 1644511149
transform -1 0 16192 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _1529_
timestamp 1644511149
transform -1 0 16928 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1530_
timestamp 1644511149
transform 1 0 16652 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1531_
timestamp 1644511149
transform 1 0 17572 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1532_
timestamp 1644511149
transform -1 0 23552 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__mux2_2  _1533_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 23920 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_4  _1534_
timestamp 1644511149
transform 1 0 23644 0 -1 7616
box -38 -48 2062 592
use sky130_fd_sc_hd__nor2_1  _1535_
timestamp 1644511149
transform -1 0 21896 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1536_
timestamp 1644511149
transform -1 0 25576 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1537_
timestamp 1644511149
transform 1 0 22356 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1538_
timestamp 1644511149
transform 1 0 22172 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_4  _1539_
timestamp 1644511149
transform 1 0 24472 0 1 6528
box -38 -48 2062 592
use sky130_fd_sc_hd__nor2_1  _1540_
timestamp 1644511149
transform -1 0 12972 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1541_
timestamp 1644511149
transform 1 0 12696 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1542_
timestamp 1644511149
transform 1 0 14076 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1543_
timestamp 1644511149
transform 1 0 13432 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1544_
timestamp 1644511149
transform -1 0 13708 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _1545_
timestamp 1644511149
transform -1 0 10764 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1546_
timestamp 1644511149
transform -1 0 7452 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1547_
timestamp 1644511149
transform -1 0 6992 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1548_
timestamp 1644511149
transform -1 0 4048 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1549_
timestamp 1644511149
transform -1 0 4324 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _1550_
timestamp 1644511149
transform 1 0 3772 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1551_
timestamp 1644511149
transform -1 0 4508 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1552_
timestamp 1644511149
transform 1 0 3772 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _1553_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 3220 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1554_
timestamp 1644511149
transform -1 0 7360 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1555_
timestamp 1644511149
transform 1 0 5152 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _1556_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 6532 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_4  _1557_
timestamp 1644511149
transform -1 0 4232 0 -1 13056
box -38 -48 2062 592
use sky130_fd_sc_hd__xnor2_4  _1558_
timestamp 1644511149
transform 1 0 1932 0 -1 23936
box -38 -48 2062 592
use sky130_fd_sc_hd__and2b_1  _1559_
timestamp 1644511149
transform -1 0 4324 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1560_
timestamp 1644511149
transform -1 0 3680 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_4  _1561_
timestamp 1644511149
transform 1 0 2668 0 -1 22848
box -38 -48 2062 592
use sky130_fd_sc_hd__nor2_1  _1562_
timestamp 1644511149
transform 1 0 3864 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1563_
timestamp 1644511149
transform 1 0 3772 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__a211o_1  _1564_
timestamp 1644511149
transform 1 0 2852 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1565_
timestamp 1644511149
transform -1 0 21252 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1566_
timestamp 1644511149
transform -1 0 20608 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1567_
timestamp 1644511149
transform -1 0 24564 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1568_
timestamp 1644511149
transform -1 0 23276 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1569_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17848 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1570_
timestamp 1644511149
transform -1 0 19596 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1571_
timestamp 1644511149
transform -1 0 23184 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1572_
timestamp 1644511149
transform -1 0 23092 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1573_
timestamp 1644511149
transform -1 0 23552 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1574_
timestamp 1644511149
transform 1 0 24380 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1575_
timestamp 1644511149
transform 1 0 24380 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1576_
timestamp 1644511149
transform 1 0 35972 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1577_
timestamp 1644511149
transform 1 0 33856 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1578_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 35052 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1579_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28152 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1580_
timestamp 1644511149
transform 1 0 28428 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1581_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29624 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1582_
timestamp 1644511149
transform 1 0 30452 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1583_
timestamp 1644511149
transform -1 0 31648 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1584_
timestamp 1644511149
transform 1 0 31096 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1585_
timestamp 1644511149
transform 1 0 31188 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1586_
timestamp 1644511149
transform -1 0 27968 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1587_
timestamp 1644511149
transform -1 0 27600 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1588_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19596 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1589_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19688 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1590_
timestamp 1644511149
transform -1 0 19872 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1591_
timestamp 1644511149
transform -1 0 17756 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1592_
timestamp 1644511149
transform -1 0 17204 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1593_
timestamp 1644511149
transform -1 0 16376 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1594_
timestamp 1644511149
transform -1 0 8372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _1595_
timestamp 1644511149
transform 1 0 6624 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1596_
timestamp 1644511149
transform -1 0 5428 0 1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_1  _1597_
timestamp 1644511149
transform 1 0 2668 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1598_
timestamp 1644511149
transform 1 0 4416 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1599_
timestamp 1644511149
transform 1 0 2852 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _1600_
timestamp 1644511149
transform -1 0 3680 0 -1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _1601_
timestamp 1644511149
transform 1 0 2208 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1602_
timestamp 1644511149
transform 1 0 4784 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1603_
timestamp 1644511149
transform 1 0 2668 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1604_
timestamp 1644511149
transform -1 0 2760 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1605_
timestamp 1644511149
transform 1 0 3772 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _1606_
timestamp 1644511149
transform 1 0 2852 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _1607_
timestamp 1644511149
transform -1 0 3312 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _1608_
timestamp 1644511149
transform -1 0 3128 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1609_
timestamp 1644511149
transform -1 0 6900 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1610_
timestamp 1644511149
transform -1 0 35696 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1611_
timestamp 1644511149
transform -1 0 24932 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1612_
timestamp 1644511149
transform 1 0 24932 0 1 8704
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1613_
timestamp 1644511149
transform 1 0 26220 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _1614_
timestamp 1644511149
transform -1 0 27876 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1615_
timestamp 1644511149
transform -1 0 30820 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1616_
timestamp 1644511149
transform 1 0 32016 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1617_
timestamp 1644511149
transform 1 0 31188 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1618_
timestamp 1644511149
transform -1 0 28888 0 -1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _1619_
timestamp 1644511149
transform 1 0 29532 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1620_
timestamp 1644511149
transform 1 0 30544 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_2  _1621_
timestamp 1644511149
transform 1 0 32844 0 -1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _1622_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 36340 0 1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_1  _1623_
timestamp 1644511149
transform -1 0 33672 0 1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_2  _1624_
timestamp 1644511149
transform -1 0 34040 0 -1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _1625_
timestamp 1644511149
transform -1 0 30912 0 1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__a22o_1  _1626_
timestamp 1644511149
transform -1 0 27416 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1627_
timestamp 1644511149
transform -1 0 25484 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1628_
timestamp 1644511149
transform -1 0 23184 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o21a_1  _1629_
timestamp 1644511149
transform 1 0 16652 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _1630_
timestamp 1644511149
transform 1 0 17572 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1631_
timestamp 1644511149
transform -1 0 16284 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1632_
timestamp 1644511149
transform 1 0 6348 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1633_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 7176 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_2  _1634_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6256 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_2  _1635_
timestamp 1644511149
transform -1 0 3312 0 -1 5440
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1636_
timestamp 1644511149
transform -1 0 3220 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_4  _1637_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 4600 0 -1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__xor2_4  _1638_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 4876 0 -1 6528
box -38 -48 2062 592
use sky130_fd_sc_hd__xnor2_4  _1639_
timestamp 1644511149
transform 1 0 2852 0 -1 14144
box -38 -48 2062 592
use sky130_fd_sc_hd__a21o_1  _1640_
timestamp 1644511149
transform -1 0 3772 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_4  _1641_
timestamp 1644511149
transform 1 0 3864 0 1 16320
box -38 -48 2062 592
use sky130_fd_sc_hd__or2_1  _1642_
timestamp 1644511149
transform 1 0 3772 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1643_
timestamp 1644511149
transform -1 0 3220 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1644_
timestamp 1644511149
transform -1 0 4048 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_2  _1645_
timestamp 1644511149
transform 1 0 3588 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1646_
timestamp 1644511149
transform -1 0 4048 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_2  _1647_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 3680 0 -1 5440
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _1648_
timestamp 1644511149
transform 1 0 28244 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a2bb2o_1  _1649_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 25760 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _1650_
timestamp 1644511149
transform 1 0 36064 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1651_
timestamp 1644511149
transform -1 0 36064 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_2  _1652_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 35512 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1653_
timestamp 1644511149
transform 1 0 35696 0 1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1654_
timestamp 1644511149
transform 1 0 36248 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _1655_
timestamp 1644511149
transform 1 0 27140 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _1656_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 28152 0 -1 6528
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _1657_
timestamp 1644511149
transform 1 0 37260 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1658_
timestamp 1644511149
transform -1 0 37260 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1659_
timestamp 1644511149
transform 1 0 37628 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1660_
timestamp 1644511149
transform -1 0 37168 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1661_
timestamp 1644511149
transform -1 0 37904 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1662_
timestamp 1644511149
transform -1 0 37904 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _1663_
timestamp 1644511149
transform 1 0 33028 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__nor2_1  _1664_
timestamp 1644511149
transform 1 0 33488 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1665_
timestamp 1644511149
transform 1 0 33488 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1666_
timestamp 1644511149
transform 1 0 33856 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1667_
timestamp 1644511149
transform -1 0 33028 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1668_
timestamp 1644511149
transform -1 0 32384 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1669_
timestamp 1644511149
transform 1 0 31280 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_1  _1670_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 23736 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1671_
timestamp 1644511149
transform -1 0 24840 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1672_
timestamp 1644511149
transform -1 0 24104 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_2  _1673_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 23920 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1674_
timestamp 1644511149
transform 1 0 16652 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1675_
timestamp 1644511149
transform 1 0 15916 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1676_
timestamp 1644511149
transform -1 0 10120 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _1677_
timestamp 1644511149
transform 1 0 9384 0 -1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _1678_
timestamp 1644511149
transform -1 0 10488 0 -1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _1679_
timestamp 1644511149
transform -1 0 5704 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1680_
timestamp 1644511149
transform -1 0 28428 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _1681_
timestamp 1644511149
transform -1 0 27876 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _1682_
timestamp 1644511149
transform -1 0 31188 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__o21a_1  _1683_
timestamp 1644511149
transform -1 0 40572 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_1  _1684_
timestamp 1644511149
transform 1 0 40940 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1685_
timestamp 1644511149
transform -1 0 40940 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _1686_
timestamp 1644511149
transform 1 0 39376 0 -1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _1687_
timestamp 1644511149
transform -1 0 37904 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1688_
timestamp 1644511149
transform 1 0 40204 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1689_
timestamp 1644511149
transform 1 0 41308 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1690_
timestamp 1644511149
transform -1 0 41676 0 1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1691_
timestamp 1644511149
transform 1 0 40848 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _1692_
timestamp 1644511149
transform 1 0 37076 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1693_
timestamp 1644511149
transform 1 0 40020 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1694_
timestamp 1644511149
transform 1 0 40664 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1695_
timestamp 1644511149
transform -1 0 40388 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1696_
timestamp 1644511149
transform -1 0 36800 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_2  _1697_
timestamp 1644511149
transform 1 0 32844 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1698_
timestamp 1644511149
transform -1 0 33488 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1699_
timestamp 1644511149
transform -1 0 32660 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1700_
timestamp 1644511149
transform -1 0 23828 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1701_
timestamp 1644511149
transform -1 0 24748 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1702_
timestamp 1644511149
transform 1 0 17664 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1703_
timestamp 1644511149
transform -1 0 9568 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a221oi_4  _1704_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 11316 0 1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__xnor2_1  _1705_
timestamp 1644511149
transform -1 0 17296 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1706_
timestamp 1644511149
transform -1 0 14536 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1707_
timestamp 1644511149
transform -1 0 15180 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1708_
timestamp 1644511149
transform -1 0 14352 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1709_
timestamp 1644511149
transform 1 0 10580 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1710_
timestamp 1644511149
transform 1 0 11224 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_1  _1711_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11500 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1712_
timestamp 1644511149
transform 1 0 12880 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _1713_
timestamp 1644511149
transform 1 0 39744 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1714_
timestamp 1644511149
transform 1 0 44988 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _1715_
timestamp 1644511149
transform -1 0 40204 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _1716_
timestamp 1644511149
transform 1 0 28428 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _1717_
timestamp 1644511149
transform -1 0 32200 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1718_
timestamp 1644511149
transform 1 0 43332 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1719_
timestamp 1644511149
transform 1 0 44988 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__a31o_1  _1720_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 40940 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1721_
timestamp 1644511149
transform -1 0 46828 0 1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1722_
timestamp 1644511149
transform -1 0 46368 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1723_
timestamp 1644511149
transform -1 0 41952 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1724_
timestamp 1644511149
transform -1 0 42872 0 -1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _1725_
timestamp 1644511149
transform -1 0 42504 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _1726_
timestamp 1644511149
transform -1 0 26496 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1727_
timestamp 1644511149
transform -1 0 16928 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1728_
timestamp 1644511149
transform 1 0 17296 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1729_
timestamp 1644511149
transform 1 0 18676 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _1730_
timestamp 1644511149
transform 1 0 19228 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1731_
timestamp 1644511149
transform 1 0 19872 0 1 3264
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _1732_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 20516 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1733_
timestamp 1644511149
transform -1 0 13248 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _1734_
timestamp 1644511149
transform 1 0 12328 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _1735_
timestamp 1644511149
transform 1 0 20700 0 1 2176
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_4  _1736_
timestamp 1644511149
transform 1 0 21160 0 1 3264
box -38 -48 2062 592
use sky130_fd_sc_hd__o31a_2  _1737_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 21160 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1738_
timestamp 1644511149
transform 1 0 25944 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _1739_
timestamp 1644511149
transform -1 0 25484 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1740_
timestamp 1644511149
transform 1 0 26956 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _1741_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 26496 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _1742_
timestamp 1644511149
transform -1 0 46552 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _1743_
timestamp 1644511149
transform -1 0 45356 0 -1 4352
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1744_
timestamp 1644511149
transform 1 0 43516 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_1  _1745_
timestamp 1644511149
transform 1 0 43976 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _1746_
timestamp 1644511149
transform 1 0 43516 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1747_
timestamp 1644511149
transform -1 0 45724 0 -1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _1748_
timestamp 1644511149
transform 1 0 28796 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1749_
timestamp 1644511149
transform -1 0 29072 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1750_
timestamp 1644511149
transform 1 0 27600 0 -1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_4  _1751_
timestamp 1644511149
transform 1 0 29164 0 -1 3264
box -38 -48 2062 592
use sky130_fd_sc_hd__a21oi_1  _1752_
timestamp 1644511149
transform 1 0 28520 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_4  _1753_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28244 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  _1754_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6440 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1755_
timestamp 1644511149
transform -1 0 8096 0 1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _1756_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11040 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1757_
timestamp 1644511149
transform 1 0 27968 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _1758_
timestamp 1644511149
transform 1 0 31280 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1759_
timestamp 1644511149
transform 1 0 21344 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1760_
timestamp 1644511149
transform 1 0 24104 0 -1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _1761_
timestamp 1644511149
transform 1 0 24380 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1762_
timestamp 1644511149
transform -1 0 28152 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1763_
timestamp 1644511149
transform 1 0 19044 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1764_
timestamp 1644511149
transform -1 0 12236 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  _1765_
timestamp 1644511149
transform -1 0 7820 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _1766_
timestamp 1644511149
transform 1 0 10212 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1767_
timestamp 1644511149
transform -1 0 24656 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _1768_
timestamp 1644511149
transform -1 0 5888 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1769_
timestamp 1644511149
transform -1 0 8188 0 -1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _1770_
timestamp 1644511149
transform 1 0 11500 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1771_
timestamp 1644511149
transform 1 0 24656 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _1772_
timestamp 1644511149
transform 1 0 24932 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1773_
timestamp 1644511149
transform 1 0 26772 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1774_
timestamp 1644511149
transform -1 0 26404 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1775_
timestamp 1644511149
transform 1 0 27232 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1776_
timestamp 1644511149
transform 1 0 27876 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1777_
timestamp 1644511149
transform -1 0 28336 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1778_
timestamp 1644511149
transform -1 0 28152 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1779_
timestamp 1644511149
transform -1 0 27876 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _1780_
timestamp 1644511149
transform -1 0 8464 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1781_
timestamp 1644511149
transform -1 0 7820 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1782_
timestamp 1644511149
transform 1 0 6900 0 1 26112
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  _1783_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 17020 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1784_
timestamp 1644511149
transform 1 0 11960 0 1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1785_
timestamp 1644511149
transform 1 0 10028 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1786_
timestamp 1644511149
transform 1 0 9200 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_2  _1787_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 10856 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _1788_
timestamp 1644511149
transform 1 0 3496 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1789_
timestamp 1644511149
transform 1 0 9200 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1790_
timestamp 1644511149
transform 1 0 23460 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _1791_
timestamp 1644511149
transform 1 0 25300 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_1  _1792_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 23920 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1793_
timestamp 1644511149
transform 1 0 19780 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1794_
timestamp 1644511149
transform 1 0 24104 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__o211a_1  _1795_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 25116 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _1796_
timestamp 1644511149
transform -1 0 29072 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1797_
timestamp 1644511149
transform -1 0 27232 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1798_
timestamp 1644511149
transform 1 0 28152 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_1  _1799_
timestamp 1644511149
transform -1 0 28612 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _1800_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28060 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_2  _1801_
timestamp 1644511149
transform 1 0 29072 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1802_
timestamp 1644511149
transform -1 0 43424 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _1803_
timestamp 1644511149
transform -1 0 11592 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1804_
timestamp 1644511149
transform -1 0 11868 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1805_
timestamp 1644511149
transform -1 0 11316 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1806_
timestamp 1644511149
transform 1 0 9936 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1807_
timestamp 1644511149
transform -1 0 10856 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1808_
timestamp 1644511149
transform 1 0 11500 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _1809_
timestamp 1644511149
transform 1 0 9936 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1810_
timestamp 1644511149
transform 1 0 6716 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_4  _1811_
timestamp 1644511149
transform 1 0 16652 0 -1 29376
box -38 -48 2062 592
use sky130_fd_sc_hd__xor2_1  _1812_
timestamp 1644511149
transform 1 0 5428 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1813_
timestamp 1644511149
transform -1 0 7728 0 1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__and3b_1  _1814_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 9292 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and3b_1  _1815_
timestamp 1644511149
transform 1 0 10304 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1816_
timestamp 1644511149
transform 1 0 5060 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nor3b_1  _1817_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 9568 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__nor4_1  _1818_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 10212 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_4  _1819_
timestamp 1644511149
transform 1 0 18308 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _1820_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 10028 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _1821_
timestamp 1644511149
transform 1 0 10580 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1822_
timestamp 1644511149
transform 1 0 10396 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _1823_
timestamp 1644511149
transform 1 0 20700 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1824_
timestamp 1644511149
transform -1 0 23276 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _1825_
timestamp 1644511149
transform 1 0 22632 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1826_
timestamp 1644511149
transform 1 0 16100 0 1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _1827_
timestamp 1644511149
transform -1 0 15732 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _1828_
timestamp 1644511149
transform 1 0 16652 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1829_
timestamp 1644511149
transform 1 0 24380 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1830_
timestamp 1644511149
transform 1 0 26772 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _1831_
timestamp 1644511149
transform 1 0 27508 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _1832_
timestamp 1644511149
transform -1 0 28244 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_2  _1833_
timestamp 1644511149
transform -1 0 27784 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1834_
timestamp 1644511149
transform -1 0 3128 0 -1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__and2_1  _1835_
timestamp 1644511149
transform -1 0 28244 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1836_
timestamp 1644511149
transform 1 0 24196 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1837_
timestamp 1644511149
transform -1 0 9660 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1838_
timestamp 1644511149
transform -1 0 8556 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1839_
timestamp 1644511149
transform -1 0 8280 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1840_
timestamp 1644511149
transform -1 0 6532 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _1841_
timestamp 1644511149
transform -1 0 7452 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _1842_
timestamp 1644511149
transform 1 0 7268 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_2  _1843_
timestamp 1644511149
transform 1 0 9568 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _1844_
timestamp 1644511149
transform 1 0 16560 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_4  _1845_
timestamp 1644511149
transform 1 0 16652 0 -1 28288
box -38 -48 2062 592
use sky130_fd_sc_hd__nor2_1  _1846_
timestamp 1644511149
transform -1 0 9200 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1847_
timestamp 1644511149
transform -1 0 13984 0 -1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__a2bb2o_1  _1848_
timestamp 1644511149
transform 1 0 14352 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1849_
timestamp 1644511149
transform 1 0 3772 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1850_
timestamp 1644511149
transform -1 0 7728 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1851_
timestamp 1644511149
transform 1 0 12052 0 -1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__and3_2  _1852_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6900 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _1853_
timestamp 1644511149
transform 1 0 12420 0 1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _1854_
timestamp 1644511149
transform 1 0 12880 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1855_
timestamp 1644511149
transform 1 0 12972 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _1856_
timestamp 1644511149
transform 1 0 13340 0 -1 31552
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1857_
timestamp 1644511149
transform 1 0 13248 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1858_
timestamp 1644511149
transform 1 0 15180 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nor3_1  _1859_
timestamp 1644511149
transform -1 0 10212 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _1860_
timestamp 1644511149
transform -1 0 15272 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _1861_
timestamp 1644511149
transform 1 0 14996 0 -1 34816
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _1862_
timestamp 1644511149
transform 1 0 24656 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1863_
timestamp 1644511149
transform 1 0 26220 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _1864_
timestamp 1644511149
transform 1 0 26772 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _1865_
timestamp 1644511149
transform -1 0 28704 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_4  _1866_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 27692 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  _1867_
timestamp 1644511149
transform 1 0 2208 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1868_
timestamp 1644511149
transform 1 0 24656 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1869_
timestamp 1644511149
transform 1 0 16652 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1870_
timestamp 1644511149
transform 1 0 15640 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__buf_4  _1871_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 37260 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1872_
timestamp 1644511149
transform -1 0 8464 0 1 33728
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1873_
timestamp 1644511149
transform -1 0 6992 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1874_
timestamp 1644511149
transform -1 0 7728 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1875_
timestamp 1644511149
transform 1 0 5612 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_2  _1876_
timestamp 1644511149
transform -1 0 7084 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1877_
timestamp 1644511149
transform -1 0 18676 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1878_
timestamp 1644511149
transform 1 0 9384 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _1879_
timestamp 1644511149
transform 1 0 11500 0 1 32640
box -38 -48 1234 592
use sky130_fd_sc_hd__o21a_2  _1880_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16192 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_4  _1881_
timestamp 1644511149
transform 1 0 12788 0 -1 32640
box -38 -48 2062 592
use sky130_fd_sc_hd__and2_1  _1882_
timestamp 1644511149
transform 1 0 14996 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _1883_
timestamp 1644511149
transform 1 0 14444 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _1884_
timestamp 1644511149
transform -1 0 16284 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o31ai_2  _1885_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 15272 0 -1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__or4_1  _1886_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 16652 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_2  _1887_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 18032 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1888_
timestamp 1644511149
transform -1 0 18492 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _1889_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 18216 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1890_
timestamp 1644511149
transform -1 0 18768 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _1891_
timestamp 1644511149
transform 1 0 5244 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _1892_
timestamp 1644511149
transform 1 0 6808 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1893_
timestamp 1644511149
transform 1 0 18492 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _1894_
timestamp 1644511149
transform -1 0 19872 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _1895_
timestamp 1644511149
transform -1 0 18768 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _1896_
timestamp 1644511149
transform 1 0 19228 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1897_
timestamp 1644511149
transform 1 0 18308 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1898_
timestamp 1644511149
transform 1 0 18124 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__or3_2  _1899_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 19596 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_2  _1900_
timestamp 1644511149
transform 1 0 18584 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_2  _1901_
timestamp 1644511149
transform 1 0 25116 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _1902_
timestamp 1644511149
transform -1 0 25484 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1903_
timestamp 1644511149
transform 1 0 27692 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _1904_
timestamp 1644511149
transform -1 0 27876 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1905_
timestamp 1644511149
transform -1 0 27600 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _1906_
timestamp 1644511149
transform 1 0 28520 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _1907_
timestamp 1644511149
transform 1 0 27968 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _1908_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 28520 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _1909_
timestamp 1644511149
transform -1 0 51612 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand3_1  _1910_
timestamp 1644511149
transform 1 0 27692 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1911_
timestamp 1644511149
transform -1 0 9844 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1912_
timestamp 1644511149
transform 1 0 11224 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1913_
timestamp 1644511149
transform 1 0 8648 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _1914_
timestamp 1644511149
transform 1 0 9844 0 1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _1915_
timestamp 1644511149
transform 1 0 9936 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1916_
timestamp 1644511149
transform -1 0 9752 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1917_
timestamp 1644511149
transform 1 0 9200 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_2  _1918_
timestamp 1644511149
transform -1 0 10856 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _1919_
timestamp 1644511149
transform 1 0 19228 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _1920_
timestamp 1644511149
transform -1 0 16100 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _1921_
timestamp 1644511149
transform -1 0 12236 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_2  _1922_
timestamp 1644511149
transform -1 0 12788 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _1923_
timestamp 1644511149
transform 1 0 10856 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _1924_
timestamp 1644511149
transform 1 0 11316 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_2  _1925_
timestamp 1644511149
transform 1 0 11684 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_4  _1926_
timestamp 1644511149
transform 1 0 12236 0 -1 34816
box -38 -48 2062 592
use sky130_fd_sc_hd__a22o_1  _1927_
timestamp 1644511149
transform 1 0 10396 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _1928_
timestamp 1644511149
transform 1 0 13340 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _1929_
timestamp 1644511149
transform 1 0 19688 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_2  _1930_
timestamp 1644511149
transform 1 0 20700 0 1 31552
box -38 -48 1234 592
use sky130_fd_sc_hd__inv_2  _1931_
timestamp 1644511149
transform 1 0 33856 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  _1932_
timestamp 1644511149
transform 1 0 34776 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_2  _1933_
timestamp 1644511149
transform -1 0 22448 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _1934_
timestamp 1644511149
transform 1 0 21712 0 1 32640
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_4  _1935_
timestamp 1644511149
transform 1 0 34684 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1936_
timestamp 1644511149
transform -1 0 24564 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__xor2_2  _1937_
timestamp 1644511149
transform -1 0 20424 0 1 28288
box -38 -48 1234 592
use sky130_fd_sc_hd__and2b_1  _1938_
timestamp 1644511149
transform -1 0 13616 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _1939_
timestamp 1644511149
transform 1 0 17020 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1940_
timestamp 1644511149
transform 1 0 24748 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _1941_
timestamp 1644511149
transform 1 0 5888 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _1942_
timestamp 1644511149
transform 1 0 7544 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1943_
timestamp 1644511149
transform -1 0 16928 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1944_
timestamp 1644511149
transform 1 0 25668 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _1945_
timestamp 1644511149
transform 1 0 19596 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1946_
timestamp 1644511149
transform -1 0 23920 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _1947_
timestamp 1644511149
transform 1 0 24472 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_2  _1948_
timestamp 1644511149
transform -1 0 26496 0 -1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _1949_
timestamp 1644511149
transform -1 0 23736 0 1 33728
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _1950_
timestamp 1644511149
transform 1 0 20056 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _1951_
timestamp 1644511149
transform -1 0 21896 0 1 34816
box -38 -48 1234 592
use sky130_fd_sc_hd__o21bai_1  _1952_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 19780 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _1953_
timestamp 1644511149
transform 1 0 19688 0 -1 36992
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_1  _1954_
timestamp 1644511149
transform 1 0 28520 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _1955_
timestamp 1644511149
transform -1 0 29716 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _1956_
timestamp 1644511149
transform -1 0 28704 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1957_
timestamp 1644511149
transform 1 0 28244 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1958_
timestamp 1644511149
transform -1 0 28704 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _1959_
timestamp 1644511149
transform -1 0 26496 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _1960_
timestamp 1644511149
transform -1 0 22816 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _1961_
timestamp 1644511149
transform 1 0 20700 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _1962_
timestamp 1644511149
transform 1 0 23000 0 -1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1963_
timestamp 1644511149
transform -1 0 23920 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_2  _1964_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22264 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _1965_
timestamp 1644511149
transform 1 0 10212 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1966_
timestamp 1644511149
transform 1 0 2024 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1967_
timestamp 1644511149
transform 1 0 7912 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _1968_
timestamp 1644511149
transform 1 0 14076 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1969_
timestamp 1644511149
transform 1 0 14996 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _1970_
timestamp 1644511149
transform -1 0 16652 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_2  _1971_
timestamp 1644511149
transform -1 0 17388 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _1972_
timestamp 1644511149
transform 1 0 10580 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__a311o_4  _1973_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 11500 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__and2_1  _1974_
timestamp 1644511149
transform -1 0 8096 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _1975_
timestamp 1644511149
transform 1 0 8372 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _1976_
timestamp 1644511149
transform -1 0 6992 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_4  _1977_
timestamp 1644511149
transform 1 0 6440 0 1 31552
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_2  _1978_
timestamp 1644511149
transform 1 0 14260 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1979_
timestamp 1644511149
transform 1 0 14720 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__a22oi_1  _1980_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 14076 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _1981_
timestamp 1644511149
transform 1 0 13064 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o211a_1  _1982_
timestamp 1644511149
transform -1 0 14812 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_4  _1983_
timestamp 1644511149
transform 1 0 14076 0 1 30464
box -38 -48 2062 592
use sky130_fd_sc_hd__xor2_2  _1984_
timestamp 1644511149
transform 1 0 29532 0 1 31552
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _1985_
timestamp 1644511149
transform 1 0 30176 0 1 32640
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_2  _1986_
timestamp 1644511149
transform 1 0 18860 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _1987_
timestamp 1644511149
transform 1 0 6992 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _1988_
timestamp 1644511149
transform 1 0 13432 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _1989_
timestamp 1644511149
transform 1 0 17848 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _1990_
timestamp 1644511149
transform 1 0 22908 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _1991_
timestamp 1644511149
transform -1 0 24196 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _1992_
timestamp 1644511149
transform 1 0 24564 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_2  _1993_
timestamp 1644511149
transform 1 0 30084 0 -1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _1994_
timestamp 1644511149
transform 1 0 31096 0 1 33728
box -38 -48 1234 592
use sky130_fd_sc_hd__and2b_1  _1995_
timestamp 1644511149
transform 1 0 21988 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_2  _1996_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 22724 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_4  _1997_
timestamp 1644511149
transform 1 0 32108 0 -1 34816
box -38 -48 2062 592
use sky130_fd_sc_hd__a21o_1  _1998_
timestamp 1644511149
transform -1 0 21804 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _1999_
timestamp 1644511149
transform 1 0 22264 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _2000_
timestamp 1644511149
transform 1 0 23828 0 -1 36992
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _2001_
timestamp 1644511149
transform 1 0 26956 0 -1 36992
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_1  _2002_
timestamp 1644511149
transform -1 0 42872 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2003_
timestamp 1644511149
transform 1 0 43516 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_2  _2004_
timestamp 1644511149
transform 1 0 42504 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_2  _2005_
timestamp 1644511149
transform -1 0 30176 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_4  _2006_
timestamp 1644511149
transform 1 0 42504 0 1 35904
box -38 -48 2062 592
use sky130_fd_sc_hd__or3_1  _2007_
timestamp 1644511149
transform 1 0 24380 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _2008_
timestamp 1644511149
transform 1 0 25668 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _2009_
timestamp 1644511149
transform 1 0 22172 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2010_
timestamp 1644511149
transform 1 0 30636 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _2011_
timestamp 1644511149
transform 1 0 29624 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__clkinv_2  _2012_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 29808 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _2013_
timestamp 1644511149
transform 1 0 4140 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2014_
timestamp 1644511149
transform 1 0 6348 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _2015_
timestamp 1644511149
transform 1 0 7544 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _2016_
timestamp 1644511149
transform 1 0 8004 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_2  _2017_
timestamp 1644511149
transform -1 0 7636 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _2018_
timestamp 1644511149
transform 1 0 30820 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _2019_
timestamp 1644511149
transform 1 0 32200 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _2020_
timestamp 1644511149
transform -1 0 16008 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _2021_
timestamp 1644511149
transform 1 0 7360 0 -1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_2  _2022_
timestamp 1644511149
transform 1 0 8096 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_2  _2023_
timestamp 1644511149
transform 1 0 7084 0 1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_4  _2024_
timestamp 1644511149
transform 1 0 7084 0 -1 32640
box -38 -48 2062 592
use sky130_fd_sc_hd__clkbuf_2  _2025_
timestamp 1644511149
transform -1 0 14812 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _2026_
timestamp 1644511149
transform 1 0 13248 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_2  _2027_
timestamp 1644511149
transform 1 0 14444 0 -1 27200
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_2  _2028_
timestamp 1644511149
transform 1 0 30728 0 1 29376
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _2029_
timestamp 1644511149
transform 1 0 32568 0 -1 30464
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _2030_
timestamp 1644511149
transform 1 0 34684 0 1 31552
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_4  _2031_
timestamp 1644511149
transform 1 0 30636 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _2032_
timestamp 1644511149
transform 1 0 21252 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2033_
timestamp 1644511149
transform 1 0 22448 0 -1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _2034_
timestamp 1644511149
transform 1 0 23644 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _2035_
timestamp 1644511149
transform 1 0 30176 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2036_
timestamp 1644511149
transform 1 0 13248 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _2037_
timestamp 1644511149
transform 1 0 16652 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_2  _2038_
timestamp 1644511149
transform 1 0 17848 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _2039_
timestamp 1644511149
transform 1 0 30360 0 1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _2040_
timestamp 1644511149
transform 1 0 32108 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _2041_
timestamp 1644511149
transform 1 0 32108 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _2042_
timestamp 1644511149
transform 1 0 33764 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _2043_
timestamp 1644511149
transform 1 0 34684 0 1 32640
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _2044_
timestamp 1644511149
transform -1 0 30728 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _2045_
timestamp 1644511149
transform -1 0 31464 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_2  _2046_
timestamp 1644511149
transform -1 0 36248 0 1 33728
box -38 -48 1234 592
use sky130_fd_sc_hd__or2b_1  _2047_
timestamp 1644511149
transform 1 0 32660 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _2048_
timestamp 1644511149
transform 1 0 23460 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2049_
timestamp 1644511149
transform -1 0 36064 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _2050_
timestamp 1644511149
transform -1 0 35328 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _2051_
timestamp 1644511149
transform 1 0 32108 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2052_
timestamp 1644511149
transform 1 0 32200 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2053_
timestamp 1644511149
transform 1 0 34684 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2054_
timestamp 1644511149
transform 1 0 34776 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_2  _2055_
timestamp 1644511149
transform 1 0 35512 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_2  _2056_
timestamp 1644511149
transform 1 0 41308 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_4  _2057_
timestamp 1644511149
transform -1 0 37536 0 1 35904
box -38 -48 2062 592
use sky130_fd_sc_hd__or2b_1  _2058_
timestamp 1644511149
transform 1 0 31280 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _2059_
timestamp 1644511149
transform -1 0 33672 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_2  _2060_
timestamp 1644511149
transform 1 0 32292 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2061_
timestamp 1644511149
transform -1 0 37444 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _2062_
timestamp 1644511149
transform 1 0 17020 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _2063_
timestamp 1644511149
transform -1 0 5244 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _2064_
timestamp 1644511149
transform 1 0 12972 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2065_
timestamp 1644511149
transform 1 0 23460 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _2066_
timestamp 1644511149
transform -1 0 24196 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _2067_
timestamp 1644511149
transform -1 0 25024 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2068_
timestamp 1644511149
transform 1 0 2760 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2069_
timestamp 1644511149
transform -1 0 3312 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _2070_
timestamp 1644511149
transform 1 0 5060 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _2071_
timestamp 1644511149
transform 1 0 8924 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__a31o_4  _2072_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 6900 0 -1 31552
box -38 -48 1326 592
use sky130_fd_sc_hd__xor2_4  _2073_
timestamp 1644511149
transform 1 0 6992 0 -1 21760
box -38 -48 2062 592
use sky130_fd_sc_hd__a22o_1  _2074_
timestamp 1644511149
transform 1 0 12972 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_2  _2075_
timestamp 1644511149
transform 1 0 14076 0 1 25024
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _2076_
timestamp 1644511149
transform 1 0 31188 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _2077_
timestamp 1644511149
transform 1 0 33580 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _2078_
timestamp 1644511149
transform 1 0 31188 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _2079_
timestamp 1644511149
transform 1 0 32292 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _2080_
timestamp 1644511149
transform 1 0 34960 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _2081_
timestamp 1644511149
transform 1 0 18860 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _2082_
timestamp 1644511149
transform 1 0 17756 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _2083_
timestamp 1644511149
transform 1 0 19780 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_2  _2084_
timestamp 1644511149
transform 1 0 20792 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _2085_
timestamp 1644511149
transform 1 0 33856 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _2086_
timestamp 1644511149
transform 1 0 20056 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _2087_
timestamp 1644511149
transform -1 0 21528 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _2088_
timestamp 1644511149
transform 1 0 20976 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _2089_
timestamp 1644511149
transform 1 0 22264 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _2090_
timestamp 1644511149
transform -1 0 23736 0 1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _2091_
timestamp 1644511149
transform -1 0 23092 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _2092_
timestamp 1644511149
transform 1 0 22724 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2093_
timestamp 1644511149
transform 1 0 23552 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _2094_
timestamp 1644511149
transform 1 0 24380 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _2095_
timestamp 1644511149
transform 1 0 34684 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2096_
timestamp 1644511149
transform 1 0 36432 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2097_
timestamp 1644511149
transform -1 0 37536 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2098_
timestamp 1644511149
transform -1 0 37444 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _2099_
timestamp 1644511149
transform 1 0 37260 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2100_
timestamp 1644511149
transform -1 0 34224 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _2101_
timestamp 1644511149
transform -1 0 35052 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _2102_
timestamp 1644511149
transform -1 0 38456 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2103_
timestamp 1644511149
transform 1 0 37996 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _2104_
timestamp 1644511149
transform 1 0 38456 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _2105_
timestamp 1644511149
transform 1 0 38916 0 -1 32640
box -38 -48 1234 592
use sky130_fd_sc_hd__or2b_1  _2106_
timestamp 1644511149
transform 1 0 35696 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__or2_1  _2107_
timestamp 1644511149
transform 1 0 34960 0 -1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2108_
timestamp 1644511149
transform -1 0 40204 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _2109_
timestamp 1644511149
transform -1 0 40296 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2110_
timestamp 1644511149
transform 1 0 37628 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2111_
timestamp 1644511149
transform 1 0 37996 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2112_
timestamp 1644511149
transform -1 0 39284 0 1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2113_
timestamp 1644511149
transform 1 0 40296 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_2  _2114_
timestamp 1644511149
transform 1 0 39284 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_2  _2115_
timestamp 1644511149
transform -1 0 36248 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_4  _2116_
timestamp 1644511149
transform 1 0 39836 0 1 35904
box -38 -48 2062 592
use sky130_fd_sc_hd__and2b_1  _2117_
timestamp 1644511149
transform 1 0 37904 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _2118_
timestamp 1644511149
transform 1 0 37444 0 1 34816
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_2  _2119_
timestamp 1644511149
transform -1 0 39284 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2120_
timestamp 1644511149
transform -1 0 41032 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _2121_
timestamp 1644511149
transform 1 0 35972 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__o31ai_2  _2122_
timestamp 1644511149
transform -1 0 38180 0 -1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__or2b_1  _2123_
timestamp 1644511149
transform 1 0 34684 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _2124_
timestamp 1644511149
transform -1 0 25760 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2125_
timestamp 1644511149
transform 1 0 24380 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_4  _2126_
timestamp 1644511149
transform 1 0 2300 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _2127_
timestamp 1644511149
transform 1 0 10672 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2128_
timestamp 1644511149
transform 1 0 24196 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _2129_
timestamp 1644511149
transform -1 0 26404 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _2130_
timestamp 1644511149
transform -1 0 26036 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _2131_
timestamp 1644511149
transform -1 0 25668 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _2132_
timestamp 1644511149
transform 1 0 34684 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _2133_
timestamp 1644511149
transform 1 0 2300 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2134_
timestamp 1644511149
transform 1 0 2116 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _2135_
timestamp 1644511149
transform 1 0 2484 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _2136_
timestamp 1644511149
transform 1 0 4140 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_4  _2137_
timestamp 1644511149
transform 1 0 3864 0 -1 21760
box -38 -48 2062 592
use sky130_fd_sc_hd__clkbuf_2  _2138_
timestamp 1644511149
transform -1 0 13616 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _2139_
timestamp 1644511149
transform 1 0 12788 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_2  _2140_
timestamp 1644511149
transform 1 0 13800 0 -1 22848
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _2141_
timestamp 1644511149
transform 1 0 37260 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _2142_
timestamp 1644511149
transform 1 0 37076 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _2143_
timestamp 1644511149
transform 1 0 37996 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _2144_
timestamp 1644511149
transform 1 0 22356 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _2145_
timestamp 1644511149
transform -1 0 22448 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _2146_
timestamp 1644511149
transform 1 0 21528 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _2147_
timestamp 1644511149
transform -1 0 23920 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_1  _2148_
timestamp 1644511149
transform 1 0 24012 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _2149_
timestamp 1644511149
transform 1 0 34776 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2150_
timestamp 1644511149
transform 1 0 20700 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2151_
timestamp 1644511149
transform 1 0 16284 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _2152_
timestamp 1644511149
transform -1 0 21068 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2153_
timestamp 1644511149
transform 1 0 32476 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2154_
timestamp 1644511149
transform 1 0 36248 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2155_
timestamp 1644511149
transform 1 0 36340 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2156_
timestamp 1644511149
transform 1 0 37536 0 1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _2157_
timestamp 1644511149
transform 1 0 38640 0 1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2158_
timestamp 1644511149
transform 1 0 39560 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _2159_
timestamp 1644511149
transform 1 0 40572 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _2160_
timestamp 1644511149
transform 1 0 38640 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _2161_
timestamp 1644511149
transform 1 0 41124 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2162_
timestamp 1644511149
transform 1 0 41676 0 1 33728
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2163_
timestamp 1644511149
transform -1 0 43240 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _2164_
timestamp 1644511149
transform 1 0 43148 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _2165_
timestamp 1644511149
transform 1 0 44988 0 -1 35904
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_4  _2166_
timestamp 1644511149
transform -1 0 47840 0 1 35904
box -38 -48 2062 592
use sky130_fd_sc_hd__a21o_2  _2167_
timestamp 1644511149
transform -1 0 38916 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_4  _2168_
timestamp 1644511149
transform -1 0 47104 0 -1 36992
box -38 -48 2062 592
use sky130_fd_sc_hd__nand2_1  _2169_
timestamp 1644511149
transform 1 0 42412 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2170_
timestamp 1644511149
transform 1 0 41676 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2171_
timestamp 1644511149
transform 1 0 38548 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2172_
timestamp 1644511149
transform 1 0 39100 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _2173_
timestamp 1644511149
transform 1 0 38088 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _2174_
timestamp 1644511149
transform 1 0 2208 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2175_
timestamp 1644511149
transform 1 0 9108 0 1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _2176_
timestamp 1644511149
transform 1 0 9936 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _2177_
timestamp 1644511149
transform 1 0 9476 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_2  _2178_
timestamp 1644511149
transform -1 0 10672 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _2179_
timestamp 1644511149
transform 1 0 33488 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_2  _2180_
timestamp 1644511149
transform 1 0 7268 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__or4b_2  _2181_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 4876 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__and2_1  _2182_
timestamp 1644511149
transform -1 0 5796 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2183_
timestamp 1644511149
transform 1 0 2852 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _2184_
timestamp 1644511149
transform 1 0 4416 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_1  _2185_
timestamp 1644511149
transform -1 0 8188 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2186_
timestamp 1644511149
transform 1 0 8004 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__or3_4  _2187_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 9660 0 -1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__a22o_1  _2188_
timestamp 1644511149
transform 1 0 12972 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _2189_
timestamp 1644511149
transform -1 0 14720 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _2190_
timestamp 1644511149
transform -1 0 35788 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _2191_
timestamp 1644511149
transform -1 0 35052 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _2192_
timestamp 1644511149
transform 1 0 34776 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _2193_
timestamp 1644511149
transform 1 0 34592 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _2194_
timestamp 1644511149
transform 1 0 37720 0 -1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _2195_
timestamp 1644511149
transform 1 0 39008 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _2196_
timestamp 1644511149
transform 1 0 19964 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _2197_
timestamp 1644511149
transform 1 0 16652 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_2  _2198_
timestamp 1644511149
transform 1 0 17296 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _2199_
timestamp 1644511149
transform 1 0 34684 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__and2_2  _2200_
timestamp 1644511149
transform -1 0 22448 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _2201_
timestamp 1644511149
transform 1 0 17020 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_2  _2202_
timestamp 1644511149
transform 1 0 19228 0 1 26112
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_2  _2203_
timestamp 1644511149
transform 1 0 30452 0 1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_1  _2204_
timestamp 1644511149
transform 1 0 37260 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _2205_
timestamp 1644511149
transform 1 0 33212 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _2206_
timestamp 1644511149
transform 1 0 10856 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _2207_
timestamp 1644511149
transform 1 0 16928 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _2208_
timestamp 1644511149
transform 1 0 27416 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _2209_
timestamp 1644511149
transform 1 0 36708 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _2210_
timestamp 1644511149
transform 1 0 38272 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _2211_
timestamp 1644511149
transform 1 0 37628 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _2212_
timestamp 1644511149
transform 1 0 38364 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2213_
timestamp 1644511149
transform 1 0 40940 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _2214_
timestamp 1644511149
transform -1 0 40572 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _2215_
timestamp 1644511149
transform -1 0 41676 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__o211ai_1  _2216_
timestamp 1644511149
transform -1 0 41676 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__nand3b_1  _2217_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 42412 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__a21bo_1  _2218_
timestamp 1644511149
transform 1 0 41860 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _2219_
timestamp 1644511149
transform -1 0 41124 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2220_
timestamp 1644511149
transform -1 0 40940 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _2221_
timestamp 1644511149
transform 1 0 42596 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _2222_
timestamp 1644511149
transform 1 0 42412 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _2223_
timestamp 1644511149
transform 1 0 43148 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _2224_
timestamp 1644511149
transform 1 0 43148 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2225_
timestamp 1644511149
transform -1 0 45264 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_2  _2226_
timestamp 1644511149
transform 1 0 45080 0 -1 32640
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _2227_
timestamp 1644511149
transform 1 0 43792 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _2228_
timestamp 1644511149
transform -1 0 43424 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2229_
timestamp 1644511149
transform -1 0 45540 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_4  _2230_
timestamp 1644511149
transform 1 0 45724 0 1 32640
box -38 -48 2062 592
use sky130_fd_sc_hd__xor2_4  _2231_
timestamp 1644511149
transform -1 0 53820 0 1 31552
box -38 -48 2062 592
use sky130_fd_sc_hd__and2_1  _2232_
timestamp 1644511149
transform -1 0 48024 0 -1 36992
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_2  _2233_
timestamp 1644511149
transform -1 0 46828 0 1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_4  _2234_
timestamp 1644511149
transform -1 0 53728 0 1 30464
box -38 -48 2062 592
use sky130_fd_sc_hd__a221oi_2  _2235_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 44620 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__a21bo_1  _2236_
timestamp 1644511149
transform 1 0 40756 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__o21ba_1  _2237_
timestamp 1644511149
transform -1 0 37996 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _2238_
timestamp 1644511149
transform 1 0 8004 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2239_
timestamp 1644511149
transform 1 0 27508 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _2240_
timestamp 1644511149
transform 1 0 28796 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _2241_
timestamp 1644511149
transform 1 0 29624 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _2242_
timestamp 1644511149
transform -1 0 30176 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _2243_
timestamp 1644511149
transform -1 0 14444 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_4  _2244_
timestamp 1644511149
transform 1 0 2300 0 -1 19584
box -38 -48 2062 592
use sky130_fd_sc_hd__a21bo_1  _2245_
timestamp 1644511149
transform -1 0 7176 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a31o_1  _2246_
timestamp 1644511149
transform -1 0 4508 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_4  _2247_
timestamp 1644511149
transform 1 0 3772 0 1 18496
box -38 -48 2062 592
use sky130_fd_sc_hd__a22o_1  _2248_
timestamp 1644511149
transform 1 0 14812 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_2  _2249_
timestamp 1644511149
transform 1 0 15824 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _2250_
timestamp 1644511149
transform 1 0 38732 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _2251_
timestamp 1644511149
transform 1 0 40020 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2252_
timestamp 1644511149
transform 1 0 40848 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2253_
timestamp 1644511149
transform 1 0 12420 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_2  _2254_
timestamp 1644511149
transform 1 0 14076 0 1 23936
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _2255_
timestamp 1644511149
transform 1 0 33764 0 -1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2256_
timestamp 1644511149
transform 1 0 17204 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2257_
timestamp 1644511149
transform 1 0 18032 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _2258_
timestamp 1644511149
transform 1 0 30268 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2259_
timestamp 1644511149
transform 1 0 40020 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2260_
timestamp 1644511149
transform 1 0 40112 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2261_
timestamp 1644511149
transform 1 0 40940 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_2  _2262_
timestamp 1644511149
transform 1 0 11500 0 -1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__and2b_1  _2263_
timestamp 1644511149
transform 1 0 16008 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _2264_
timestamp 1644511149
transform 1 0 10672 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2265_
timestamp 1644511149
transform 1 0 18032 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2266_
timestamp 1644511149
transform 1 0 17572 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2267_
timestamp 1644511149
transform -1 0 18768 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_2  _2268_
timestamp 1644511149
transform 1 0 19044 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _2269_
timestamp 1644511149
transform 1 0 39928 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _2270_
timestamp 1644511149
transform 1 0 41768 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2271_
timestamp 1644511149
transform 1 0 41584 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2272_
timestamp 1644511149
transform 1 0 42596 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_1  _2273_
timestamp 1644511149
transform 1 0 43424 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2274_
timestamp 1644511149
transform 1 0 44068 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _2275_
timestamp 1644511149
transform 1 0 37168 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2276_
timestamp 1644511149
transform 1 0 44988 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2277_
timestamp 1644511149
transform 1 0 42872 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _2278_
timestamp 1644511149
transform -1 0 45356 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2279_
timestamp 1644511149
transform -1 0 44528 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2280_
timestamp 1644511149
transform 1 0 44988 0 1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__o2bb2a_1  _2281_
timestamp 1644511149
transform -1 0 45724 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_2  _2282_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 44896 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _2283_
timestamp 1644511149
transform 1 0 44436 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__o21bai_2  _2284_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 45080 0 1 31552
box -38 -48 866 592
use sky130_fd_sc_hd__o31a_1  _2285_
timestamp 1644511149
transform -1 0 46000 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2286_
timestamp 1644511149
transform -1 0 52164 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2287_
timestamp 1644511149
transform 1 0 50876 0 1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_2  _2288_
timestamp 1644511149
transform 1 0 52716 0 -1 30464
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2289_
timestamp 1644511149
transform -1 0 53176 0 -1 32640
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_2  _2290_
timestamp 1644511149
transform 1 0 51612 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_4  _2291_
timestamp 1644511149
transform -1 0 53544 0 1 29376
box -38 -48 2062 592
use sky130_fd_sc_hd__a21oi_4  _2292_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 51060 0 -1 30464
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _2293_
timestamp 1644511149
transform 1 0 47840 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2294_
timestamp 1644511149
transform -1 0 45724 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2295_
timestamp 1644511149
transform 1 0 41860 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__or2b_1  _2296_
timestamp 1644511149
transform 1 0 43700 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _2297_
timestamp 1644511149
transform -1 0 31924 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _2298_
timestamp 1644511149
transform 1 0 10396 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _2299_
timestamp 1644511149
transform 1 0 28060 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__mux2_1  _2300_
timestamp 1644511149
transform -1 0 27692 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_1  _2301_
timestamp 1644511149
transform 1 0 31004 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _2302_
timestamp 1644511149
transform -1 0 32752 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _2303_
timestamp 1644511149
transform 1 0 26496 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _2304_
timestamp 1644511149
transform 1 0 27232 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a211oi_2  _2305_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 8004 0 -1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__o21a_1  _2306_
timestamp 1644511149
transform -1 0 7636 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_2  _2307_
timestamp 1644511149
transform 1 0 4968 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2308_
timestamp 1644511149
transform 1 0 1840 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2309_
timestamp 1644511149
transform 1 0 5796 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_4  _2310_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 7452 0 -1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__or3_1  _2311_
timestamp 1644511149
transform 1 0 7636 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a32o_1  _2312_
timestamp 1644511149
transform 1 0 13064 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__o21ai_1  _2313_
timestamp 1644511149
transform 1 0 30912 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _2314_
timestamp 1644511149
transform 1 0 30728 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and3_2  _2315_
timestamp 1644511149
transform 1 0 32568 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _2316_
timestamp 1644511149
transform 1 0 31556 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _2317_
timestamp 1644511149
transform 1 0 40296 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__or3b_1  _2318_
timestamp 1644511149
transform 1 0 42504 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__o21bai_1  _2319_
timestamp 1644511149
transform 1 0 42504 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  _2320_
timestamp 1644511149
transform 1 0 23368 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__nor2_1  _2321_
timestamp 1644511149
transform -1 0 20792 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _2322_
timestamp 1644511149
transform 1 0 14904 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _2323_
timestamp 1644511149
transform 1 0 21160 0 1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _2324_
timestamp 1644511149
transform -1 0 22448 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2325_
timestamp 1644511149
transform 1 0 27876 0 -1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2326_
timestamp 1644511149
transform 1 0 17296 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2327_
timestamp 1644511149
transform 1 0 19136 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _2328_
timestamp 1644511149
transform 1 0 26588 0 1 22848
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2329_
timestamp 1644511149
transform 1 0 29532 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2330_
timestamp 1644511149
transform -1 0 29072 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2331_
timestamp 1644511149
transform 1 0 30176 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__and2b_1  _2332_
timestamp 1644511149
transform 1 0 17112 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _2333_
timestamp 1644511149
transform 1 0 17572 0 -1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _2334_
timestamp 1644511149
transform -1 0 19596 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_1  _2335_
timestamp 1644511149
transform -1 0 18768 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__a221o_2  _2336_
timestamp 1644511149
transform 1 0 19228 0 1 20672
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_2  _2337_
timestamp 1644511149
transform 1 0 30452 0 -1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _2338_
timestamp 1644511149
transform 1 0 31280 0 1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__and3_1  _2339_
timestamp 1644511149
transform 1 0 43700 0 -1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _2340_
timestamp 1644511149
transform -1 0 43976 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__a211oi_2  _2341_
timestamp 1644511149
transform -1 0 45172 0 -1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__o211a_1  _2342_
timestamp 1644511149
transform -1 0 45724 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__a211oi_1  _2343_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 45724 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _2344_
timestamp 1644511149
transform -1 0 46552 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2345_
timestamp 1644511149
transform 1 0 47564 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2346_
timestamp 1644511149
transform -1 0 45356 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _2347_
timestamp 1644511149
transform 1 0 44712 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _2348_
timestamp 1644511149
transform 1 0 47196 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2349_
timestamp 1644511149
transform 1 0 49220 0 -1 29376
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2350_
timestamp 1644511149
transform -1 0 47932 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_1  _2351_
timestamp 1644511149
transform 1 0 48300 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _2352_
timestamp 1644511149
transform 1 0 48116 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_1  _2353_
timestamp 1644511149
transform 1 0 49312 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _2354_
timestamp 1644511149
transform 1 0 48392 0 -1 32640
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_4  _2355_
timestamp 1644511149
transform -1 0 50416 0 -1 33728
box -38 -48 2062 592
use sky130_fd_sc_hd__xor2_2  _2356_
timestamp 1644511149
transform -1 0 48760 0 1 34816
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _2357_
timestamp 1644511149
transform -1 0 49036 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  _2358_
timestamp 1644511149
transform 1 0 48484 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__a31o_1  _2359_
timestamp 1644511149
transform -1 0 48944 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_1  _2360_
timestamp 1644511149
transform 1 0 43516 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_4  _2361_
timestamp 1644511149
transform 1 0 12420 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _2362_
timestamp 1644511149
transform -1 0 8004 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2363_
timestamp 1644511149
transform -1 0 7728 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2364_
timestamp 1644511149
transform 1 0 8924 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_4  _2365_
timestamp 1644511149
transform -1 0 11040 0 -1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__and3_2  _2366_
timestamp 1644511149
transform 1 0 10212 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__or3_1  _2367_
timestamp 1644511149
transform 1 0 33028 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _2368_
timestamp 1644511149
transform -1 0 26220 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _2369_
timestamp 1644511149
transform 1 0 27600 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _2370_
timestamp 1644511149
transform -1 0 28520 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2371_
timestamp 1644511149
transform -1 0 27508 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _2372_
timestamp 1644511149
transform -1 0 34040 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _2373_
timestamp 1644511149
transform -1 0 35052 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _2374_
timestamp 1644511149
transform 1 0 33856 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _2375_
timestamp 1644511149
transform 1 0 31280 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _2376_
timestamp 1644511149
transform 1 0 32108 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2377_
timestamp 1644511149
transform -1 0 33304 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__and3_1  _2378_
timestamp 1644511149
transform 1 0 32660 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _2379_
timestamp 1644511149
transform 1 0 32292 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _2380_
timestamp 1644511149
transform 1 0 34316 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _2381_
timestamp 1644511149
transform -1 0 34224 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_2  _2382_
timestamp 1644511149
transform -1 0 35052 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _2383_
timestamp 1644511149
transform 1 0 34684 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_1  _2384_
timestamp 1644511149
transform 1 0 44896 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _2385_
timestamp 1644511149
transform -1 0 45540 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _2386_
timestamp 1644511149
transform 1 0 35420 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _2387_
timestamp 1644511149
transform 1 0 20240 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _2388_
timestamp 1644511149
transform 1 0 20516 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2389_
timestamp 1644511149
transform 1 0 21528 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _2390_
timestamp 1644511149
transform 1 0 36800 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _2391_
timestamp 1644511149
transform 1 0 34316 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _2392_
timestamp 1644511149
transform 1 0 20976 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  _2393_
timestamp 1644511149
transform -1 0 21344 0 -1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__or2_4  _2394_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 9476 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2395_
timestamp 1644511149
transform 1 0 24380 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2396_
timestamp 1644511149
transform -1 0 24656 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _2397_
timestamp 1644511149
transform 1 0 23000 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _2398_
timestamp 1644511149
transform 1 0 35880 0 1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _2399_
timestamp 1644511149
transform 1 0 38088 0 -1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_2  _2400_
timestamp 1644511149
transform 1 0 40204 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _2401_
timestamp 1644511149
transform 1 0 19228 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2402_
timestamp 1644511149
transform 1 0 19320 0 1 19584
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  _2403_
timestamp 1644511149
transform -1 0 20332 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _2404_
timestamp 1644511149
transform 1 0 18216 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_2  _2405_
timestamp 1644511149
transform 1 0 19228 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _2406_
timestamp 1644511149
transform 1 0 40296 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _2407_
timestamp 1644511149
transform 1 0 41860 0 1 20672
box -38 -48 1234 592
use sky130_fd_sc_hd__nand3_1  _2408_
timestamp 1644511149
transform -1 0 46920 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _2409_
timestamp 1644511149
transform -1 0 46184 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _2410_
timestamp 1644511149
transform 1 0 46276 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _2411_
timestamp 1644511149
transform -1 0 46552 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _2412_
timestamp 1644511149
transform 1 0 47564 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _2413_
timestamp 1644511149
transform 1 0 27600 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _2414_
timestamp 1644511149
transform 1 0 30360 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _2415_
timestamp 1644511149
transform 1 0 6348 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _2416_
timestamp 1644511149
transform 1 0 7084 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _2417_
timestamp 1644511149
transform 1 0 30912 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _2418_
timestamp 1644511149
transform 1 0 30728 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2419_
timestamp 1644511149
transform 1 0 46828 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _2420_
timestamp 1644511149
transform 1 0 47748 0 1 23936
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _2421_
timestamp 1644511149
transform -1 0 47104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _2422_
timestamp 1644511149
transform -1 0 49588 0 -1 26112
box -38 -48 1234 592
use sky130_fd_sc_hd__and2b_1  _2423_
timestamp 1644511149
transform 1 0 48208 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2424_
timestamp 1644511149
transform -1 0 48576 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _2425_
timestamp 1644511149
transform 1 0 48208 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _2426_
timestamp 1644511149
transform 1 0 48484 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2427_
timestamp 1644511149
transform 1 0 49128 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _2428_
timestamp 1644511149
transform 1 0 49220 0 1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2429_
timestamp 1644511149
transform -1 0 49496 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _2430_
timestamp 1644511149
transform -1 0 49220 0 1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__a311o_1  _2431_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 49036 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _2432_
timestamp 1644511149
transform 1 0 49404 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2433_
timestamp 1644511149
transform -1 0 50232 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _2434_
timestamp 1644511149
transform -1 0 47840 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__a21boi_2  _2435_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 45816 0 -1 21760
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _2436_
timestamp 1644511149
transform 1 0 32476 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2437_
timestamp 1644511149
transform 1 0 35972 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _2438_
timestamp 1644511149
transform 1 0 36432 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _2439_
timestamp 1644511149
transform -1 0 36340 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _2440_
timestamp 1644511149
transform -1 0 36616 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _2441_
timestamp 1644511149
transform 1 0 6808 0 1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__inv_2  _2442_
timestamp 1644511149
transform -1 0 7084 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__a2111o_1  _2443_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 8004 0 1 18496
box -38 -48 866 592
use sky130_fd_sc_hd__nand2_1  _2444_
timestamp 1644511149
transform -1 0 9200 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__and3_1  _2445_
timestamp 1644511149
transform 1 0 8096 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2446_
timestamp 1644511149
transform -1 0 10856 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2447_
timestamp 1644511149
transform -1 0 10304 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2448_
timestamp 1644511149
transform -1 0 9476 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _2449_
timestamp 1644511149
transform -1 0 9568 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _2450_
timestamp 1644511149
transform 1 0 9200 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  _2451_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 9936 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _2452_
timestamp 1644511149
transform -1 0 28428 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _2453_
timestamp 1644511149
transform -1 0 30176 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2454_
timestamp 1644511149
transform -1 0 29440 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _2455_
timestamp 1644511149
transform -1 0 30912 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _2456_
timestamp 1644511149
transform 1 0 38272 0 -1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _2457_
timestamp 1644511149
transform 1 0 44620 0 -1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _2458_
timestamp 1644511149
transform 1 0 45448 0 -1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_2  _2459_
timestamp 1644511149
transform -1 0 22172 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _2460_
timestamp 1644511149
transform 1 0 24380 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2461_
timestamp 1644511149
transform -1 0 25024 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_2  _2462_
timestamp 1644511149
transform 1 0 25576 0 1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_2  _2463_
timestamp 1644511149
transform -1 0 23460 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _2464_
timestamp 1644511149
transform 1 0 21620 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_2  _2465_
timestamp 1644511149
transform 1 0 21804 0 -1 19584
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _2466_
timestamp 1644511149
transform 1 0 37904 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _2467_
timestamp 1644511149
transform 1 0 40204 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2468_
timestamp 1644511149
transform 1 0 19688 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2469_
timestamp 1644511149
transform -1 0 19320 0 -1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _2470_
timestamp 1644511149
transform -1 0 17940 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _2471_
timestamp 1644511149
transform 1 0 19504 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_2  _2472_
timestamp 1644511149
transform 1 0 20148 0 1 17408
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _2473_
timestamp 1644511149
transform 1 0 40756 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2474_
timestamp 1644511149
transform 1 0 41676 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2475_
timestamp 1644511149
transform 1 0 42320 0 1 18496
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2476_
timestamp 1644511149
transform 1 0 43792 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_2  _2477_
timestamp 1644511149
transform 1 0 46460 0 1 19584
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _2478_
timestamp 1644511149
transform 1 0 47932 0 -1 21760
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_1  _2479_
timestamp 1644511149
transform 1 0 38272 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__and2b_1  _2480_
timestamp 1644511149
transform 1 0 42412 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _2481_
timestamp 1644511149
transform 1 0 6716 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__and2b_1  _2482_
timestamp 1644511149
transform 1 0 12420 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  _2483_
timestamp 1644511149
transform 1 0 14260 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__o21bai_1  _2484_
timestamp 1644511149
transform 1 0 7360 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_4  _2485_
timestamp 1644511149
transform -1 0 8004 0 1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _2486_
timestamp 1644511149
transform 1 0 12880 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2487_
timestamp 1644511149
transform -1 0 14352 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_4  _2488_
timestamp 1644511149
transform -1 0 16008 0 -1 19584
box -38 -48 1602 592
use sky130_fd_sc_hd__o21ai_2  _2489_
timestamp 1644511149
transform 1 0 43424 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _2490_
timestamp 1644511149
transform 1 0 43332 0 -1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2491_
timestamp 1644511149
transform 1 0 49220 0 1 20672
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_2  _2492_
timestamp 1644511149
transform 1 0 49220 0 -1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _2493_
timestamp 1644511149
transform 1 0 50140 0 1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _2494_
timestamp 1644511149
transform -1 0 51244 0 -1 25024
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_1  _2495_
timestamp 1644511149
transform 1 0 50140 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2496_
timestamp 1644511149
transform -1 0 49404 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2497_
timestamp 1644511149
transform -1 0 50968 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _2498_
timestamp 1644511149
transform 1 0 51060 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _2499_
timestamp 1644511149
transform 1 0 52072 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _2500_
timestamp 1644511149
transform -1 0 51520 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _2501_
timestamp 1644511149
transform 1 0 51244 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _2502_
timestamp 1644511149
transform -1 0 53084 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2503_
timestamp 1644511149
transform 1 0 52716 0 -1 33728
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2504_
timestamp 1644511149
transform 1 0 53452 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__o211ai_4  _2505_
timestamp 1644511149
transform 1 0 49220 0 -1 34816
box -38 -48 1602 592
use sky130_fd_sc_hd__nand2_1  _2506_
timestamp 1644511149
transform 1 0 51980 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _2507_
timestamp 1644511149
transform 1 0 52992 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _2508_
timestamp 1644511149
transform 1 0 51152 0 1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2509_
timestamp 1644511149
transform -1 0 50600 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2510_
timestamp 1644511149
transform 1 0 50968 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _2511_
timestamp 1644511149
transform 1 0 48300 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _2512_
timestamp 1644511149
transform 1 0 49680 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2513_
timestamp 1644511149
transform -1 0 46092 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2514_
timestamp 1644511149
transform 1 0 47564 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _2515_
timestamp 1644511149
transform 1 0 37260 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_2  _2516_
timestamp 1644511149
transform 1 0 37260 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2517_
timestamp 1644511149
transform 1 0 42780 0 -1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_1  _2518_
timestamp 1644511149
transform 1 0 26956 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2519_
timestamp 1644511149
transform -1 0 26312 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_2  _2520_
timestamp 1644511149
transform 1 0 25852 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__and3_1  _2521_
timestamp 1644511149
transform 1 0 11500 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__buf_2  _2522_
timestamp 1644511149
transform 1 0 10672 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _2523_
timestamp 1644511149
transform -1 0 12696 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__or3_4  _2524_
timestamp 1644511149
transform 1 0 13248 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  _2525_
timestamp 1644511149
transform 1 0 29900 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _2526_
timestamp 1644511149
transform 1 0 30636 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _2527_
timestamp 1644511149
transform 1 0 31004 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _2528_
timestamp 1644511149
transform 1 0 30820 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _2529_
timestamp 1644511149
transform 1 0 42872 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _2530_
timestamp 1644511149
transform -1 0 43056 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _2531_
timestamp 1644511149
transform 1 0 43884 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _2532_
timestamp 1644511149
transform -1 0 44068 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__or2b_1  _2533_
timestamp 1644511149
transform 1 0 44988 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _2534_
timestamp 1644511149
transform 1 0 44160 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _2535_
timestamp 1644511149
transform 1 0 45264 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _2536_
timestamp 1644511149
transform -1 0 24840 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _2537_
timestamp 1644511149
transform 1 0 28152 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__and2_2  _2538_
timestamp 1644511149
transform 1 0 12420 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _2539_
timestamp 1644511149
transform 1 0 25852 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2540_
timestamp 1644511149
transform -1 0 28428 0 1 16320
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _2541_
timestamp 1644511149
transform -1 0 27784 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2542_
timestamp 1644511149
transform 1 0 26404 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_2  _2543_
timestamp 1644511149
transform 1 0 35972 0 1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_2  _2544_
timestamp 1644511149
transform 1 0 22540 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _2545_
timestamp 1644511149
transform -1 0 23920 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _2546_
timestamp 1644511149
transform -1 0 23828 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _2547_
timestamp 1644511149
transform -1 0 23460 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_2  _2548_
timestamp 1644511149
transform 1 0 23000 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _2549_
timestamp 1644511149
transform 1 0 38456 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _2550_
timestamp 1644511149
transform 1 0 45724 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _2551_
timestamp 1644511149
transform 1 0 19412 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2552_
timestamp 1644511149
transform 1 0 20516 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _2553_
timestamp 1644511149
transform 1 0 17020 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _2554_
timestamp 1644511149
transform -1 0 18308 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _2555_
timestamp 1644511149
transform -1 0 21344 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_2  _2556_
timestamp 1644511149
transform 1 0 19596 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _2557_
timestamp 1644511149
transform 1 0 40572 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _2558_
timestamp 1644511149
transform 1 0 47932 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _2559_
timestamp 1644511149
transform -1 0 48576 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _2560_
timestamp 1644511149
transform -1 0 49404 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o211ai_1  _2561_
timestamp 1644511149
transform 1 0 50416 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _2562_
timestamp 1644511149
transform -1 0 50048 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2563_
timestamp 1644511149
transform 1 0 40480 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _2564_
timestamp 1644511149
transform 1 0 15456 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  _2565_
timestamp 1644511149
transform 1 0 21160 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _2566_
timestamp 1644511149
transform -1 0 14904 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a2bb2o_1  _2567_
timestamp 1644511149
transform 1 0 13340 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a221oi_4  _2568_
timestamp 1644511149
transform 1 0 14352 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__a21oi_2  _2569_
timestamp 1644511149
transform 1 0 42780 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _2570_
timestamp 1644511149
transform 1 0 42964 0 1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2571_
timestamp 1644511149
transform 1 0 48760 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__and3_2  _2572_
timestamp 1644511149
transform 1 0 51336 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _2573_
timestamp 1644511149
transform -1 0 50784 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__a211oi_4  _2574_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 50968 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__o211a_1  _2575_
timestamp 1644511149
transform -1 0 51888 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__nor3_2  _2576_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 52716 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__o21a_1  _2577_
timestamp 1644511149
transform -1 0 52256 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_4  _2578_
timestamp 1644511149
transform 1 0 52072 0 1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__o211a_1  _2579_
timestamp 1644511149
transform -1 0 53452 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _2580_
timestamp 1644511149
transform 1 0 50140 0 1 25024
box -38 -48 498 592
use sky130_fd_sc_hd__o21a_1  _2581_
timestamp 1644511149
transform -1 0 53268 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2582_
timestamp 1644511149
transform -1 0 53268 0 -1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__nor3_2  _2583_
timestamp 1644511149
transform 1 0 52624 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__o211ai_1  _2584_
timestamp 1644511149
transform -1 0 53268 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _2585_
timestamp 1644511149
transform 1 0 53636 0 -1 26112
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _2586_
timestamp 1644511149
transform -1 0 53176 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__or2_2  _2587_
timestamp 1644511149
transform 1 0 53360 0 -1 27200
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _2588_
timestamp 1644511149
transform -1 0 51796 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__a31oi_4  _2589_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 52164 0 1 33728
box -38 -48 1602 592
use sky130_fd_sc_hd__xor2_4  _2590_
timestamp 1644511149
transform -1 0 54832 0 1 27200
box -38 -48 2062 592
use sky130_fd_sc_hd__inv_2  _2591_
timestamp 1644511149
transform 1 0 54556 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__a31o_1  _2592_
timestamp 1644511149
transform -1 0 56028 0 1 25024
box -38 -48 682 592
use sky130_fd_sc_hd__o211a_1  _2593_
timestamp 1644511149
transform -1 0 50876 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_1  _2594_
timestamp 1644511149
transform 1 0 48944 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _2595_
timestamp 1644511149
transform 1 0 32476 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _2596_
timestamp 1644511149
transform -1 0 25116 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _2597_
timestamp 1644511149
transform 1 0 28520 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _2598_
timestamp 1644511149
transform -1 0 30176 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _2599_
timestamp 1644511149
transform -1 0 37996 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _2600_
timestamp 1644511149
transform -1 0 39192 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nand3_2  _2601_
timestamp 1644511149
transform -1 0 38456 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__a22o_1  _2602_
timestamp 1644511149
transform 1 0 23276 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2603_
timestamp 1644511149
transform -1 0 23920 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _2604_
timestamp 1644511149
transform -1 0 24932 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _2605_
timestamp 1644511149
transform 1 0 38364 0 -1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__a21o_1  _2606_
timestamp 1644511149
transform -1 0 49956 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _2607_
timestamp 1644511149
transform 1 0 48668 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _2608_
timestamp 1644511149
transform 1 0 19228 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_2  _2609_
timestamp 1644511149
transform 1 0 19596 0 -1 16320
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _2610_
timestamp 1644511149
transform 1 0 40388 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _2611_
timestamp 1644511149
transform 1 0 50324 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _2612_
timestamp 1644511149
transform -1 0 50508 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_2  _2613_
timestamp 1644511149
transform -1 0 10212 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_2  _2614_
timestamp 1644511149
transform 1 0 33028 0 -1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__nand4_1  _2615_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 32568 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _2616_
timestamp 1644511149
transform 1 0 32108 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _2617_
timestamp 1644511149
transform -1 0 32568 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _2618_
timestamp 1644511149
transform 1 0 33212 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_2  _2619_
timestamp 1644511149
transform -1 0 35328 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__a21o_1  _2620_
timestamp 1644511149
transform -1 0 44804 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _2621_
timestamp 1644511149
transform 1 0 45172 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _2622_
timestamp 1644511149
transform 1 0 46276 0 -1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _2623_
timestamp 1644511149
transform -1 0 44712 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_1  _2624_
timestamp 1644511149
transform 1 0 47196 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _2625_
timestamp 1644511149
transform 1 0 52716 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _2626_
timestamp 1644511149
transform 1 0 52716 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2627_
timestamp 1644511149
transform -1 0 54556 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _2628_
timestamp 1644511149
transform 1 0 52716 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__and2_1  _2629_
timestamp 1644511149
transform 1 0 46736 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2630_
timestamp 1644511149
transform 1 0 48944 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _2631_
timestamp 1644511149
transform 1 0 14444 0 -1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2632_
timestamp 1644511149
transform 1 0 14076 0 1 15232
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _2633_
timestamp 1644511149
transform 1 0 14076 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _2634_
timestamp 1644511149
transform 1 0 14996 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_2  _2635_
timestamp 1644511149
transform 1 0 50232 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _2636_
timestamp 1644511149
transform 1 0 51244 0 -1 17408
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2637_
timestamp 1644511149
transform 1 0 51796 0 1 16320
box -38 -48 498 592
use sky130_fd_sc_hd__or3b_1  _2638_
timestamp 1644511149
transform -1 0 54004 0 1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__o21bai_1  _2639_
timestamp 1644511149
transform 1 0 53176 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__o211ai_1  _2640_
timestamp 1644511149
transform 1 0 52256 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__a211o_1  _2641_
timestamp 1644511149
transform -1 0 53820 0 1 18496
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _2642_
timestamp 1644511149
transform -1 0 54740 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _2643_
timestamp 1644511149
transform -1 0 54004 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__o211ai_1  _2644_
timestamp 1644511149
transform 1 0 53820 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _2645_
timestamp 1644511149
transform -1 0 55844 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_1  _2646_
timestamp 1644511149
transform -1 0 54464 0 -1 21760
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2647_
timestamp 1644511149
transform -1 0 54832 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2648_
timestamp 1644511149
transform 1 0 55292 0 1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2649_
timestamp 1644511149
transform 1 0 55936 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _2650_
timestamp 1644511149
transform 1 0 55660 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2651_
timestamp 1644511149
transform 1 0 56396 0 1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__o21ba_1  _2652_
timestamp 1644511149
transform -1 0 56028 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _2653_
timestamp 1644511149
transform 1 0 56764 0 -1 27200
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _2654_
timestamp 1644511149
transform -1 0 55936 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__o211ai_2  _2655_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 55384 0 -1 22848
box -38 -48 958 592
use sky130_fd_sc_hd__nand2_2  _2656_
timestamp 1644511149
transform 1 0 56120 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__a21bo_1  _2657_
timestamp 1644511149
transform 1 0 53544 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _2658_
timestamp 1644511149
transform -1 0 53728 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _2659_
timestamp 1644511149
transform 1 0 53452 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_1  _2660_
timestamp 1644511149
transform 1 0 46276 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__o31a_1  _2661_
timestamp 1644511149
transform -1 0 53360 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2662_
timestamp 1644511149
transform 1 0 28336 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2663_
timestamp 1644511149
transform -1 0 29256 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _2664_
timestamp 1644511149
transform -1 0 30544 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_1  _2665_
timestamp 1644511149
transform 1 0 37996 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_4  _2666_
timestamp 1644511149
transform -1 0 36616 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _2667_
timestamp 1644511149
transform -1 0 25024 0 1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_2  _2668_
timestamp 1644511149
transform -1 0 24840 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_2  _2669_
timestamp 1644511149
transform 1 0 35144 0 1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _2670_
timestamp 1644511149
transform 1 0 40572 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _2671_
timestamp 1644511149
transform -1 0 41032 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _2672_
timestamp 1644511149
transform -1 0 20608 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _2673_
timestamp 1644511149
transform -1 0 21528 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _2674_
timestamp 1644511149
transform 1 0 19872 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_2  _2675_
timestamp 1644511149
transform 1 0 20056 0 -1 15232
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _2676_
timestamp 1644511149
transform 1 0 40572 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _2677_
timestamp 1644511149
transform 1 0 42228 0 1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__a21o_1  _2678_
timestamp 1644511149
transform -1 0 46368 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__and3_2  _2679_
timestamp 1644511149
transform 1 0 33028 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _2680_
timestamp 1644511149
transform 1 0 34316 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_2  _2681_
timestamp 1644511149
transform 1 0 33304 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a2111oi_4  _2682_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 36708 0 1 14144
box -38 -48 2062 592
use sky130_fd_sc_hd__a22o_1  _2683_
timestamp 1644511149
transform 1 0 36064 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_1  _2684_
timestamp 1644511149
transform 1 0 43884 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__or3_1  _2685_
timestamp 1644511149
transform 1 0 43976 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2686_
timestamp 1644511149
transform 1 0 44988 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_2  _2687_
timestamp 1644511149
transform 1 0 46552 0 1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _2688_
timestamp 1644511149
transform 1 0 48208 0 1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _2689_
timestamp 1644511149
transform 1 0 52716 0 -1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_1  _2690_
timestamp 1644511149
transform -1 0 50508 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _2691_
timestamp 1644511149
transform 1 0 15088 0 -1 17408
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2692_
timestamp 1644511149
transform 1 0 14168 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _2693_
timestamp 1644511149
transform 1 0 15272 0 1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_2  _2694_
timestamp 1644511149
transform 1 0 53728 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _2695_
timestamp 1644511149
transform 1 0 53360 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2696_
timestamp 1644511149
transform 1 0 54372 0 1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _2697_
timestamp 1644511149
transform 1 0 55660 0 1 14144
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _2698_
timestamp 1644511149
transform 1 0 56120 0 1 16320
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _2699_
timestamp 1644511149
transform 1 0 56212 0 -1 17408
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _2700_
timestamp 1644511149
transform 1 0 56304 0 1 18496
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_1  _2701_
timestamp 1644511149
transform 1 0 56120 0 -1 21760
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2702_
timestamp 1644511149
transform -1 0 57224 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_2  _2703_
timestamp 1644511149
transform 1 0 56948 0 -1 22848
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_4  _2704_
timestamp 1644511149
transform 1 0 56212 0 1 22848
box -38 -48 2062 592
use sky130_fd_sc_hd__xnor2_2  _2705_
timestamp 1644511149
transform -1 0 56120 0 -1 29376
box -38 -48 1234 592
use sky130_fd_sc_hd__a21oi_1  _2706_
timestamp 1644511149
transform 1 0 55660 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2707_
timestamp 1644511149
transform 1 0 55936 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o32a_1  _2708_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 55292 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__or2_1  _2709_
timestamp 1644511149
transform -1 0 55568 0 -1 30464
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2710_
timestamp 1644511149
transform -1 0 56212 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__and2_4  _2711_
timestamp 1644511149
transform -1 0 55568 0 -1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  _2712_
timestamp 1644511149
transform 1 0 2484 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2713_
timestamp 1644511149
transform -1 0 56856 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _2714_
timestamp 1644511149
transform 1 0 52992 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _2715_
timestamp 1644511149
transform -1 0 55568 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _2716_
timestamp 1644511149
transform -1 0 45540 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _2717_
timestamp 1644511149
transform 1 0 37628 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _2718_
timestamp 1644511149
transform -1 0 37628 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _2719_
timestamp 1644511149
transform 1 0 38548 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _2720_
timestamp 1644511149
transform -1 0 39284 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2721_
timestamp 1644511149
transform -1 0 42412 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _2722_
timestamp 1644511149
transform 1 0 44804 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__or3_2  _2723_
timestamp 1644511149
transform 1 0 13340 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2724_
timestamp 1644511149
transform 1 0 29072 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _2725_
timestamp 1644511149
transform -1 0 30268 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2726_
timestamp 1644511149
transform 1 0 29808 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _2727_
timestamp 1644511149
transform -1 0 38272 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _2728_
timestamp 1644511149
transform 1 0 38640 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _2729_
timestamp 1644511149
transform -1 0 28336 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _2730_
timestamp 1644511149
transform 1 0 24380 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _2731_
timestamp 1644511149
transform 1 0 24472 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2732_
timestamp 1644511149
transform 1 0 24840 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_2  _2733_
timestamp 1644511149
transform 1 0 25944 0 1 13056
box -38 -48 1234 592
use sky130_fd_sc_hd__a21o_1  _2734_
timestamp 1644511149
transform -1 0 38732 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__nand3_1  _2735_
timestamp 1644511149
transform -1 0 38732 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _2736_
timestamp 1644511149
transform -1 0 20240 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _2737_
timestamp 1644511149
transform 1 0 20884 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _2738_
timestamp 1644511149
transform 1 0 21620 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _2739_
timestamp 1644511149
transform -1 0 20792 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _2740_
timestamp 1644511149
transform 1 0 20700 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_2  _2741_
timestamp 1644511149
transform 1 0 21804 0 -1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_1  _2742_
timestamp 1644511149
transform 1 0 40940 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_2  _2743_
timestamp 1644511149
transform -1 0 43884 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_1  _2744_
timestamp 1644511149
transform -1 0 43700 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _2745_
timestamp 1644511149
transform 1 0 45908 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__a21oi_1  _2746_
timestamp 1644511149
transform -1 0 46092 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2747_
timestamp 1644511149
transform -1 0 46828 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2748_
timestamp 1644511149
transform 1 0 47564 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nor3b_1  _2749_
timestamp 1644511149
transform -1 0 49128 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2750_
timestamp 1644511149
transform -1 0 49312 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__and2b_1  _2751_
timestamp 1644511149
transform -1 0 42964 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a21oi_2  _2752_
timestamp 1644511149
transform 1 0 41124 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2753_
timestamp 1644511149
transform 1 0 15088 0 1 15232
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _2754_
timestamp 1644511149
transform 1 0 14168 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2755_
timestamp 1644511149
transform -1 0 16192 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__a221o_1  _2756_
timestamp 1644511149
transform 1 0 16376 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__a21oi_4  _2757_
timestamp 1644511149
transform -1 0 17848 0 -1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _2758_
timestamp 1644511149
transform 1 0 50600 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nor3_1  _2759_
timestamp 1644511149
transform -1 0 51520 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _2760_
timestamp 1644511149
transform -1 0 52164 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_1  _2761_
timestamp 1644511149
transform -1 0 54648 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__o211a_1  _2762_
timestamp 1644511149
transform -1 0 55752 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__or3_1  _2763_
timestamp 1644511149
transform 1 0 56764 0 1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _2764_
timestamp 1644511149
transform 1 0 56580 0 -1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _2765_
timestamp 1644511149
transform -1 0 58144 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_1  _2766_
timestamp 1644511149
transform -1 0 56856 0 -1 16320
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _2767_
timestamp 1644511149
transform 1 0 56580 0 1 15232
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _2768_
timestamp 1644511149
transform 1 0 57868 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2769_
timestamp 1644511149
transform 1 0 56764 0 -1 19584
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2770_
timestamp 1644511149
transform 1 0 57868 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2771_
timestamp 1644511149
transform 1 0 57868 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__a21oi_1  _2772_
timestamp 1644511149
transform -1 0 57040 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__or2_1  _2773_
timestamp 1644511149
transform -1 0 56764 0 1 23936
box -38 -48 498 592
use sky130_fd_sc_hd__a311o_1  _2774_
timestamp 1644511149
transform -1 0 56120 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__nand3_1  _2775_
timestamp 1644511149
transform -1 0 58236 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _2776_
timestamp 1644511149
transform -1 0 57408 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__and3_1  _2777_
timestamp 1644511149
transform -1 0 57408 0 -1 28288
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _2778_
timestamp 1644511149
transform -1 0 57684 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__or2b_2  _2779_
timestamp 1644511149
transform -1 0 57408 0 -1 29376
box -38 -48 682 592
use sky130_fd_sc_hd__a21boi_1  _2780_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 55292 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_2  _2781_
timestamp 1644511149
transform -1 0 56488 0 1 31552
box -38 -48 1234 592
use sky130_fd_sc_hd__a221o_1  _2782_
timestamp 1644511149
transform -1 0 56948 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__o31a_1  _2783_
timestamp 1644511149
transform 1 0 56488 0 1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__nand2_1  _2784_
timestamp 1644511149
transform -1 0 57316 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2785_
timestamp 1644511149
transform 1 0 56764 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o21bai_2  _2786_
timestamp 1644511149
transform 1 0 56304 0 -1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__nor2_2  _2787_
timestamp 1644511149
transform 1 0 50784 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or2_2  _2788_
timestamp 1644511149
transform -1 0 52348 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__a31o_1  _2789_
timestamp 1644511149
transform -1 0 46460 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _2790_
timestamp 1644511149
transform 1 0 39100 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2791_
timestamp 1644511149
transform 1 0 38548 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2792_
timestamp 1644511149
transform -1 0 41952 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__a21o_1  _2793_
timestamp 1644511149
transform -1 0 32752 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _2794_
timestamp 1644511149
transform -1 0 30728 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _2795_
timestamp 1644511149
transform -1 0 31188 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2796_
timestamp 1644511149
transform -1 0 30912 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _2797_
timestamp 1644511149
transform -1 0 34868 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2798_
timestamp 1644511149
transform 1 0 34684 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or3_1  _2799_
timestamp 1644511149
transform 1 0 32476 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  _2800_
timestamp 1644511149
transform 1 0 25484 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _2801_
timestamp 1644511149
transform 1 0 24932 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _2802_
timestamp 1644511149
transform -1 0 30176 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2803_
timestamp 1644511149
transform -1 0 29072 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a21oi_1  _2804_
timestamp 1644511149
transform -1 0 34040 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__and3_1  _2805_
timestamp 1644511149
transform 1 0 33580 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__or4_2  _2806_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 34868 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__o22ai_2  _2807_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 34684 0 1 10880
box -38 -48 958 592
use sky130_fd_sc_hd__nor2_1  _2808_
timestamp 1644511149
transform -1 0 20148 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _2809_
timestamp 1644511149
transform -1 0 22264 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _2810_
timestamp 1644511149
transform -1 0 21804 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_2  _2811_
timestamp 1644511149
transform -1 0 20792 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_1  _2812_
timestamp 1644511149
transform 1 0 40480 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__nand3_1  _2813_
timestamp 1644511149
transform 1 0 40940 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_1  _2814_
timestamp 1644511149
transform 1 0 41676 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_1  _2815_
timestamp 1644511149
transform 1 0 41676 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_2  _2816_
timestamp 1644511149
transform 1 0 42504 0 -1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _2817_
timestamp 1644511149
transform 1 0 47564 0 -1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _2818_
timestamp 1644511149
transform -1 0 49404 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2819_
timestamp 1644511149
transform 1 0 16652 0 -1 14144
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _2820_
timestamp 1644511149
transform 1 0 15272 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _2821_
timestamp 1644511149
transform 1 0 17480 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _2822_
timestamp 1644511149
transform 1 0 14536 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _2823_
timestamp 1644511149
transform 1 0 15732 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _2824_
timestamp 1644511149
transform 1 0 18584 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_4  _2825_
timestamp 1644511149
transform 1 0 19228 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_2  _2826_
timestamp 1644511149
transform 1 0 48484 0 -1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _2827_
timestamp 1644511149
transform 1 0 49220 0 -1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _2828_
timestamp 1644511149
transform 1 0 51060 0 -1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _2829_
timestamp 1644511149
transform 1 0 52716 0 -1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _2830_
timestamp 1644511149
transform 1 0 56120 0 1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__nor2_1  _2831_
timestamp 1644511149
transform -1 0 57592 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2832_
timestamp 1644511149
transform -1 0 57224 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2833_
timestamp 1644511149
transform 1 0 56764 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__xnor2_2  _2834_
timestamp 1644511149
transform -1 0 57408 0 -1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_2  _2835_
timestamp 1644511149
transform 1 0 55936 0 1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__a31oi_2  _2836_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 58144 0 1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__o31ai_4  _2837_
timestamp 1644511149
transform 1 0 55292 0 1 29376
box -38 -48 1602 592
use sky130_fd_sc_hd__xor2_1  _2838_
timestamp 1644511149
transform 1 0 56764 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _2839_
timestamp 1644511149
transform -1 0 56396 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2840_
timestamp 1644511149
transform -1 0 48760 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__and2b_1  _2841_
timestamp 1644511149
transform 1 0 47748 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__a21o_1  _2842_
timestamp 1644511149
transform 1 0 48668 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__o21ba_1  _2843_
timestamp 1644511149
transform -1 0 43056 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  _2844_
timestamp 1644511149
transform -1 0 21344 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _2845_
timestamp 1644511149
transform 1 0 21712 0 1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_2  _2846_
timestamp 1644511149
transform 1 0 22356 0 -1 11968
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_2  _2847_
timestamp 1644511149
transform 1 0 37260 0 -1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_4  _2848_
timestamp 1644511149
transform 1 0 12052 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a22o_1  _2849_
timestamp 1644511149
transform 1 0 29164 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2850_
timestamp 1644511149
transform -1 0 30544 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _2851_
timestamp 1644511149
transform -1 0 31740 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _2852_
timestamp 1644511149
transform 1 0 32568 0 1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_4  _2853_
timestamp 1644511149
transform -1 0 36800 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__a211oi_4  _2854_
timestamp 1644511149
transform -1 0 35696 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__a22o_1  _2855_
timestamp 1644511149
transform -1 0 28612 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2856_
timestamp 1644511149
transform -1 0 28152 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__xnor2_1  _2857_
timestamp 1644511149
transform 1 0 32200 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__xor2_2  _2858_
timestamp 1644511149
transform 1 0 34684 0 1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _2859_
timestamp 1644511149
transform 1 0 37444 0 -1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_1  _2860_
timestamp 1644511149
transform 1 0 42412 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _2861_
timestamp 1644511149
transform 1 0 44896 0 -1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__a22o_1  _2862_
timestamp 1644511149
transform 1 0 15732 0 1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2863_
timestamp 1644511149
transform 1 0 15548 0 -1 15232
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_4  _2864_
timestamp 1644511149
transform 1 0 16744 0 1 14144
box -38 -48 866 592
use sky130_fd_sc_hd__a21oi_2  _2865_
timestamp 1644511149
transform 1 0 42596 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and3_1  _2866_
timestamp 1644511149
transform 1 0 42688 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2867_
timestamp 1644511149
transform 1 0 43976 0 -1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__xor2_1  _2868_
timestamp 1644511149
transform 1 0 45816 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2869_
timestamp 1644511149
transform 1 0 48300 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2870_
timestamp 1644511149
transform 1 0 49036 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__a22oi_2  _2871_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 52532 0 1 7616
box -38 -48 958 592
use sky130_fd_sc_hd__xor2_1  _2872_
timestamp 1644511149
transform 1 0 51520 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_1  _2873_
timestamp 1644511149
transform 1 0 55108 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  _2874_
timestamp 1644511149
transform 1 0 54280 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2b_1  _2875_
timestamp 1644511149
transform 1 0 54004 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__o21ai_1  _2876_
timestamp 1644511149
transform 1 0 56764 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_2  _2877_
timestamp 1644511149
transform 1 0 56672 0 -1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _2878_
timestamp 1644511149
transform 1 0 57960 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__o21ba_1  _2879_
timestamp 1644511149
transform 1 0 56212 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _2880_
timestamp 1644511149
transform -1 0 54740 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _2881_
timestamp 1644511149
transform 1 0 54280 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2882_
timestamp 1644511149
transform 1 0 53728 0 -1 6528
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _2883_
timestamp 1644511149
transform 1 0 55936 0 -1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__a21o_1  _2884_
timestamp 1644511149
transform -1 0 57316 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__xor2_1  _2885_
timestamp 1644511149
transform 1 0 56764 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__or2_1  _2886_
timestamp 1644511149
transform 1 0 55936 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2887_
timestamp 1644511149
transform 1 0 56212 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_1  _2888_
timestamp 1644511149
transform -1 0 55936 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__o211a_4  _2889_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 56028 0 -1 11968
box -38 -48 1326 592
use sky130_fd_sc_hd__nor2_1  _2890_
timestamp 1644511149
transform -1 0 51704 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__or2_1  _2891_
timestamp 1644511149
transform 1 0 45172 0 1 6528
box -38 -48 498 592
use sky130_fd_sc_hd__o21ai_4  _2892_
timestamp 1644511149
transform -1 0 46552 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__and2_1  _2893_
timestamp 1644511149
transform 1 0 34408 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2894_
timestamp 1644511149
transform -1 0 37904 0 1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__a22o_1  _2895_
timestamp 1644511149
transform 1 0 16008 0 1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__a22o_1  _2896_
timestamp 1644511149
transform 1 0 15548 0 -1 14144
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_2  _2897_
timestamp 1644511149
transform 1 0 16652 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__o21ba_2  _2898_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 35880 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__or3b_1  _2899_
timestamp 1644511149
transform 1 0 36156 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_2  _2900_
timestamp 1644511149
transform 1 0 36432 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__or2_2  _2901_
timestamp 1644511149
transform 1 0 39652 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2902_
timestamp 1644511149
transform 1 0 39100 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _2903_
timestamp 1644511149
transform 1 0 12512 0 -1 14144
box -38 -48 498 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2904_
timestamp 1644511149
transform -1 0 28704 0 -1 13056
box -38 -48 958 592
use sky130_fd_sc_hd__a22o_1  _2905_
timestamp 1644511149
transform -1 0 26036 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a21oi_1  _2906_
timestamp 1644511149
transform 1 0 25300 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_1  _2907_
timestamp 1644511149
transform 1 0 22172 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_2  _2908_
timestamp 1644511149
transform -1 0 12972 0 1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__nand2_1  _2909_
timestamp 1644511149
transform 1 0 12972 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_2  _2910_
timestamp 1644511149
transform 1 0 12236 0 1 13056
box -38 -48 866 592
use sky130_fd_sc_hd__xor2_4  _2911_
timestamp 1644511149
transform 1 0 11592 0 -1 11968
box -38 -48 2062 592
use sky130_fd_sc_hd__buf_4  _2912_
timestamp 1644511149
transform -1 0 36708 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  _2913_
timestamp 1644511149
transform -1 0 21252 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _2914_
timestamp 1644511149
transform 1 0 22724 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _2915_
timestamp 1644511149
transform -1 0 24564 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _2916_
timestamp 1644511149
transform -1 0 23920 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _2917_
timestamp 1644511149
transform -1 0 23368 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_1  _2918_
timestamp 1644511149
transform -1 0 19872 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__xnor2_2  _2919_
timestamp 1644511149
transform -1 0 15272 0 1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_4  _2920_
timestamp 1644511149
transform 1 0 12144 0 -1 9792
box -38 -48 2062 592
use sky130_fd_sc_hd__xnor2_2  _2921_
timestamp 1644511149
transform 1 0 39836 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_4  _2922_
timestamp 1644511149
transform 1 0 40388 0 1 8704
box -38 -48 2062 592
use sky130_fd_sc_hd__xor2_2  _2923_
timestamp 1644511149
transform -1 0 46184 0 1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__xor2_1  _2924_
timestamp 1644511149
transform 1 0 45448 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__o2bb2a_1  _2925_
timestamp 1644511149
transform 1 0 48392 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _2926_
timestamp 1644511149
transform 1 0 48944 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_4  _2927_
timestamp 1644511149
transform -1 0 52256 0 -1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _2928_
timestamp 1644511149
transform 1 0 51704 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _2929_
timestamp 1644511149
transform -1 0 51796 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _2930_
timestamp 1644511149
transform 1 0 9200 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__xnor2_4  _2931_
timestamp 1644511149
transform -1 0 10580 0 -1 14144
box -38 -48 2062 592
use sky130_fd_sc_hd__and2_1  _2932_
timestamp 1644511149
transform -1 0 9384 0 1 35904
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2933_
timestamp 1644511149
transform -1 0 8464 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _2934_
timestamp 1644511149
transform 1 0 8740 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _2935_
timestamp 1644511149
transform 1 0 54096 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_1  _2936_
timestamp 1644511149
transform 1 0 54740 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__nand2_1  _2937_
timestamp 1644511149
transform 1 0 54556 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__a32o_4  _2938_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 56856 0 1 6528
box -38 -48 1602 592
use sky130_fd_sc_hd__xor2_1  _2939_
timestamp 1644511149
transform 1 0 5244 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__or2b_4  _2940_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 48576 0 1 9792
box -38 -48 866 592
use sky130_fd_sc_hd__and2_1  _2941_
timestamp 1644511149
transform 1 0 11960 0 1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2942_
timestamp 1644511149
transform -1 0 12696 0 1 9792
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2943_
timestamp 1644511149
transform -1 0 15272 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _2944_
timestamp 1644511149
transform -1 0 17940 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _2945_
timestamp 1644511149
transform -1 0 17112 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _2946_
timestamp 1644511149
transform 1 0 15180 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__o21ai_2  _2947_
timestamp 1644511149
transform -1 0 12420 0 -1 10880
box -38 -48 682 592
use sky130_fd_sc_hd__or3_1  _2948_
timestamp 1644511149
transform -1 0 13248 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__nand2_1  _2949_
timestamp 1644511149
transform -1 0 11776 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  _2950_
timestamp 1644511149
transform -1 0 18308 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  _2951_
timestamp 1644511149
transform -1 0 30268 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _2952_
timestamp 1644511149
transform 1 0 32108 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__a22o_1  _2953_
timestamp 1644511149
transform 1 0 28152 0 -1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__a221o_2  _2954_
timestamp 1644511149
transform 1 0 29348 0 -1 10880
box -38 -48 866 592
use sky130_fd_sc_hd__xnor2_4  _2955_
timestamp 1644511149
transform -1 0 34132 0 -1 10880
box -38 -48 2062 592
use sky130_fd_sc_hd__xnor2_2  _2956_
timestamp 1644511149
transform -1 0 17572 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__or2_1  _2957_
timestamp 1644511149
transform -1 0 19688 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2958_
timestamp 1644511149
transform 1 0 19228 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  _2959_
timestamp 1644511149
transform -1 0 26588 0 1 9792
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  _2960_
timestamp 1644511149
transform -1 0 26312 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__a22o_1  _2961_
timestamp 1644511149
transform -1 0 24196 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_1  _2962_
timestamp 1644511149
transform 1 0 18676 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_2  _2963_
timestamp 1644511149
transform -1 0 15364 0 1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__xnor2_2  _2964_
timestamp 1644511149
transform -1 0 15272 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__buf_2  _2965_
timestamp 1644511149
transform -1 0 38732 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_1  _2966_
timestamp 1644511149
transform 1 0 11408 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _2967_
timestamp 1644511149
transform 1 0 10212 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2968_
timestamp 1644511149
transform -1 0 11132 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  _2969_
timestamp 1644511149
transform 1 0 37904 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_1  _2970_
timestamp 1644511149
transform -1 0 40388 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o31a_2  _2971_
timestamp 1644511149
transform 1 0 39008 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__xor2_1  _2972_
timestamp 1644511149
transform -1 0 9568 0 1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__xnor2_1  _2973_
timestamp 1644511149
transform 1 0 8924 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__a22oi_4  _2974_ pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform 1 0 44804 0 -1 9792
box -38 -48 1602 592
use sky130_fd_sc_hd__nor2_1  _2975_
timestamp 1644511149
transform -1 0 10212 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _2976_
timestamp 1644511149
transform -1 0 9568 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2977_
timestamp 1644511149
transform -1 0 9384 0 -1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__and2_1  _2978_
timestamp 1644511149
transform 1 0 8004 0 1 11968
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _2979_
timestamp 1644511149
transform 1 0 8280 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  _2980_
timestamp 1644511149
transform -1 0 6808 0 -1 13056
box -38 -48 498 592
use sky130_fd_sc_hd__or2_1  _2981_
timestamp 1644511149
transform 1 0 53636 0 -1 10880
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_2  input1
timestamp 1644511149
transform 1 0 1748 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input2
timestamp 1644511149
transform 1 0 57868 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input3
timestamp 1644511149
transform -1 0 58236 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input4
timestamp 1644511149
transform -1 0 58236 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__buf_4  input5
timestamp 1644511149
transform 1 0 42412 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input6
timestamp 1644511149
transform 1 0 28428 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input7
timestamp 1644511149
transform 1 0 30360 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input8
timestamp 1644511149
transform 1 0 1380 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 1644511149
transform -1 0 58236 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input10
timestamp 1644511149
transform -1 0 57408 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1644511149
transform 1 0 57960 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input12
timestamp 1644511149
transform -1 0 26128 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input13
timestamp 1644511149
transform 1 0 36156 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input14
timestamp 1644511149
transform 1 0 1380 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1644511149
transform -1 0 8096 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  input16
timestamp 1644511149
transform -1 0 58236 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input17
timestamp 1644511149
transform 1 0 24380 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input18
timestamp 1644511149
transform 1 0 1748 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input19
timestamp 1644511149
transform 1 0 1748 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  input20 pdk5/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1644511149
transform -1 0 58236 0 1 7616
box -38 -48 866 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input21
timestamp 1644511149
transform 1 0 9752 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_4  input22
timestamp 1644511149
transform -1 0 58236 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input23
timestamp 1644511149
transform -1 0 58236 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input24
timestamp 1644511149
transform 1 0 1748 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input25
timestamp 1644511149
transform 1 0 19964 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input26
timestamp 1644511149
transform -1 0 58236 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input27
timestamp 1644511149
transform -1 0 31648 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input28
timestamp 1644511149
transform -1 0 56488 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input29
timestamp 1644511149
transform -1 0 58236 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1644511149
transform -1 0 41952 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1644511149
transform -1 0 34224 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input32
timestamp 1644511149
transform 1 0 9752 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input33
timestamp 1644511149
transform -1 0 58236 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  input34
timestamp 1644511149
transform 1 0 20056 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_2  input35
timestamp 1644511149
transform 1 0 1748 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input36
timestamp 1644511149
transform 1 0 24748 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  input37
timestamp 1644511149
transform 1 0 1380 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  input38
timestamp 1644511149
transform 1 0 29900 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1644511149
transform -1 0 1656 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  input40
timestamp 1644511149
transform 1 0 37628 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input41
timestamp 1644511149
transform 1 0 1748 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input42
timestamp 1644511149
transform -1 0 12696 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input43
timestamp 1644511149
transform 1 0 1748 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input44
timestamp 1644511149
transform 1 0 2576 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_6  input45
timestamp 1644511149
transform 1 0 56120 0 1 36992
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_4  input46
timestamp 1644511149
transform -1 0 48484 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  input47
timestamp 1644511149
transform 1 0 21988 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input48
timestamp 1644511149
transform -1 0 58236 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__buf_6  input49
timestamp 1644511149
transform -1 0 54832 0 1 2176
box -38 -48 866 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1644511149
transform -1 0 1656 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1644511149
transform -1 0 1656 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input52
timestamp 1644511149
transform -1 0 8464 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input53
timestamp 1644511149
transform 1 0 15272 0 1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input54
timestamp 1644511149
transform 1 0 26956 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input55
timestamp 1644511149
transform -1 0 58236 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input56
timestamp 1644511149
transform 1 0 27784 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input57
timestamp 1644511149
transform 1 0 50508 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input58
timestamp 1644511149
transform 1 0 48852 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input59
timestamp 1644511149
transform 1 0 14260 0 1 36992
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input60
timestamp 1644511149
transform -1 0 22540 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input61
timestamp 1644511149
transform 1 0 34684 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input62
timestamp 1644511149
transform -1 0 1656 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input63
timestamp 1644511149
transform 1 0 4140 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_4  input64
timestamp 1644511149
transform -1 0 58236 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output65
timestamp 1644511149
transform 1 0 52716 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output66
timestamp 1644511149
transform -1 0 12052 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output67
timestamp 1644511149
transform -1 0 50692 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output68
timestamp 1644511149
transform -1 0 46184 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output69
timestamp 1644511149
transform -1 0 32660 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output70
timestamp 1644511149
transform -1 0 40204 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output71
timestamp 1644511149
transform 1 0 54188 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output72
timestamp 1644511149
transform -1 0 48116 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output73
timestamp 1644511149
transform 1 0 57868 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output74
timestamp 1644511149
transform -1 0 1748 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output75
timestamp 1644511149
transform -1 0 40940 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output76
timestamp 1644511149
transform -1 0 18492 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output77
timestamp 1644511149
transform 1 0 57868 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output78
timestamp 1644511149
transform 1 0 57868 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output79
timestamp 1644511149
transform 1 0 6348 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output80
timestamp 1644511149
transform -1 0 1748 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output81
timestamp 1644511149
transform -1 0 1748 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output82
timestamp 1644511149
transform 1 0 38088 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output83
timestamp 1644511149
transform -1 0 2484 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output84
timestamp 1644511149
transform 1 0 16652 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output85
timestamp 1644511149
transform -1 0 4324 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output86
timestamp 1644511149
transform 1 0 14076 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1644511149
transform 1 0 43884 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1644511149
transform 1 0 57868 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output89
timestamp 1644511149
transform 1 0 57868 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1644511149
transform -1 0 1748 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1644511149
transform -1 0 1748 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output92
timestamp 1644511149
transform 1 0 52716 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output93
timestamp 1644511149
transform -1 0 18492 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output94
timestamp 1644511149
transform 1 0 57868 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output95
timestamp 1644511149
transform -1 0 1748 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1644511149
transform -1 0 41124 0 1 2176
box -38 -48 406 592
<< labels >>
rlabel metal2 s 5814 0 5870 800 6 CLK
port 0 nsew signal input
rlabel metal2 s 44454 39200 44510 40000 6 RST
port 1 nsew signal input
rlabel metal3 s 0 23128 800 23248 6 az[0]
port 2 nsew signal input
rlabel metal2 s 57978 39200 58034 40000 6 az[10]
port 3 nsew signal input
rlabel metal3 s 59200 31288 60000 31408 6 az[11]
port 4 nsew signal input
rlabel metal3 s 59200 20408 60000 20528 6 az[12]
port 5 nsew signal input
rlabel metal2 s 41878 0 41934 800 6 az[13]
port 6 nsew signal input
rlabel metal2 s 28354 39200 28410 40000 6 az[14]
port 7 nsew signal input
rlabel metal2 s 30286 39200 30342 40000 6 az[15]
port 8 nsew signal input
rlabel metal3 s 0 19048 800 19168 6 az[16]
port 9 nsew signal input
rlabel metal3 s 59200 37408 60000 37528 6 az[17]
port 10 nsew signal input
rlabel metal3 s 59200 1368 60000 1488 6 az[18]
port 11 nsew signal input
rlabel metal3 s 59200 29248 60000 29368 6 az[19]
port 12 nsew signal input
rlabel metal2 s 25778 39200 25834 40000 6 az[1]
port 13 nsew signal input
rlabel metal2 s 36082 0 36138 800 6 az[20]
port 14 nsew signal input
rlabel metal3 s 0 2048 800 2168 6 az[21]
port 15 nsew signal input
rlabel metal2 s 7746 39200 7802 40000 6 az[22]
port 16 nsew signal input
rlabel metal3 s 59200 35368 60000 35488 6 az[23]
port 17 nsew signal input
rlabel metal2 s 23846 39200 23902 40000 6 az[24]
port 18 nsew signal input
rlabel metal3 s 0 25168 800 25288 6 az[25]
port 19 nsew signal input
rlabel metal3 s 0 33328 800 33448 6 az[26]
port 20 nsew signal input
rlabel metal3 s 59200 8168 60000 8288 6 az[27]
port 21 nsew signal input
rlabel metal2 s 9678 0 9734 800 6 az[28]
port 22 nsew signal input
rlabel metal3 s 59200 16328 60000 16448 6 az[29]
port 23 nsew signal input
rlabel metal3 s 59200 3408 60000 3528 6 az[2]
port 24 nsew signal input
rlabel metal3 s 0 6128 800 6248 6 az[30]
port 25 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 az[31]
port 26 nsew signal input
rlabel metal3 s 59200 27208 60000 27328 6 az[3]
port 27 nsew signal input
rlabel metal2 s 31574 0 31630 800 6 az[4]
port 28 nsew signal input
rlabel metal2 s 56046 0 56102 800 6 az[5]
port 29 nsew signal input
rlabel metal3 s 59200 33328 60000 33448 6 az[6]
port 30 nsew signal input
rlabel metal2 s 41878 39200 41934 40000 6 az[7]
port 31 nsew signal input
rlabel metal2 s 34150 39200 34206 40000 6 az[8]
port 32 nsew signal input
rlabel metal2 s 9678 39200 9734 40000 6 az[9]
port 33 nsew signal input
rlabel metal2 s 52182 39200 52238 40000 6 mac[0]
port 34 nsew signal tristate
rlabel metal2 s 11610 0 11666 800 6 mac[10]
port 35 nsew signal tristate
rlabel metal2 s 50250 0 50306 800 6 mac[11]
port 36 nsew signal tristate
rlabel metal2 s 45742 0 45798 800 6 mac[12]
port 37 nsew signal tristate
rlabel metal2 s 32218 39200 32274 40000 6 mac[13]
port 38 nsew signal tristate
rlabel metal2 s 38014 39200 38070 40000 6 mac[14]
port 39 nsew signal tristate
rlabel metal2 s 54114 39200 54170 40000 6 mac[15]
port 40 nsew signal tristate
rlabel metal2 s 47674 0 47730 800 6 mac[16]
port 41 nsew signal tristate
rlabel metal3 s 59200 25168 60000 25288 6 mac[17]
port 42 nsew signal tristate
rlabel metal3 s 0 36048 800 36168 6 mac[18]
port 43 nsew signal tristate
rlabel metal2 s 39946 39200 40002 40000 6 mac[19]
port 44 nsew signal tristate
rlabel metal2 s 18050 0 18106 800 6 mac[1]
port 45 nsew signal tristate
rlabel metal2 s 57978 0 58034 800 6 mac[20]
port 46 nsew signal tristate
rlabel metal3 s 59200 14288 60000 14408 6 mac[21]
port 47 nsew signal tristate
rlabel metal2 s 5814 39200 5870 40000 6 mac[22]
port 48 nsew signal tristate
rlabel metal2 s 18 39200 74 40000 6 mac[23]
port 49 nsew signal tristate
rlabel metal3 s 0 38088 800 38208 6 mac[24]
port 50 nsew signal tristate
rlabel metal2 s 38014 0 38070 800 6 mac[25]
port 51 nsew signal tristate
rlabel metal2 s 1950 39200 2006 40000 6 mac[26]
port 52 nsew signal tristate
rlabel metal2 s 16118 39200 16174 40000 6 mac[27]
port 53 nsew signal tristate
rlabel metal2 s 3882 0 3938 800 6 mac[28]
port 54 nsew signal tristate
rlabel metal2 s 13542 0 13598 800 6 mac[29]
port 55 nsew signal tristate
rlabel metal2 s 43810 0 43866 800 6 mac[2]
port 56 nsew signal tristate
rlabel metal3 s 59200 10208 60000 10328 6 mac[30]
port 57 nsew signal tristate
rlabel metal2 s 59910 0 59966 800 6 mac[31]
port 58 nsew signal tristate
rlabel metal3 s 0 8168 800 8288 6 mac[3]
port 59 nsew signal tristate
rlabel metal3 s 0 4088 800 4208 6 mac[4]
port 60 nsew signal tristate
rlabel metal2 s 52182 0 52238 800 6 mac[5]
port 61 nsew signal tristate
rlabel metal2 s 18050 39200 18106 40000 6 mac[6]
port 62 nsew signal tristate
rlabel metal3 s 59200 6128 60000 6248 6 mac[7]
port 63 nsew signal tristate
rlabel metal3 s 0 29248 800 29368 6 mac[8]
port 64 nsew signal tristate
rlabel metal2 s 39946 0 40002 800 6 mac[9]
port 65 nsew signal tristate
rlabel metal3 s 59200 23128 60000 23248 6 mx[0]
port 66 nsew signal input
rlabel metal2 s 19982 39200 20038 40000 6 mx[10]
port 67 nsew signal input
rlabel metal3 s 0 31288 800 31408 6 mx[11]
port 68 nsew signal input
rlabel metal2 s 23846 0 23902 800 6 mx[12]
port 69 nsew signal input
rlabel metal2 s 18 0 74 800 6 mx[13]
port 70 nsew signal input
rlabel metal2 s 29642 0 29698 800 6 mx[14]
port 71 nsew signal input
rlabel metal3 s 0 10208 800 10328 6 mx[15]
port 72 nsew signal input
rlabel metal2 s 36082 39200 36138 40000 6 mx[1]
port 73 nsew signal input
rlabel metal3 s 0 16328 800 16448 6 mx[2]
port 74 nsew signal input
rlabel metal2 s 12254 39200 12310 40000 6 mx[3]
port 75 nsew signal input
rlabel metal3 s 0 27208 800 27328 6 mx[4]
port 76 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 mx[5]
port 77 nsew signal input
rlabel metal2 s 56046 39200 56102 40000 6 mx[6]
port 78 nsew signal input
rlabel metal2 s 46386 39200 46442 40000 6 mx[7]
port 79 nsew signal input
rlabel metal2 s 21914 0 21970 800 6 mx[8]
port 80 nsew signal input
rlabel metal2 s 59910 39200 59966 40000 6 mx[9]
port 81 nsew signal input
rlabel metal2 s 54114 0 54170 800 6 my[0]
port 82 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 my[10]
port 83 nsew signal input
rlabel metal3 s 0 21088 800 21208 6 my[11]
port 84 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 my[12]
port 85 nsew signal input
rlabel metal2 s 15474 0 15530 800 6 my[13]
port 86 nsew signal input
rlabel metal2 s 25778 0 25834 800 6 my[14]
port 87 nsew signal input
rlabel metal3 s 59200 18368 60000 18488 6 my[15]
port 88 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 my[1]
port 89 nsew signal input
rlabel metal2 s 50250 39200 50306 40000 6 my[2]
port 90 nsew signal input
rlabel metal2 s 48318 39200 48374 40000 6 my[3]
port 91 nsew signal input
rlabel metal2 s 14186 39200 14242 40000 6 my[4]
port 92 nsew signal input
rlabel metal2 s 21914 39200 21970 40000 6 my[5]
port 93 nsew signal input
rlabel metal2 s 34150 0 34206 800 6 my[6]
port 94 nsew signal input
rlabel metal3 s 0 14288 800 14408 6 my[7]
port 95 nsew signal input
rlabel metal2 s 3882 39200 3938 40000 6 my[8]
port 96 nsew signal input
rlabel metal3 s 59200 12248 60000 12368 6 my[9]
port 97 nsew signal input
rlabel metal4 s 4208 2128 4528 37584 6 vccd1
port 98 nsew power input
rlabel metal4 s 34928 2128 35248 37584 6 vccd1
port 98 nsew power input
rlabel metal4 s 19568 2128 19888 37584 6 vssd1
port 99 nsew ground input
rlabel metal4 s 50288 2128 50608 37584 6 vssd1
port 99 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 60000 40000
<< end >>
