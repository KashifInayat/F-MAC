magic
tech sky130A
magscale 1 2
timestamp 1647889168
<< obsli1 >>
rect 1104 2159 58880 37553
<< obsm1 >>
rect 14 1708 59970 37664
<< metal2 >>
rect 18 39200 74 40000
rect 1950 39200 2006 40000
rect 3882 39200 3938 40000
rect 5814 39200 5870 40000
rect 7746 39200 7802 40000
rect 9678 39200 9734 40000
rect 12254 39200 12310 40000
rect 14186 39200 14242 40000
rect 16118 39200 16174 40000
rect 18050 39200 18106 40000
rect 19982 39200 20038 40000
rect 21914 39200 21970 40000
rect 23846 39200 23902 40000
rect 25778 39200 25834 40000
rect 28354 39200 28410 40000
rect 30286 39200 30342 40000
rect 32218 39200 32274 40000
rect 34150 39200 34206 40000
rect 36082 39200 36138 40000
rect 38014 39200 38070 40000
rect 39946 39200 40002 40000
rect 41878 39200 41934 40000
rect 44454 39200 44510 40000
rect 46386 39200 46442 40000
rect 48318 39200 48374 40000
rect 50250 39200 50306 40000
rect 52182 39200 52238 40000
rect 54114 39200 54170 40000
rect 56046 39200 56102 40000
rect 57978 39200 58034 40000
rect 59910 39200 59966 40000
rect 18 0 74 800
rect 1950 0 2006 800
rect 3882 0 3938 800
rect 5814 0 5870 800
rect 7746 0 7802 800
rect 9678 0 9734 800
rect 11610 0 11666 800
rect 13542 0 13598 800
rect 15474 0 15530 800
rect 18050 0 18106 800
rect 19982 0 20038 800
rect 21914 0 21970 800
rect 23846 0 23902 800
rect 25778 0 25834 800
rect 27710 0 27766 800
rect 29642 0 29698 800
rect 31574 0 31630 800
rect 34150 0 34206 800
rect 36082 0 36138 800
rect 38014 0 38070 800
rect 39946 0 40002 800
rect 41878 0 41934 800
rect 43810 0 43866 800
rect 45742 0 45798 800
rect 47674 0 47730 800
rect 50250 0 50306 800
rect 52182 0 52238 800
rect 54114 0 54170 800
rect 56046 0 56102 800
rect 57978 0 58034 800
rect 59910 0 59966 800
<< obsm2 >>
rect 130 39144 1894 39250
rect 2062 39144 3826 39250
rect 3994 39144 5758 39250
rect 5926 39144 7690 39250
rect 7858 39144 9622 39250
rect 9790 39144 12198 39250
rect 12366 39144 14130 39250
rect 14298 39144 16062 39250
rect 16230 39144 17994 39250
rect 18162 39144 19926 39250
rect 20094 39144 21858 39250
rect 22026 39144 23790 39250
rect 23958 39144 25722 39250
rect 25890 39144 28298 39250
rect 28466 39144 30230 39250
rect 30398 39144 32162 39250
rect 32330 39144 34094 39250
rect 34262 39144 36026 39250
rect 36194 39144 37958 39250
rect 38126 39144 39890 39250
rect 40058 39144 41822 39250
rect 41990 39144 44398 39250
rect 44566 39144 46330 39250
rect 46498 39144 48262 39250
rect 48430 39144 50194 39250
rect 50362 39144 52126 39250
rect 52294 39144 54058 39250
rect 54226 39144 55990 39250
rect 56158 39144 57922 39250
rect 58090 39144 59854 39250
rect 20 856 59964 39144
rect 130 734 1894 856
rect 2062 734 3826 856
rect 3994 734 5758 856
rect 5926 734 7690 856
rect 7858 734 9622 856
rect 9790 734 11554 856
rect 11722 734 13486 856
rect 13654 734 15418 856
rect 15586 734 17994 856
rect 18162 734 19926 856
rect 20094 734 21858 856
rect 22026 734 23790 856
rect 23958 734 25722 856
rect 25890 734 27654 856
rect 27822 734 29586 856
rect 29754 734 31518 856
rect 31686 734 34094 856
rect 34262 734 36026 856
rect 36194 734 37958 856
rect 38126 734 39890 856
rect 40058 734 41822 856
rect 41990 734 43754 856
rect 43922 734 45686 856
rect 45854 734 47618 856
rect 47786 734 50194 856
rect 50362 734 52126 856
rect 52294 734 54058 856
rect 54226 734 55990 856
rect 56158 734 57922 856
rect 58090 734 59854 856
<< metal3 >>
rect 0 38088 800 38208
rect 59200 37408 60000 37528
rect 0 36048 800 36168
rect 59200 35368 60000 35488
rect 0 33328 800 33448
rect 59200 33328 60000 33448
rect 0 31288 800 31408
rect 59200 31288 60000 31408
rect 0 29248 800 29368
rect 59200 29248 60000 29368
rect 0 27208 800 27328
rect 59200 27208 60000 27328
rect 0 25168 800 25288
rect 59200 25168 60000 25288
rect 0 23128 800 23248
rect 59200 23128 60000 23248
rect 0 21088 800 21208
rect 59200 20408 60000 20528
rect 0 19048 800 19168
rect 59200 18368 60000 18488
rect 0 16328 800 16448
rect 59200 16328 60000 16448
rect 0 14288 800 14408
rect 59200 14288 60000 14408
rect 0 12248 800 12368
rect 59200 12248 60000 12368
rect 0 10208 800 10328
rect 59200 10208 60000 10328
rect 0 8168 800 8288
rect 59200 8168 60000 8288
rect 0 6128 800 6248
rect 59200 6128 60000 6248
rect 0 4088 800 4208
rect 59200 3408 60000 3528
rect 0 2048 800 2168
rect 59200 1368 60000 1488
<< obsm3 >>
rect 880 38008 59200 38181
rect 800 37608 59200 38008
rect 800 37328 59120 37608
rect 800 36248 59200 37328
rect 880 35968 59200 36248
rect 800 35568 59200 35968
rect 800 35288 59120 35568
rect 800 33528 59200 35288
rect 880 33248 59120 33528
rect 800 31488 59200 33248
rect 880 31208 59120 31488
rect 800 29448 59200 31208
rect 880 29168 59120 29448
rect 800 27408 59200 29168
rect 880 27128 59120 27408
rect 800 25368 59200 27128
rect 880 25088 59120 25368
rect 800 23328 59200 25088
rect 880 23048 59120 23328
rect 800 21288 59200 23048
rect 880 21008 59200 21288
rect 800 20608 59200 21008
rect 800 20328 59120 20608
rect 800 19248 59200 20328
rect 880 18968 59200 19248
rect 800 18568 59200 18968
rect 800 18288 59120 18568
rect 800 16528 59200 18288
rect 880 16248 59120 16528
rect 800 14488 59200 16248
rect 880 14208 59120 14488
rect 800 12448 59200 14208
rect 880 12168 59120 12448
rect 800 10408 59200 12168
rect 880 10128 59120 10408
rect 800 8368 59200 10128
rect 880 8088 59120 8368
rect 800 6328 59200 8088
rect 880 6048 59120 6328
rect 800 4288 59200 6048
rect 880 4008 59200 4288
rect 800 3608 59200 4008
rect 800 3328 59120 3608
rect 800 2248 59200 3328
rect 880 1968 59200 2248
rect 800 1568 59200 1968
rect 800 1395 59120 1568
<< metal4 >>
rect 4208 2128 4528 37584
rect 19568 2128 19888 37584
rect 34928 2128 35248 37584
rect 50288 2128 50608 37584
<< obsm4 >>
rect 21219 15267 23677 26621
<< labels >>
rlabel metal2 s 5814 0 5870 800 6 CLK
port 1 nsew signal input
rlabel metal2 s 44454 39200 44510 40000 6 RST
port 2 nsew signal input
rlabel metal3 s 0 23128 800 23248 6 az[0]
port 3 nsew signal input
rlabel metal2 s 57978 39200 58034 40000 6 az[10]
port 4 nsew signal input
rlabel metal3 s 59200 31288 60000 31408 6 az[11]
port 5 nsew signal input
rlabel metal3 s 59200 20408 60000 20528 6 az[12]
port 6 nsew signal input
rlabel metal2 s 41878 0 41934 800 6 az[13]
port 7 nsew signal input
rlabel metal2 s 28354 39200 28410 40000 6 az[14]
port 8 nsew signal input
rlabel metal2 s 30286 39200 30342 40000 6 az[15]
port 9 nsew signal input
rlabel metal3 s 0 19048 800 19168 6 az[16]
port 10 nsew signal input
rlabel metal3 s 59200 37408 60000 37528 6 az[17]
port 11 nsew signal input
rlabel metal3 s 59200 1368 60000 1488 6 az[18]
port 12 nsew signal input
rlabel metal3 s 59200 29248 60000 29368 6 az[19]
port 13 nsew signal input
rlabel metal2 s 25778 39200 25834 40000 6 az[1]
port 14 nsew signal input
rlabel metal2 s 36082 0 36138 800 6 az[20]
port 15 nsew signal input
rlabel metal3 s 0 2048 800 2168 6 az[21]
port 16 nsew signal input
rlabel metal2 s 7746 39200 7802 40000 6 az[22]
port 17 nsew signal input
rlabel metal3 s 59200 35368 60000 35488 6 az[23]
port 18 nsew signal input
rlabel metal2 s 23846 39200 23902 40000 6 az[24]
port 19 nsew signal input
rlabel metal3 s 0 25168 800 25288 6 az[25]
port 20 nsew signal input
rlabel metal3 s 0 33328 800 33448 6 az[26]
port 21 nsew signal input
rlabel metal3 s 59200 8168 60000 8288 6 az[27]
port 22 nsew signal input
rlabel metal2 s 9678 0 9734 800 6 az[28]
port 23 nsew signal input
rlabel metal3 s 59200 16328 60000 16448 6 az[29]
port 24 nsew signal input
rlabel metal3 s 59200 3408 60000 3528 6 az[2]
port 25 nsew signal input
rlabel metal3 s 0 6128 800 6248 6 az[30]
port 26 nsew signal input
rlabel metal2 s 19982 0 20038 800 6 az[31]
port 27 nsew signal input
rlabel metal3 s 59200 27208 60000 27328 6 az[3]
port 28 nsew signal input
rlabel metal2 s 31574 0 31630 800 6 az[4]
port 29 nsew signal input
rlabel metal2 s 56046 0 56102 800 6 az[5]
port 30 nsew signal input
rlabel metal3 s 59200 33328 60000 33448 6 az[6]
port 31 nsew signal input
rlabel metal2 s 41878 39200 41934 40000 6 az[7]
port 32 nsew signal input
rlabel metal2 s 34150 39200 34206 40000 6 az[8]
port 33 nsew signal input
rlabel metal2 s 9678 39200 9734 40000 6 az[9]
port 34 nsew signal input
rlabel metal2 s 52182 39200 52238 40000 6 mac[0]
port 35 nsew signal output
rlabel metal2 s 11610 0 11666 800 6 mac[10]
port 36 nsew signal output
rlabel metal2 s 50250 0 50306 800 6 mac[11]
port 37 nsew signal output
rlabel metal2 s 45742 0 45798 800 6 mac[12]
port 38 nsew signal output
rlabel metal2 s 32218 39200 32274 40000 6 mac[13]
port 39 nsew signal output
rlabel metal2 s 38014 39200 38070 40000 6 mac[14]
port 40 nsew signal output
rlabel metal2 s 54114 39200 54170 40000 6 mac[15]
port 41 nsew signal output
rlabel metal2 s 47674 0 47730 800 6 mac[16]
port 42 nsew signal output
rlabel metal3 s 59200 25168 60000 25288 6 mac[17]
port 43 nsew signal output
rlabel metal3 s 0 36048 800 36168 6 mac[18]
port 44 nsew signal output
rlabel metal2 s 39946 39200 40002 40000 6 mac[19]
port 45 nsew signal output
rlabel metal2 s 18050 0 18106 800 6 mac[1]
port 46 nsew signal output
rlabel metal2 s 57978 0 58034 800 6 mac[20]
port 47 nsew signal output
rlabel metal3 s 59200 14288 60000 14408 6 mac[21]
port 48 nsew signal output
rlabel metal2 s 5814 39200 5870 40000 6 mac[22]
port 49 nsew signal output
rlabel metal2 s 18 39200 74 40000 6 mac[23]
port 50 nsew signal output
rlabel metal3 s 0 38088 800 38208 6 mac[24]
port 51 nsew signal output
rlabel metal2 s 38014 0 38070 800 6 mac[25]
port 52 nsew signal output
rlabel metal2 s 1950 39200 2006 40000 6 mac[26]
port 53 nsew signal output
rlabel metal2 s 16118 39200 16174 40000 6 mac[27]
port 54 nsew signal output
rlabel metal2 s 3882 0 3938 800 6 mac[28]
port 55 nsew signal output
rlabel metal2 s 13542 0 13598 800 6 mac[29]
port 56 nsew signal output
rlabel metal2 s 43810 0 43866 800 6 mac[2]
port 57 nsew signal output
rlabel metal3 s 59200 10208 60000 10328 6 mac[30]
port 58 nsew signal output
rlabel metal2 s 59910 0 59966 800 6 mac[31]
port 59 nsew signal output
rlabel metal3 s 0 8168 800 8288 6 mac[3]
port 60 nsew signal output
rlabel metal3 s 0 4088 800 4208 6 mac[4]
port 61 nsew signal output
rlabel metal2 s 52182 0 52238 800 6 mac[5]
port 62 nsew signal output
rlabel metal2 s 18050 39200 18106 40000 6 mac[6]
port 63 nsew signal output
rlabel metal3 s 59200 6128 60000 6248 6 mac[7]
port 64 nsew signal output
rlabel metal3 s 0 29248 800 29368 6 mac[8]
port 65 nsew signal output
rlabel metal2 s 39946 0 40002 800 6 mac[9]
port 66 nsew signal output
rlabel metal3 s 59200 23128 60000 23248 6 mx[0]
port 67 nsew signal input
rlabel metal2 s 19982 39200 20038 40000 6 mx[10]
port 68 nsew signal input
rlabel metal3 s 0 31288 800 31408 6 mx[11]
port 69 nsew signal input
rlabel metal2 s 23846 0 23902 800 6 mx[12]
port 70 nsew signal input
rlabel metal2 s 18 0 74 800 6 mx[13]
port 71 nsew signal input
rlabel metal2 s 29642 0 29698 800 6 mx[14]
port 72 nsew signal input
rlabel metal3 s 0 10208 800 10328 6 mx[15]
port 73 nsew signal input
rlabel metal2 s 36082 39200 36138 40000 6 mx[1]
port 74 nsew signal input
rlabel metal3 s 0 16328 800 16448 6 mx[2]
port 75 nsew signal input
rlabel metal2 s 12254 39200 12310 40000 6 mx[3]
port 76 nsew signal input
rlabel metal3 s 0 27208 800 27328 6 mx[4]
port 77 nsew signal input
rlabel metal2 s 1950 0 2006 800 6 mx[5]
port 78 nsew signal input
rlabel metal2 s 56046 39200 56102 40000 6 mx[6]
port 79 nsew signal input
rlabel metal2 s 46386 39200 46442 40000 6 mx[7]
port 80 nsew signal input
rlabel metal2 s 21914 0 21970 800 6 mx[8]
port 81 nsew signal input
rlabel metal2 s 59910 39200 59966 40000 6 mx[9]
port 82 nsew signal input
rlabel metal2 s 54114 0 54170 800 6 my[0]
port 83 nsew signal input
rlabel metal3 s 0 12248 800 12368 6 my[10]
port 84 nsew signal input
rlabel metal3 s 0 21088 800 21208 6 my[11]
port 85 nsew signal input
rlabel metal2 s 7746 0 7802 800 6 my[12]
port 86 nsew signal input
rlabel metal2 s 15474 0 15530 800 6 my[13]
port 87 nsew signal input
rlabel metal2 s 25778 0 25834 800 6 my[14]
port 88 nsew signal input
rlabel metal3 s 59200 18368 60000 18488 6 my[15]
port 89 nsew signal input
rlabel metal2 s 27710 0 27766 800 6 my[1]
port 90 nsew signal input
rlabel metal2 s 50250 39200 50306 40000 6 my[2]
port 91 nsew signal input
rlabel metal2 s 48318 39200 48374 40000 6 my[3]
port 92 nsew signal input
rlabel metal2 s 14186 39200 14242 40000 6 my[4]
port 93 nsew signal input
rlabel metal2 s 21914 39200 21970 40000 6 my[5]
port 94 nsew signal input
rlabel metal2 s 34150 0 34206 800 6 my[6]
port 95 nsew signal input
rlabel metal3 s 0 14288 800 14408 6 my[7]
port 96 nsew signal input
rlabel metal2 s 3882 39200 3938 40000 6 my[8]
port 97 nsew signal input
rlabel metal3 s 59200 12248 60000 12368 6 my[9]
port 98 nsew signal input
rlabel metal4 s 4208 2128 4528 37584 6 vccd1
port 99 nsew power input
rlabel metal4 s 34928 2128 35248 37584 6 vccd1
port 99 nsew power input
rlabel metal4 s 19568 2128 19888 37584 6 vssd1
port 100 nsew ground input
rlabel metal4 s 50288 2128 50608 37584 6 vssd1
port 100 nsew ground input
<< properties >>
string FIXED_BBOX 0 0 60000 40000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 5091264
string GDS_FILE /home/engrkashif/work/mpw5/caravel_user_project/openlane/mac_top/runs/mac_top/results/finishing/mac_top.magic.gds
string GDS_START 803600
<< end >>

