* NGSPICE file created from user_proj_example.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_1 abstract view
.subckt sky130_fd_sc_hd__nor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_2 abstract view
.subckt sky130_fd_sc_hd__clkbuf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_2 abstract view
.subckt sky130_fd_sc_hd__xnor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_1 abstract view
.subckt sky130_fd_sc_hd__a21o_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_2 abstract view
.subckt sky130_fd_sc_hd__o211ai_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_2 abstract view
.subckt sky130_fd_sc_hd__a21oi_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_1 abstract view
.subckt sky130_fd_sc_hd__xnor2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_1 abstract view
.subckt sky130_fd_sc_hd__a31o_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_1 abstract view
.subckt sky130_fd_sc_hd__a22o_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_1 abstract view
.subckt sky130_fd_sc_hd__xor2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_1 abstract view
.subckt sky130_fd_sc_hd__or3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_1 abstract view
.subckt sky130_fd_sc_hd__and3_1 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_1 abstract view
.subckt sky130_fd_sc_hd__or2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_1 abstract view
.subckt sky130_fd_sc_hd__a21oi_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_1 abstract view
.subckt sky130_fd_sc_hd__a221o_1 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22o_2 abstract view
.subckt sky130_fd_sc_hd__a22o_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3b_1 abstract view
.subckt sky130_fd_sc_hd__or3b_1 A B C_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor2_2 abstract view
.subckt sky130_fd_sc_hd__nor2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21bo_1 abstract view
.subckt sky130_fd_sc_hd__a21bo_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_1 abstract view
.subckt sky130_fd_sc_hd__a211o_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_1 abstract view
.subckt sky130_fd_sc_hd__o21a_1 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_1 abstract view
.subckt sky130_fd_sc_hd__o21bai_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_2 abstract view
.subckt sky130_fd_sc_hd__and3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_1 abstract view
.subckt sky130_fd_sc_hd__or2b_1 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xnor2_4 abstract view
.subckt sky130_fd_sc_hd__xnor2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_2 abstract view
.subckt sky130_fd_sc_hd__xor2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_1 abstract view
.subckt sky130_fd_sc_hd__nand2_1 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_2 abstract view
.subckt sky130_fd_sc_hd__a211o_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_2 abstract view
.subckt sky130_fd_sc_hd__nand3b_2 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dlymetal6s2s_1 abstract view
.subckt sky130_fd_sc_hd__dlymetal6s2s_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_1 abstract view
.subckt sky130_fd_sc_hd__a211oi_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_2 abstract view
.subckt sky130_fd_sc_hd__and2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_1 abstract view
.subckt sky130_fd_sc_hd__o21ba_1 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_1 abstract view
.subckt sky130_fd_sc_hd__nand3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_1 abstract view
.subckt sky130_fd_sc_hd__nor3_1 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_1 abstract view
.subckt sky130_fd_sc_hd__o211a_1 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_2 abstract view
.subckt sky130_fd_sc_hd__or2_2 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_1 abstract view
.subckt sky130_fd_sc_hd__o21ai_1 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3b_1 abstract view
.subckt sky130_fd_sc_hd__and3b_1 A_N B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22ai_4 abstract view
.subckt sky130_fd_sc_hd__o22ai_4 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2bb2o_1 abstract view
.subckt sky130_fd_sc_hd__a2bb2o_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_4 abstract view
.subckt sky130_fd_sc_hd__o21ai_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221oi_4 abstract view
.subckt sky130_fd_sc_hd__a221oi_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_4 abstract view
.subckt sky130_fd_sc_hd__nand4_4 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_1 abstract view
.subckt sky130_fd_sc_hd__a22oi_1 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2b_2 abstract view
.subckt sky130_fd_sc_hd__or2b_2 A B_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a31o_2 abstract view
.subckt sky130_fd_sc_hd__a31o_2 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21o_2 abstract view
.subckt sky130_fd_sc_hd__a21o_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_2 abstract view
.subckt sky130_fd_sc_hd__a221o_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21oi_4 abstract view
.subckt sky130_fd_sc_hd__a21oi_4 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_2 abstract view
.subckt sky130_fd_sc_hd__or3_2 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_1 abstract view
.subckt sky130_fd_sc_hd__a311o_1 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o2bb2a_1 abstract view
.subckt sky130_fd_sc_hd__o2bb2a_1 A1_N A2_N B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_2 abstract view
.subckt sky130_fd_sc_hd__o31ai_2 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_2 abstract view
.subckt sky130_fd_sc_hd__nand3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_2 abstract view
.subckt sky130_fd_sc_hd__nand2_2 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_1 abstract view
.subckt sky130_fd_sc_hd__mux2_1 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_8 abstract view
.subckt sky130_fd_sc_hd__clkbuf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_4 abstract view
.subckt sky130_fd_sc_hd__a21boi_4 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_1 abstract view
.subckt sky130_fd_sc_hd__or4_1 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__xor2_4 abstract view
.subckt sky130_fd_sc_hd__xor2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_6 abstract view
.subckt sky130_fd_sc_hd__buf_6 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ai_2 abstract view
.subckt sky130_fd_sc_hd__o21ai_2 A1 A2 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a311o_4 abstract view
.subckt sky130_fd_sc_hd__a311o_4 A1 A2 A3 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3b_1 abstract view
.subckt sky130_fd_sc_hd__nand3b_1 A_N B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4_4 abstract view
.subckt sky130_fd_sc_hd__or4_4 A B C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21a_2 abstract view
.subckt sky130_fd_sc_hd__o21a_2 A1 A2 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_1 abstract view
.subckt sky130_fd_sc_hd__o211ai_1 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_4 abstract view
.subckt sky130_fd_sc_hd__buf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21bai_2 abstract view
.subckt sky130_fd_sc_hd__o21bai_2 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a21boi_1 abstract view
.subckt sky130_fd_sc_hd__a21boi_1 A1 A2 B1_N VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a221o_4 abstract view
.subckt sky130_fd_sc_hd__a221o_4 A1 A2 B1 B2 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_1 abstract view
.subckt sky130_fd_sc_hd__a32o_1 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31ai_4 abstract view
.subckt sky130_fd_sc_hd__o31ai_4 A1 A2 A3 B1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o31a_1 abstract view
.subckt sky130_fd_sc_hd__o31a_1 A1 A2 A3 B1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__mux2_2 abstract view
.subckt sky130_fd_sc_hd__mux2_2 A0 A1 S VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_2 abstract view
.subckt sky130_fd_sc_hd__a211oi_2 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nor3_2 abstract view
.subckt sky130_fd_sc_hd__nor3_2 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_4 abstract view
.subckt sky130_fd_sc_hd__clkinv_4 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211oi_4 abstract view
.subckt sky130_fd_sc_hd__a211oi_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_2 abstract view
.subckt sky130_fd_sc_hd__and2b_2 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or3_4 abstract view
.subckt sky130_fd_sc_hd__or3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or4b_2 abstract view
.subckt sky130_fd_sc_hd__or4b_2 A B C D_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkinv_2 abstract view
.subckt sky130_fd_sc_hd__clkinv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_2 abstract view
.subckt sky130_fd_sc_hd__o22a_2 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o21ba_4 abstract view
.subckt sky130_fd_sc_hd__o21ba_4 A1 A2 B1_N VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o22a_1 abstract view
.subckt sky130_fd_sc_hd__o22a_1 A1 A2 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211a_2 abstract view
.subckt sky130_fd_sc_hd__o211a_2 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand3_4 abstract view
.subckt sky130_fd_sc_hd__nand3_4 A B C VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and4bb_1 abstract view
.subckt sky130_fd_sc_hd__and4bb_1 A_N B_N C D VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_2 abstract view
.subckt sky130_fd_sc_hd__a2111o_2 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a22oi_2 abstract view
.subckt sky130_fd_sc_hd__a22oi_2 A1 A2 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a211o_4 abstract view
.subckt sky130_fd_sc_hd__a211o_4 A1 A2 B1 C1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o32ai_4 abstract view
.subckt sky130_fd_sc_hd__o32ai_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand4_1 abstract view
.subckt sky130_fd_sc_hd__nand4_1 A B C D VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o221ai_2 abstract view
.subckt sky130_fd_sc_hd__o221ai_2 A1 A2 B1 B2 C1 VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a2111o_1 abstract view
.subckt sky130_fd_sc_hd__a2111o_1 A1 A2 B1 C1 D1 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__o211ai_4 abstract view
.subckt sky130_fd_sc_hd__o211ai_4 A1 A2 B1 C1 VGND VNB VPB VPWR Y
.ends

.subckt user_proj_example io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ irq[0] irq[1] irq[2] la_data_in[0] la_data_in[100] la_data_in[101] la_data_in[102]
+ la_data_in[103] la_data_in[104] la_data_in[105] la_data_in[106] la_data_in[107]
+ la_data_in[108] la_data_in[109] la_data_in[10] la_data_in[110] la_data_in[111] la_data_in[112]
+ la_data_in[113] la_data_in[114] la_data_in[115] la_data_in[116] la_data_in[117]
+ la_data_in[118] la_data_in[119] la_data_in[11] la_data_in[120] la_data_in[121] la_data_in[122]
+ la_data_in[123] la_data_in[124] la_data_in[125] la_data_in[126] la_data_in[127]
+ la_data_in[12] la_data_in[13] la_data_in[14] la_data_in[15] la_data_in[16] la_data_in[17]
+ la_data_in[18] la_data_in[19] la_data_in[1] la_data_in[20] la_data_in[21] la_data_in[22]
+ la_data_in[23] la_data_in[24] la_data_in[25] la_data_in[26] la_data_in[27] la_data_in[28]
+ la_data_in[29] la_data_in[2] la_data_in[30] la_data_in[31] la_data_in[32] la_data_in[33]
+ la_data_in[34] la_data_in[35] la_data_in[36] la_data_in[37] la_data_in[38] la_data_in[39]
+ la_data_in[3] la_data_in[40] la_data_in[41] la_data_in[42] la_data_in[43] la_data_in[44]
+ la_data_in[45] la_data_in[46] la_data_in[47] la_data_in[48] la_data_in[49] la_data_in[4]
+ la_data_in[50] la_data_in[51] la_data_in[52] la_data_in[53] la_data_in[54] la_data_in[55]
+ la_data_in[56] la_data_in[57] la_data_in[58] la_data_in[59] la_data_in[5] la_data_in[60]
+ la_data_in[61] la_data_in[62] la_data_in[63] la_data_in[64] la_data_in[65] la_data_in[66]
+ la_data_in[67] la_data_in[68] la_data_in[69] la_data_in[6] la_data_in[70] la_data_in[71]
+ la_data_in[72] la_data_in[73] la_data_in[74] la_data_in[75] la_data_in[76] la_data_in[77]
+ la_data_in[78] la_data_in[79] la_data_in[7] la_data_in[80] la_data_in[81] la_data_in[82]
+ la_data_in[83] la_data_in[84] la_data_in[85] la_data_in[86] la_data_in[87] la_data_in[88]
+ la_data_in[89] la_data_in[8] la_data_in[90] la_data_in[91] la_data_in[92] la_data_in[93]
+ la_data_in[94] la_data_in[95] la_data_in[96] la_data_in[97] la_data_in[98] la_data_in[99]
+ la_data_in[9] la_data_out[0] la_data_out[100] la_data_out[101] la_data_out[102]
+ la_data_out[103] la_data_out[104] la_data_out[105] la_data_out[106] la_data_out[107]
+ la_data_out[108] la_data_out[109] la_data_out[10] la_data_out[110] la_data_out[111]
+ la_data_out[112] la_data_out[113] la_data_out[114] la_data_out[115] la_data_out[116]
+ la_data_out[117] la_data_out[118] la_data_out[119] la_data_out[11] la_data_out[120]
+ la_data_out[121] la_data_out[122] la_data_out[123] la_data_out[124] la_data_out[125]
+ la_data_out[126] la_data_out[127] la_data_out[12] la_data_out[13] la_data_out[14]
+ la_data_out[15] la_data_out[16] la_data_out[17] la_data_out[18] la_data_out[19]
+ la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22] la_data_out[23] la_data_out[24]
+ la_data_out[25] la_data_out[26] la_data_out[27] la_data_out[28] la_data_out[29]
+ la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32] la_data_out[33] la_data_out[34]
+ la_data_out[35] la_data_out[36] la_data_out[37] la_data_out[38] la_data_out[39]
+ la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42] la_data_out[43] la_data_out[44]
+ la_data_out[45] la_data_out[46] la_data_out[47] la_data_out[48] la_data_out[49]
+ la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52] la_data_out[53] la_data_out[54]
+ la_data_out[55] la_data_out[56] la_data_out[57] la_data_out[58] la_data_out[59]
+ la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62] la_data_out[63] la_data_out[64]
+ la_data_out[65] la_data_out[66] la_data_out[67] la_data_out[68] la_data_out[69]
+ la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72] la_data_out[73] la_data_out[74]
+ la_data_out[75] la_data_out[76] la_data_out[77] la_data_out[78] la_data_out[79]
+ la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82] la_data_out[83] la_data_out[84]
+ la_data_out[85] la_data_out[86] la_data_out[87] la_data_out[88] la_data_out[89]
+ la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92] la_data_out[93] la_data_out[94]
+ la_data_out[95] la_data_out[96] la_data_out[97] la_data_out[98] la_data_out[99]
+ la_data_out[9] la_oenb[0] la_oenb[100] la_oenb[101] la_oenb[102] la_oenb[103] la_oenb[104]
+ la_oenb[105] la_oenb[106] la_oenb[107] la_oenb[108] la_oenb[109] la_oenb[10] la_oenb[110]
+ la_oenb[111] la_oenb[112] la_oenb[113] la_oenb[114] la_oenb[115] la_oenb[116] la_oenb[117]
+ la_oenb[118] la_oenb[119] la_oenb[11] la_oenb[120] la_oenb[121] la_oenb[122] la_oenb[123]
+ la_oenb[124] la_oenb[125] la_oenb[126] la_oenb[127] la_oenb[12] la_oenb[13] la_oenb[14]
+ la_oenb[15] la_oenb[16] la_oenb[17] la_oenb[18] la_oenb[19] la_oenb[1] la_oenb[20]
+ la_oenb[21] la_oenb[22] la_oenb[23] la_oenb[24] la_oenb[25] la_oenb[26] la_oenb[27]
+ la_oenb[28] la_oenb[29] la_oenb[2] la_oenb[30] la_oenb[31] la_oenb[32] la_oenb[33]
+ la_oenb[34] la_oenb[35] la_oenb[36] la_oenb[37] la_oenb[38] la_oenb[39] la_oenb[3]
+ la_oenb[40] la_oenb[41] la_oenb[42] la_oenb[43] la_oenb[44] la_oenb[45] la_oenb[46]
+ la_oenb[47] la_oenb[48] la_oenb[49] la_oenb[4] la_oenb[50] la_oenb[51] la_oenb[52]
+ la_oenb[53] la_oenb[54] la_oenb[55] la_oenb[56] la_oenb[57] la_oenb[58] la_oenb[59]
+ la_oenb[5] la_oenb[60] la_oenb[61] la_oenb[62] la_oenb[63] la_oenb[64] la_oenb[65]
+ la_oenb[66] la_oenb[67] la_oenb[68] la_oenb[69] la_oenb[6] la_oenb[70] la_oenb[71]
+ la_oenb[72] la_oenb[73] la_oenb[74] la_oenb[75] la_oenb[76] la_oenb[77] la_oenb[78]
+ la_oenb[79] la_oenb[7] la_oenb[80] la_oenb[81] la_oenb[82] la_oenb[83] la_oenb[84]
+ la_oenb[85] la_oenb[86] la_oenb[87] la_oenb[88] la_oenb[89] la_oenb[8] la_oenb[90]
+ la_oenb[91] la_oenb[92] la_oenb[93] la_oenb[94] la_oenb[95] la_oenb[96] la_oenb[97]
+ la_oenb[98] la_oenb[99] la_oenb[9] vccd1 vssd1 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0]
+ wbs_adr_i[10] wbs_adr_i[11] wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15]
+ wbs_adr_i[16] wbs_adr_i[17] wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20]
+ wbs_adr_i[21] wbs_adr_i[22] wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26]
+ wbs_adr_i[27] wbs_adr_i[28] wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31]
+ wbs_adr_i[3] wbs_adr_i[4] wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9]
+ wbs_cyc_i wbs_dat_i[0] wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14]
+ wbs_dat_i[15] wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1]
+ wbs_dat_i[20] wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25]
+ wbs_dat_i[26] wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30]
+ wbs_dat_i[31] wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8]
+ wbs_dat_i[9] wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13]
+ wbs_dat_o[14] wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19]
+ wbs_dat_o[1] wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24]
+ wbs_dat_o[25] wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2]
+ wbs_dat_o[30] wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6]
+ wbs_dat_o[7] wbs_dat_o[8] wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3]
+ wbs_stb_i wbs_we_i
XTAP_199 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_188 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_177 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2106_ _2163_/A _2106_/B vssd1 vssd1 vccd1 vccd1 _2107_/B sky130_fd_sc_hd__nor2_1
XFILLER_39_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2037_ _2037_/A vssd1 vssd1 vccd1 vccd1 _2037_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__2455__A _2629_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3181__275 vssd1 vssd1 vccd1 vccd1 _3181__275/HI wbs_dat_o[3] sky130_fd_sc_hd__conb_1
XFILLER_23_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2939_ _2939_/A _2939_/B vssd1 vssd1 vccd1 vccd1 _2963_/B sky130_fd_sc_hd__xnor2_2
XFILLER_50_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2812__B _2812_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3165__259 vssd1 vssd1 vccd1 vccd1 _3165__259/HI la_data_out[116] sky130_fd_sc_hd__conb_1
XFILLER_24_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3059__153 vssd1 vssd1 vccd1 vccd1 _3059__153/HI io_out[19] sky130_fd_sc_hd__conb_1
X_2724_ _2725_/A _2725_/B _2599_/A vssd1 vssd1 vccd1 vccd1 _2724_/X sky130_fd_sc_hd__a21o_1
X_2655_ _2605_/X _2585_/X _2653_/X _2654_/Y vssd1 vssd1 vccd1 vccd1 _2657_/B sky130_fd_sc_hd__o211ai_2
X_1606_ _1643_/B _1606_/B vssd1 vssd1 vccd1 vccd1 _1621_/B sky130_fd_sc_hd__nor2_1
X_2586_ _2585_/A _2585_/B _2585_/C vssd1 vssd1 vccd1 vccd1 _2586_/Y sky130_fd_sc_hd__a21oi_2
X_1537_ _1521_/A _1521_/B _1536_/X vssd1 vssd1 vccd1 vccd1 _1559_/B sky130_fd_sc_hd__a21oi_2
XANTENNA__2185__A input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2807__B _2807_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2440_ _2363_/A _2440_/B vssd1 vssd1 vccd1 vccd1 _2451_/A sky130_fd_sc_hd__and2b_1
XFILLER_5_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2371_ _2371_/A _2371_/B vssd1 vssd1 vccd1 vccd1 _2371_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_64_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2707_ _2620_/A _2620_/B _2620_/C vssd1 vssd1 vccd1 vccd1 _2712_/A sky130_fd_sc_hd__a21oi_2
X_2638_ _2544_/A _2544_/B _2544_/C _2766_/A vssd1 vssd1 vccd1 vccd1 _2639_/B sky130_fd_sc_hd__a31o_1
XFILLER_59_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2569_ _2567_/X _2685_/A _2757_/A _2568_/X vssd1 vssd1 vccd1 vccd1 _2569_/X sky130_fd_sc_hd__a22o_1
XFILLER_28_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3187__281 vssd1 vssd1 vccd1 vccd1 _3187__281/HI wbs_dat_o[9] sky130_fd_sc_hd__conb_1
XFILLER_28_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input55_A la_data_in[59] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2818__A _2818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1639__A1 _1588_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1940_ _2043_/A _1944_/B vssd1 vssd1 vccd1 vccd1 _2036_/B sky130_fd_sc_hd__xor2_1
XFILLER_9_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1871_ _1871_/A _1903_/A _1905_/C vssd1 vssd1 vccd1 vccd1 _1876_/B sky130_fd_sc_hd__or3_1
XFILLER_6_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1616__B _1616_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2423_ _2492_/A _2492_/B vssd1 vssd1 vccd1 vccd1 _2494_/B sky130_fd_sc_hd__xnor2_2
X_2354_ _2354_/A _2354_/B _2354_/C vssd1 vssd1 vccd1 vccd1 _2354_/X sky130_fd_sc_hd__and3_1
X_2285_ _2309_/A _2285_/B vssd1 vssd1 vccd1 vccd1 _2361_/B sky130_fd_sc_hd__xnor2_1
XFILLER_64_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_507 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_518 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_529 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2070_ _2070_/A _2070_/B vssd1 vssd1 vccd1 vccd1 _2111_/A sky130_fd_sc_hd__nor2_1
XFILLER_62_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2972_ _2972_/A vssd1 vssd1 vccd1 vccd1 _2977_/A sky130_fd_sc_hd__clkbuf_4
X_1923_ _1923_/A _1972_/A vssd1 vssd1 vccd1 vccd1 _1923_/X sky130_fd_sc_hd__or2_1
XFILLER_15_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1854_ _2013_/A _2020_/A _1879_/B vssd1 vssd1 vccd1 vccd1 _1854_/Y sky130_fd_sc_hd__a21oi_1
X_1785_ _1813_/A _1785_/B vssd1 vssd1 vccd1 vccd1 _1786_/A sky130_fd_sc_hd__or2_1
XANTENNA__2760__A2 _2684_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2406_ _2406_/A _2406_/B vssd1 vssd1 vccd1 vccd1 _2684_/A sky130_fd_sc_hd__and2_1
X_2337_ _2337_/A vssd1 vssd1 vccd1 vccd1 _2567_/A sky130_fd_sc_hd__buf_2
X_2268_ _1929_/Y _2557_/A _2150_/A _1984_/A _2267_/X vssd1 vssd1 vccd1 vccd1 _2269_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_53_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2199_ _2199_/A _2199_/B _2199_/C vssd1 vssd1 vccd1 vccd1 _2201_/B sky130_fd_sc_hd__and3_1
XFILLER_37_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2751__A2 _2931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2368__A _2369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input18_A la_data_in[25] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2267__B2 _1979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1570_ _1530_/B _1568_/X _1569_/Y _1487_/B vssd1 vssd1 vccd1 vccd1 _1571_/B sky130_fd_sc_hd__a22o_2
XFILLER_6_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3092__186 vssd1 vssd1 vccd1 vccd1 _3092__186/HI la_data_out[11] sky130_fd_sc_hd__conb_1
XTAP_304 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_315 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_326 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_337 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_348 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_359 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2122_ _2059_/X _2062_/B _2060_/A vssd1 vssd1 vccd1 vccd1 _2123_/B sky130_fd_sc_hd__a21o_1
XFILLER_13_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2053_ _2053_/A _2053_/B _1954_/B vssd1 vssd1 vccd1 vccd1 _2066_/B sky130_fd_sc_hd__or3b_1
XFILLER_19_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2955_ _2955_/A _2955_/B vssd1 vssd1 vccd1 vccd1 _2960_/A sky130_fd_sc_hd__nor2_2
X_2886_ _2886_/A _2886_/B vssd1 vssd1 vccd1 vccd1 _2887_/B sky130_fd_sc_hd__xnor2_1
X_1906_ _1906_/A vssd1 vssd1 vccd1 vccd1 _2008_/A sky130_fd_sc_hd__inv_2
X_1837_ _1837_/A _1849_/B vssd1 vssd1 vccd1 vccd1 _1841_/A sky130_fd_sc_hd__xor2_1
X_1768_ _2013_/A vssd1 vssd1 vccd1 vccd1 _1821_/A sky130_fd_sc_hd__clkbuf_2
X_1699_ _2983_/A _1699_/B vssd1 vssd1 vccd1 vccd1 _1731_/B sky130_fd_sc_hd__xnor2_2
XTAP_860 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2188__A _2188_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1820__A _1979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput75 _2175_/Y vssd1 vssd1 vccd1 vccd1 la_data_out[74] sky130_fd_sc_hd__buf_2
XFILLER_0_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput86 _2903_/X vssd1 vssd1 vccd1 vccd1 la_data_out[85] sky130_fd_sc_hd__buf_2
XFILLER_48_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3020__114 vssd1 vssd1 vccd1 vccd1 _3020__114/HI io_oeb[17] sky130_fd_sc_hd__conb_1
XFILLER_12_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2412__B2 _2567_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2740_ _2740_/A vssd1 vssd1 vccd1 vccd1 _2740_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_8_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2671_ _2657_/A _2657_/C _2657_/B vssd1 vssd1 vccd1 vccd1 _2731_/A sky130_fd_sc_hd__a21bo_1
X_1622_ _1622_/A _1622_/B vssd1 vssd1 vccd1 vccd1 _1643_/A sky130_fd_sc_hd__and2_1
XFILLER_8_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1553_ _2939_/A _1553_/B vssd1 vssd1 vccd1 vccd1 _1590_/B sky130_fd_sc_hd__xnor2_2
XFILLER_4_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_134 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_156 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_145 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2479__A1 _2416_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_189 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_178 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_167 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2105_ _2105_/A _2105_/B vssd1 vssd1 vccd1 vccd1 _2106_/B sky130_fd_sc_hd__nor2_1
XANTENNA__2736__A _2919_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2036_ _2036_/A _2036_/B vssd1 vssd1 vccd1 vccd1 _2037_/A sky130_fd_sc_hd__and2_1
XFILLER_23_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2938_ _2863_/X _2930_/X _2932_/Y _2937_/X vssd1 vssd1 vccd1 vccd1 _2939_/B sky130_fd_sc_hd__a211o_1
X_2869_ _2819_/A _2468_/Y _2868_/Y vssd1 vssd1 vccd1 vccd1 _2870_/B sky130_fd_sc_hd__o21a_1
XFILLER_58_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_690 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2881__A1 _2083_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2633__A1 _2629_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2723_ _2723_/A _2723_/B vssd1 vssd1 vccd1 vccd1 _2728_/A sky130_fd_sc_hd__xor2_1
X_3098__192 vssd1 vssd1 vccd1 vccd1 _3098__192/HI la_data_out[17] sky130_fd_sc_hd__conb_1
X_2654_ _2653_/A _2653_/B _2652_/X vssd1 vssd1 vccd1 vccd1 _2654_/Y sky130_fd_sc_hd__o21bai_1
X_1605_ _1605_/A _1605_/B vssd1 vssd1 vccd1 vccd1 _1606_/B sky130_fd_sc_hd__and2_1
X_2585_ _2585_/A _2585_/B _2585_/C vssd1 vssd1 vccd1 vccd1 _2585_/X sky130_fd_sc_hd__and3_2
X_1536_ _2920_/A _2986_/A _1555_/B vssd1 vssd1 vccd1 vccd1 _1536_/X sky130_fd_sc_hd__and3_1
XFILLER_59_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2185__B _2185_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2019_ _2086_/A vssd1 vssd1 vccd1 vccd1 _2254_/A sky130_fd_sc_hd__buf_2
XFILLER_23_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1545__A _1605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3132__226 vssd1 vssd1 vccd1 vccd1 _3132__226/HI la_data_out[51] sky130_fd_sc_hd__conb_1
X_2370_ _2370_/A _2369_/X vssd1 vssd1 vccd1 vccd1 _2371_/B sky130_fd_sc_hd__or2b_1
XFILLER_49_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2854__A1 _2723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3026__120 vssd1 vssd1 vccd1 vccd1 _3026__120/HI io_oeb[23] sky130_fd_sc_hd__conb_1
XFILLER_17_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2706_ _2732_/A _2706_/B vssd1 vssd1 vccd1 vccd1 _2733_/A sky130_fd_sc_hd__xnor2_2
X_2637_ _2637_/A _2637_/B vssd1 vssd1 vccd1 vccd1 _2674_/A sky130_fd_sc_hd__and2_1
X_2568_ _2568_/A vssd1 vssd1 vccd1 vccd1 _2568_/X sky130_fd_sc_hd__clkbuf_2
X_1519_ _1539_/A _1539_/B vssd1 vssd1 vccd1 vccd1 _1555_/B sky130_fd_sc_hd__xnor2_4
X_2499_ input6/X _2647_/A _2498_/Y vssd1 vssd1 vccd1 vccd1 _2578_/A sky130_fd_sc_hd__a21oi_2
XFILLER_28_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input48_A la_data_in[52] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1870_ _1870_/A _1870_/B vssd1 vssd1 vccd1 vccd1 _1905_/C sky130_fd_sc_hd__and2_1
XFILLER_42_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2422_ _2818_/A _2422_/B vssd1 vssd1 vccd1 vccd1 _2492_/B sky130_fd_sc_hd__xnor2_4
XFILLER_43_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2353_ _2353_/A _2353_/B vssd1 vssd1 vccd1 vccd1 _2354_/C sky130_fd_sc_hd__xor2_2
X_2284_ _2284_/A _2284_/B vssd1 vssd1 vccd1 vccd1 _2285_/B sky130_fd_sc_hd__and2_1
XFILLER_37_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1999_ _1999_/A _2006_/C vssd1 vssd1 vccd1 vccd1 _2000_/B sky130_fd_sc_hd__xnor2_1
XFILLER_20_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2919__A _2919_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_519 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_508 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2971_ _2971_/A _2971_/B vssd1 vssd1 vccd1 vccd1 _2987_/A sky130_fd_sc_hd__nand2_1
X_1922_ _1816_/A _1916_/X _1919_/X _1921_/Y vssd1 vssd1 vccd1 vccd1 _1965_/A sky130_fd_sc_hd__a211o_2
X_1853_ _1975_/A vssd1 vssd1 vccd1 vccd1 _2020_/A sky130_fd_sc_hd__clkbuf_2
X_1784_ _1784_/A _1784_/B vssd1 vssd1 vccd1 vccd1 _1785_/B sky130_fd_sc_hd__nor2_1
X_3138__232 vssd1 vssd1 vccd1 vccd1 _3138__232/HI la_data_out[57] sky130_fd_sc_hd__conb_1
X_2405_ _2402_/X _2685_/A _2757_/A _2404_/X vssd1 vssd1 vccd1 vccd1 _2408_/A sky130_fd_sc_hd__a22o_1
XANTENNA__2739__A _2739_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2336_ _2775_/A _2819_/A vssd1 vssd1 vccd1 vccd1 _2336_/Y sky130_fd_sc_hd__nor2_1
X_2267_ _2021_/A _2096_/A _2099_/A _1979_/A vssd1 vssd1 vccd1 vccd1 _2267_/X sky130_fd_sc_hd__a22o_1
XFILLER_52_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2198_ _2197_/B _2197_/C _2254_/A vssd1 vssd1 vccd1 vccd1 _2199_/C sky130_fd_sc_hd__a21o_1
XANTENNA__2474__A _2546_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1818__A _1972_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2751__A3 _2931_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1553__A _2939_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2975__B1 _2973_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2990__A3 _2985_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_305 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_316 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_327 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_338 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_349 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2121_ _2121_/A _2120_/X vssd1 vssd1 vccd1 vccd1 _2123_/A sky130_fd_sc_hd__or2b_1
XFILLER_39_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2052_ _2052_/A _2052_/B vssd1 vssd1 vccd1 vccd1 _2112_/A sky130_fd_sc_hd__or2_1
XFILLER_19_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2954_ _2954_/A _2954_/B vssd1 vssd1 vccd1 vccd1 _2955_/B sky130_fd_sc_hd__nor2_1
X_2885_ _2944_/A _2885_/B vssd1 vssd1 vccd1 vccd1 _2886_/B sky130_fd_sc_hd__or2_1
X_1905_ _1906_/A _1905_/B _1905_/C vssd1 vssd1 vccd1 vccd1 _2006_/A sky130_fd_sc_hd__nand3b_2
X_1836_ _2086_/A _1836_/B vssd1 vssd1 vccd1 vccd1 _1849_/B sky130_fd_sc_hd__xnor2_1
X_1767_ input1/X vssd1 vssd1 vccd1 vccd1 _2013_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_1698_ _1736_/A _1698_/B vssd1 vssd1 vccd1 vccd1 _1703_/A sky130_fd_sc_hd__nor2_1
XTAP_861 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_850 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2188__B _2188_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2319_ _2192_/B _2192_/C _2258_/A _2192_/A vssd1 vssd1 vccd1 vccd1 _2325_/B sky130_fd_sc_hd__a211oi_1
XFILLER_57_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput65 _1766_/Y vssd1 vssd1 vccd1 vccd1 la_data_out[64] sky130_fd_sc_hd__buf_2
Xoutput76 _2244_/Y vssd1 vssd1 vccd1 vccd1 la_data_out[75] sky130_fd_sc_hd__buf_2
Xoutput87 _2960_/X vssd1 vssd1 vccd1 vccd1 la_data_out[86] sky130_fd_sc_hd__buf_2
XANTENNA_input30_A la_data_in[36] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2670_ _2663_/A _2603_/A _2719_/A _2663_/C vssd1 vssd1 vccd1 vccd1 _2670_/Y sky130_fd_sc_hd__o211ai_2
X_1621_ _1608_/B _1621_/B vssd1 vssd1 vccd1 vccd1 _1647_/A sky130_fd_sc_hd__and2b_1
X_3100__194 vssd1 vssd1 vccd1 vccd1 _3100__194/HI la_data_out[19] sky130_fd_sc_hd__conb_1
X_1552_ _1515_/X _2930_/X _1549_/Y _1551_/X vssd1 vssd1 vccd1 vccd1 _1553_/B sky130_fd_sc_hd__a211o_1
XTAP_135 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_157 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_146 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_179 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_168 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2104_ _2105_/A _2105_/B vssd1 vssd1 vccd1 vccd1 _2163_/A sky130_fd_sc_hd__and2_2
X_2035_ _2402_/A _2549_/A _2550_/A _2404_/A vssd1 vssd1 vccd1 vccd1 _2039_/A sky130_fd_sc_hd__a22o_1
XFILLER_22_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2937_ _2933_/X _2934_/X _2935_/X _2936_/X vssd1 vssd1 vccd1 vccd1 _2937_/X sky130_fd_sc_hd__a22o_1
XFILLER_50_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2868_ _2933_/A _2820_/X _2867_/X vssd1 vssd1 vccd1 vccd1 _2868_/Y sky130_fd_sc_hd__a21oi_1
X_1819_ _1926_/A vssd1 vssd1 vccd1 vccd1 _1979_/A sky130_fd_sc_hd__buf_2
X_2799_ _2797_/X _2799_/B vssd1 vssd1 vccd1 vccd1 _2801_/A sky130_fd_sc_hd__and2b_1
XFILLER_58_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_680 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_691 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3043__137 vssd1 vssd1 vccd1 vccd1 _3043__137/HI io_out[3] sky130_fd_sc_hd__conb_1
XFILLER_13_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1669__A0 input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2722_ _2722_/A _2722_/B vssd1 vssd1 vccd1 vccd1 _2723_/B sky130_fd_sc_hd__nor2_1
XFILLER_8_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2653_ _2653_/A _2653_/B _2652_/X vssd1 vssd1 vccd1 vccd1 _2653_/X sky130_fd_sc_hd__or3b_1
X_1604_ _1605_/A _1605_/B vssd1 vssd1 vccd1 vccd1 _1643_/B sky130_fd_sc_hd__nor2_1
X_2584_ _2657_/A _2584_/B vssd1 vssd1 vccd1 vccd1 _2585_/C sky130_fd_sc_hd__nor2_1
X_1535_ _2971_/A _1524_/B _1524_/A vssd1 vssd1 vccd1 vccd1 _1563_/B sky130_fd_sc_hd__o21ba_1
XFILLER_55_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2018_ _2018_/A vssd1 vssd1 vccd1 vccd1 _2032_/A sky130_fd_sc_hd__inv_2
XANTENNA__2085__B1 _2083_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2482__A _2577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2388__A1 _2608_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1561__A _1561_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2392__A _2629_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3171__265 vssd1 vssd1 vccd1 vccd1 _3171__265/HI la_data_out[122] sky130_fd_sc_hd__conb_1
XANTENNA__2551__B2 _2608_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2567__A _2567_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2705_ _2705_/A _2705_/B vssd1 vssd1 vccd1 vccd1 _2706_/B sky130_fd_sc_hd__xor2_2
X_2636_ _2636_/A _2636_/B _2636_/C vssd1 vssd1 vccd1 vccd1 _2637_/B sky130_fd_sc_hd__nand3_1
XANTENNA__2542__A1 _2543_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2567_ _2567_/A vssd1 vssd1 vccd1 vccd1 _2567_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_1518_ _2939_/A _1518_/B vssd1 vssd1 vccd1 vccd1 _1539_/B sky130_fd_sc_hd__xnor2_2
X_2498_ input6/X _2647_/A _2433_/A vssd1 vssd1 vccd1 vccd1 _2498_/Y sky130_fd_sc_hd__o21bai_1
XFILLER_28_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1556__A _1588_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1662__A2_N _2921_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3155__249 vssd1 vssd1 vccd1 vccd1 _3155__249/HI la_data_out[106] sky130_fd_sc_hd__conb_1
XFILLER_3_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3049__143 vssd1 vssd1 vccd1 vccd1 _3049__143/HI io_out[9] sky130_fd_sc_hd__conb_1
XFILLER_64_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2421_ _2758_/A _2609_/A _2419_/Y _2420_/X vssd1 vssd1 vccd1 vccd1 _2422_/B sky130_fd_sc_hd__a211o_1
X_2352_ _2623_/A _2352_/B vssd1 vssd1 vccd1 vccd1 _2353_/B sky130_fd_sc_hd__xnor2_2
XFILLER_36_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2283_ _2283_/A _2283_/B vssd1 vssd1 vccd1 vccd1 _2284_/B sky130_fd_sc_hd__nand2_1
XFILLER_37_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1998_ _2053_/B _1998_/B vssd1 vssd1 vccd1 vccd1 _2006_/C sky130_fd_sc_hd__xor2_1
XANTENNA__2763__A1 _2843_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2619_ _2620_/A _2620_/B _2620_/C vssd1 vssd1 vccd1 vccd1 _2624_/A sky130_fd_sc_hd__a21o_1
XFILLER_55_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA_input60_A la_data_in[63] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_509 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2809__A2 _2737_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2970_ _2970_/A _2970_/B _2970_/C vssd1 vssd1 vccd1 vccd1 _2971_/B sky130_fd_sc_hd__or3_1
XFILLER_15_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1921_ _1821_/A _2410_/A _2181_/B vssd1 vssd1 vccd1 vccd1 _1921_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_30_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1852_ input1/X _1879_/B _1975_/A vssd1 vssd1 vccd1 vccd1 _1852_/X sky130_fd_sc_hd__and3_1
XFILLER_30_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1783_ _1784_/A _1784_/B vssd1 vssd1 vccd1 vccd1 _1813_/A sky130_fd_sc_hd__and2_1
X_3177__271 vssd1 vssd1 vccd1 vccd1 _3177__271/HI wbs_ack_o sky130_fd_sc_hd__conb_1
X_2404_ _2404_/A vssd1 vssd1 vccd1 vccd1 _2404_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_57_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2335_ _2335_/A vssd1 vssd1 vccd1 vccd1 _2819_/A sky130_fd_sc_hd__buf_2
X_2266_ _2266_/A _2266_/B vssd1 vssd1 vccd1 vccd1 _2271_/A sky130_fd_sc_hd__xnor2_2
X_2197_ _2254_/A _2197_/B _2197_/C vssd1 vssd1 vccd1 vccd1 _2199_/B sky130_fd_sc_hd__nand3_1
XFILLER_25_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_52_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2474__B _2474_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2681__B1 _2258_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2975__B2 _2557_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_306 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_317 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_328 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_339 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2120_ _2120_/A _2120_/B vssd1 vssd1 vccd1 vccd1 _2120_/X sky130_fd_sc_hd__or2_1
X_2051_ _2051_/A _2067_/B vssd1 vssd1 vccd1 vccd1 _2112_/B sky130_fd_sc_hd__xor2_1
XFILLER_35_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2953_ _2954_/A _2954_/B vssd1 vssd1 vccd1 vccd1 _2955_/A sky130_fd_sc_hd__and2_1
XFILLER_22_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1904_ _1953_/B _1903_/C _1903_/A vssd1 vssd1 vccd1 vccd1 _1905_/B sky130_fd_sc_hd__a21o_1
XFILLER_15_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2884_ _2884_/A _2884_/B _2884_/C vssd1 vssd1 vccd1 vccd1 _2885_/B sky130_fd_sc_hd__and3_1
X_1835_ _1890_/A _2028_/A _2142_/A _1800_/A _1834_/X vssd1 vssd1 vccd1 vccd1 _1836_/B
+ sky130_fd_sc_hd__a221o_1
X_1766_ _1788_/A _1766_/B vssd1 vssd1 vccd1 vccd1 _1766_/Y sky130_fd_sc_hd__nor2_1
XFILLER_7_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1697_ _1697_/A _1697_/B _1697_/C vssd1 vssd1 vccd1 vccd1 _1698_/B sky130_fd_sc_hd__nor3_1
XTAP_862 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_851 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_840 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2318_ _2469_/A _2316_/X _2386_/A _2608_/A vssd1 vssd1 vccd1 vccd1 _2329_/B sky130_fd_sc_hd__a22o_1
X_2249_ _2464_/A vssd1 vssd1 vccd1 vccd1 _2385_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_25_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2957__B2 _2901_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1548__B _1548_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2709__A1 _1929_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput66 _1789_/Y vssd1 vssd1 vccd1 vccd1 la_data_out[65] sky130_fd_sc_hd__buf_2
Xoutput77 _2302_/Y vssd1 vssd1 vccd1 vccd1 la_data_out[76] sky130_fd_sc_hd__buf_2
Xoutput88 _1490_/X vssd1 vssd1 vccd1 vccd1 la_data_out[87] sky130_fd_sc_hd__buf_2
XFILLER_0_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input23_A la_data_in[2] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1620_ _1620_/A _1620_/B vssd1 vssd1 vccd1 vccd1 _1620_/Y sky130_fd_sc_hd__nor2_1
X_1551_ _1550_/X _2934_/X _2935_/X _2814_/X vssd1 vssd1 vccd1 vccd1 _1551_/X sky130_fd_sc_hd__a22o_1
XTAP_136 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_147 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_169 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_158 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2103_ _2209_/A _2103_/B vssd1 vssd1 vccd1 vccd1 _2105_/B sky130_fd_sc_hd__xnor2_1
XFILLER_54_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2034_ _2034_/A vssd1 vssd1 vccd1 vccd1 _2402_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_22_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2936_ _2936_/A vssd1 vssd1 vccd1 vccd1 _2936_/X sky130_fd_sc_hd__clkbuf_2
X_2867_ _2814_/A _2748_/X _2749_/X _2740_/X vssd1 vssd1 vccd1 vccd1 _2867_/X sky130_fd_sc_hd__a22o_1
X_1818_ _1972_/A vssd1 vssd1 vccd1 vccd1 _1926_/A sky130_fd_sc_hd__clkbuf_2
X_2798_ _2797_/B _2797_/C _2797_/A vssd1 vssd1 vccd1 vccd1 _2799_/B sky130_fd_sc_hd__a21o_1
X_1749_ _1749_/A _1749_/B vssd1 vssd1 vccd1 vccd1 _1750_/B sky130_fd_sc_hd__nor2_1
XFILLER_2_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_670 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2927__B _2927_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_681 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_692 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3082__176 vssd1 vssd1 vccd1 vccd1 _3082__176/HI la_data_out[1] sky130_fd_sc_hd__conb_1
XFILLER_14_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1602__B2 _1555_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1602__A1 _1557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2853__A _2901_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2721_ _2793_/B _2719_/Y _2669_/X _2670_/Y vssd1 vssd1 vccd1 vccd1 _2722_/B sky130_fd_sc_hd__o211a_1
XFILLER_8_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2652_ _2716_/A _2652_/B vssd1 vssd1 vccd1 vccd1 _2652_/X sky130_fd_sc_hd__and2_1
X_1603_ _1622_/A _1622_/B vssd1 vssd1 vccd1 vccd1 _1605_/B sky130_fd_sc_hd__xnor2_1
X_2583_ _2583_/A _2583_/B _2583_/C vssd1 vssd1 vccd1 vccd1 _2584_/B sky130_fd_sc_hd__and3_1
X_1534_ _1573_/B _1614_/A vssd1 vssd1 vccd1 vccd1 _1534_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__1932__A _2086_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2017_ _2269_/A _2088_/B vssd1 vssd1 vccd1 vccd1 _2018_/A sky130_fd_sc_hd__xnor2_1
XFILLER_42_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2919_ _2919_/A _2919_/B vssd1 vssd1 vccd1 vccd1 _2920_/A sky130_fd_sc_hd__or2_2
XFILLER_12_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3010__104 vssd1 vssd1 vccd1 vccd1 _3010__104/HI io_oeb[7] sky130_fd_sc_hd__conb_1
XFILLER_37_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1927__A _1972_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2704_ _2704_/A _2766_/B vssd1 vssd1 vccd1 vccd1 _2705_/B sky130_fd_sc_hd__xnor2_2
X_2635_ _2636_/B _2636_/C _2636_/A vssd1 vssd1 vccd1 vccd1 _2637_/A sky130_fd_sc_hd__a21o_1
XANTENNA__2542__A2 _2543_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2566_ _2775_/A _2827_/A vssd1 vssd1 vccd1 vccd1 _2566_/Y sky130_fd_sc_hd__nor2_1
X_1517_ _2933_/X _2930_/X _1513_/Y _1516_/X vssd1 vssd1 vccd1 vccd1 _1518_/B sky130_fd_sc_hd__a211o_1
X_2497_ input7/X vssd1 vssd1 vccd1 vccd1 _2647_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_4_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3194__288 vssd1 vssd1 vccd1 vccd1 _3194__288/HI wbs_dat_o[16] sky130_fd_sc_hd__conb_1
XANTENNA__1572__A _1616_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3088__182 vssd1 vssd1 vccd1 vccd1 _3088__182/HI la_data_out[7] sky130_fd_sc_hd__conb_1
XFILLER_34_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2420_ _2552_/A _2549_/A _2550_/A _2559_/A vssd1 vssd1 vccd1 vccd1 _2420_/X sky130_fd_sc_hd__a22o_1
X_2351_ _2404_/A _2685_/A _2483_/A _2430_/A _2350_/X vssd1 vssd1 vccd1 vccd1 _2352_/B
+ sky130_fd_sc_hd__a221o_1
X_2282_ _2283_/A _2283_/B vssd1 vssd1 vccd1 vccd1 _2284_/A sky130_fd_sc_hd__or2_1
XFILLER_29_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1997_ _2008_/A _2008_/B _1996_/X vssd1 vssd1 vccd1 vccd1 _1998_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__2763__A2 _2762_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2618_ _2824_/A _2618_/B vssd1 vssd1 vccd1 vccd1 _2620_/C sky130_fd_sc_hd__xnor2_2
XFILLER_0_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2549_ _2549_/A vssd1 vssd1 vccd1 vccd1 _2549_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_18_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3122__216 vssd1 vssd1 vccd1 vccd1 _3122__216/HI la_data_out[41] sky130_fd_sc_hd__conb_1
XFILLER_24_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3016__110 vssd1 vssd1 vccd1 vccd1 _3016__110/HI io_oeb[13] sky130_fd_sc_hd__conb_1
XFILLER_59_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input53_A la_data_in[57] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1920_ _2079_/A vssd1 vssd1 vccd1 vccd1 _2410_/A sky130_fd_sc_hd__buf_2
X_1851_ _1974_/A vssd1 vssd1 vccd1 vccd1 _1975_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_30_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1782_ _1805_/B _1782_/B vssd1 vssd1 vccd1 vccd1 _1784_/B sky130_fd_sc_hd__xor2_2
X_2403_ _2403_/A vssd1 vssd1 vccd1 vccd1 _2757_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__2101__A _2501_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2334_ _2400_/A _2333_/B _2332_/X vssd1 vssd1 vccd1 vccd1 _2354_/B sky130_fd_sc_hd__o21bai_1
XFILLER_57_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2265_ _1916_/X _1987_/A _2083_/X _2037_/A _2264_/X vssd1 vssd1 vccd1 vccd1 _2266_/B
+ sky130_fd_sc_hd__a221o_1
X_2196_ _2416_/A _2539_/A _2195_/X vssd1 vssd1 vccd1 vccd1 _2197_/C sky130_fd_sc_hd__a21oi_2
XFILLER_1_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2681__B2 _2557_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_52_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2011__A _2926_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1744__B _1745_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_307 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_318 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_329 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2050_ _1992_/A _1992_/B _2049_/Y vssd1 vssd1 vccd1 vccd1 _2067_/B sky130_fd_sc_hd__a21o_1
XFILLER_19_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2952_ _2952_/A _2952_/B vssd1 vssd1 vccd1 vccd1 _2954_/B sky130_fd_sc_hd__xnor2_4
X_1903_ _1903_/A _1953_/B _1903_/C vssd1 vssd1 vccd1 vccd1 _1906_/A sky130_fd_sc_hd__and3_1
X_2883_ _2884_/A _2884_/B _2884_/C vssd1 vssd1 vccd1 vccd1 _2944_/A sky130_fd_sc_hd__a21oi_2
XFILLER_30_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1834_ _2501_/A _1884_/B _1884_/A vssd1 vssd1 vccd1 vccd1 _1834_/X sky130_fd_sc_hd__and3b_1
X_1765_ _2393_/A _2434_/A _1775_/C vssd1 vssd1 vccd1 vccd1 _1766_/B sky130_fd_sc_hd__a21oi_1
X_1696_ _1697_/A _1697_/B _1697_/C vssd1 vssd1 vccd1 vccd1 _1736_/A sky130_fd_sc_hd__o21a_1
XTAP_852 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_841 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_830 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_863 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2317_ _2321_/A vssd1 vssd1 vccd1 vccd1 _2608_/A sky130_fd_sc_hd__buf_2
XANTENNA__2766__A _2766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2248_ _2380_/B vssd1 vssd1 vccd1 vccd1 _2464_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_38_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2179_ _2179_/A _2146_/B vssd1 vssd1 vccd1 vccd1 _2201_/A sky130_fd_sc_hd__or2b_1
XFILLER_53_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput67 _1815_/X vssd1 vssd1 vccd1 vccd1 la_data_out[66] sky130_fd_sc_hd__buf_2
XFILLER_0_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput78 _2371_/Y vssd1 vssd1 vccd1 vccd1 la_data_out[77] sky130_fd_sc_hd__buf_2
Xoutput89 _1534_/Y vssd1 vssd1 vccd1 vccd1 la_data_out[88] sky130_fd_sc_hd__buf_2
XANTENNA__2342__B1 _2141_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input16_A la_data_in[23] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3128__222 vssd1 vssd1 vccd1 vccd1 _3128__222/HI la_data_out[47] sky130_fd_sc_hd__conb_1
XFILLER_44_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_31_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1550_ _2922_/X vssd1 vssd1 vccd1 vccd1 _1550_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA_output84_A _2801_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_137 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_148 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_159 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2102_ _2273_/A _2411_/A _2560_/A _1807_/A _2101_/Y vssd1 vssd1 vccd1 vccd1 _2103_/B
+ sky130_fd_sc_hd__a221o_1
X_2033_ _2108_/A _2108_/B vssd1 vssd1 vccd1 vccd1 _2048_/A sky130_fd_sc_hd__xor2_1
XFILLER_35_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2935_ _2935_/A vssd1 vssd1 vccd1 vccd1 _2935_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_22_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2866_ _2939_/A _2866_/B vssd1 vssd1 vccd1 vccd1 _2912_/A sky130_fd_sc_hd__xnor2_2
X_1817_ _1817_/A vssd1 vssd1 vccd1 vccd1 _1984_/A sky130_fd_sc_hd__clkbuf_2
X_2797_ _2797_/A _2797_/B _2797_/C vssd1 vssd1 vccd1 vccd1 _2797_/X sky130_fd_sc_hd__and3_1
X_1748_ _1692_/A _1722_/Y _1747_/X vssd1 vssd1 vccd1 vccd1 _1749_/B sky130_fd_sc_hd__a21oi_1
X_1679_ _1711_/A _1679_/B vssd1 vssd1 vccd1 vccd1 _1681_/B sky130_fd_sc_hd__or2_1
XANTENNA_input8_A la_data_in[16] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_660 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_671 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_682 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_693 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2720_ _2669_/X _2670_/Y _2793_/B _2719_/Y vssd1 vssd1 vccd1 vccd1 _2722_/A sky130_fd_sc_hd__a211oi_1
XFILLER_8_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2651_ _2651_/A _2651_/B _2651_/C vssd1 vssd1 vccd1 vccd1 _2652_/B sky130_fd_sc_hd__or3_1
X_1602_ _1557_/A _1557_/B _1589_/B _1555_/B vssd1 vssd1 vccd1 vccd1 _1622_/B sky130_fd_sc_hd__o22ai_4
XFILLER_59_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2582_ _2583_/A _2583_/B _2583_/C vssd1 vssd1 vccd1 vccd1 _2657_/A sky130_fd_sc_hd__a21oi_2
X_1533_ _1533_/A _1533_/B vssd1 vssd1 vccd1 vccd1 _1614_/A sky130_fd_sc_hd__xnor2_1
XFILLER_55_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2016_ _1816_/A _1968_/C _2013_/X _2015_/Y vssd1 vssd1 vccd1 vccd1 _2088_/B sky130_fd_sc_hd__a211o_2
XFILLER_50_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2918_ _2992_/A _2918_/B vssd1 vssd1 vccd1 vccd1 _2942_/A sky130_fd_sc_hd__and2b_1
XFILLER_50_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2849_ _2850_/A _2896_/A vssd1 vssd1 vccd1 vccd1 _2904_/A sky130_fd_sc_hd__nor2_1
XFILLER_2_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2545__B1 _2544_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_490 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2954__A _2954_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2839__A1 _2026_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1927__B _1974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_13_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2703_ _2703_/A _2703_/B vssd1 vssd1 vccd1 vccd1 _2766_/B sky130_fd_sc_hd__nand2_1
X_2634_ _2814_/A _2811_/C _2633_/X vssd1 vssd1 vccd1 vccd1 _2636_/C sky130_fd_sc_hd__a21oi_2
X_2565_ _2623_/A vssd1 vssd1 vccd1 vccd1 _2862_/A sky130_fd_sc_hd__clkbuf_4
X_1516_ _1514_/X _2934_/X _2935_/X _1515_/X vssd1 vssd1 vccd1 vccd1 _1516_/X sky130_fd_sc_hd__a22o_1
X_3033__127 vssd1 vssd1 vccd1 vccd1 _3033__127/HI io_oeb[30] sky130_fd_sc_hd__conb_1
X_2496_ _2496_/A vssd1 vssd1 vccd1 vccd1 _2913_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_55_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1572__B _1616_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2350_ _1859_/Y _2827_/A _2403_/A _2273_/A vssd1 vssd1 vccd1 vccd1 _2350_/X sky130_fd_sc_hd__a2bb2o_1
X_2281_ _2281_/A _2281_/B vssd1 vssd1 vccd1 vccd1 _2283_/B sky130_fd_sc_hd__xnor2_1
XFILLER_64_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1996_ _2053_/A _1954_/B vssd1 vssd1 vccd1 vccd1 _1996_/X sky130_fd_sc_hd__or2b_1
X_2617_ _2819_/A _2965_/A _2616_/Y vssd1 vssd1 vccd1 vccd1 _2618_/B sky130_fd_sc_hd__o21a_1
XFILLER_0_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2548_ _2548_/A _2548_/B _2548_/C vssd1 vssd1 vccd1 vccd1 _2573_/B sky130_fd_sc_hd__or3_1
X_2479_ _2416_/A _2411_/A _2560_/A _2686_/A vssd1 vssd1 vccd1 vccd1 _2479_/X sky130_fd_sc_hd__a22o_1
XFILLER_55_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2009__A _2009_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3161__255 vssd1 vssd1 vccd1 vccd1 _3161__255/HI la_data_out[112] sky130_fd_sc_hd__conb_1
XFILLER_34_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3202__296 vssd1 vssd1 vccd1 vccd1 _3202__296/HI wbs_dat_o[24] sky130_fd_sc_hd__conb_1
XANTENNA__1508__A_N _1561_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input46_A la_data_in[50] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1850_ _1841_/A _1850_/B vssd1 vssd1 vccd1 vccd1 _1870_/A sky130_fd_sc_hd__and2b_1
X_1781_ _2181_/B _1800_/A vssd1 vssd1 vccd1 vccd1 _1782_/B sky130_fd_sc_hd__nand2_1
X_3003__97 vssd1 vssd1 vccd1 vccd1 _3003__97/HI io_oeb[0] sky130_fd_sc_hd__conb_1
XFILLER_6_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2402_ _2402_/A vssd1 vssd1 vccd1 vccd1 _2402_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_41_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2333_ _2400_/A _2333_/B _2332_/X vssd1 vssd1 vccd1 vccd1 _2354_/A sky130_fd_sc_hd__or3b_1
XANTENNA__1940__B _1944_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2264_ _1968_/C _1942_/A _1946_/A _1919_/C vssd1 vssd1 vccd1 vccd1 _2264_/X sky130_fd_sc_hd__a22o_1
X_2195_ _2131_/A _2316_/A _2386_/A _2071_/A vssd1 vssd1 vccd1 vccd1 _2195_/X sky130_fd_sc_hd__a22o_1
XFILLER_37_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3145__239 vssd1 vssd1 vccd1 vccd1 _3145__239/HI la_data_out[96] sky130_fd_sc_hd__conb_1
XFILLER_25_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1979_ _1979_/A _2022_/A vssd1 vssd1 vccd1 vccd1 _1979_/Y sky130_fd_sc_hd__nand2_1
X_3039__133 vssd1 vssd1 vccd1 vccd1 _3039__133/HI io_oeb[36] sky130_fd_sc_hd__conb_1
XFILLER_20_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_308 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_319 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2951_ _3000_/B _2951_/B vssd1 vssd1 vccd1 vccd1 _2952_/B sky130_fd_sc_hd__and2b_1
XANTENNA__1488__A _1488_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1902_ _1953_/A _1901_/B _1901_/C vssd1 vssd1 vccd1 vccd1 _1903_/C sky130_fd_sc_hd__a21o_1
XFILLER_15_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2882_ _2882_/A _2882_/B vssd1 vssd1 vccd1 vccd1 _2884_/C sky130_fd_sc_hd__nor2_1
X_1833_ input9/X input8/X vssd1 vssd1 vccd1 vccd1 _2501_/A sky130_fd_sc_hd__xnor2_4
X_1764_ _1764_/A _1764_/B vssd1 vssd1 vccd1 vccd1 _1764_/Y sky130_fd_sc_hd__xnor2_1
X_1695_ _2880_/X _2973_/Y _1694_/X vssd1 vssd1 vccd1 vccd1 _1697_/C sky130_fd_sc_hd__a21o_1
XTAP_853 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_842 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_831 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_820 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_864 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2316_ _2316_/A vssd1 vssd1 vccd1 vccd1 _2316_/X sky130_fd_sc_hd__clkbuf_2
X_2247_ _2623_/A _2185_/B _2201_/B vssd1 vssd1 vccd1 vccd1 _2308_/A sky130_fd_sc_hd__o21ba_1
XFILLER_38_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2178_ _2178_/A _2178_/B vssd1 vssd1 vccd1 vccd1 _2178_/Y sky130_fd_sc_hd__nand2_1
XFILLER_25_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput79 _2449_/Y vssd1 vssd1 vccd1 vccd1 la_data_out[78] sky130_fd_sc_hd__buf_2
XFILLER_0_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
Xoutput68 _1847_/X vssd1 vssd1 vccd1 vccd1 la_data_out[67] sky130_fd_sc_hd__buf_2
XANTENNA__2342__A1 _2410_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1580__B _2926_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3167__261 vssd1 vssd1 vccd1 vccd1 _3167__261/HI la_data_out[118] sky130_fd_sc_hd__conb_1
XFILLER_29_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2030__B1 _2026_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_138 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_149 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2101_ _2501_/A _2335_/A vssd1 vssd1 vccd1 vccd1 _2101_/Y sky130_fd_sc_hd__nor2_1
XFILLER_39_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2032_ _2032_/A _2032_/B vssd1 vssd1 vccd1 vccd1 _2108_/B sky130_fd_sc_hd__xnor2_1
XFILLER_35_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2934_ _2934_/A vssd1 vssd1 vccd1 vccd1 _2934_/X sky130_fd_sc_hd__clkbuf_2
X_2865_ _2258_/Y _2684_/X _2930_/A _2913_/A _2864_/X vssd1 vssd1 vccd1 vccd1 _2866_/B
+ sky130_fd_sc_hd__a221o_1
X_1816_ _1816_/A vssd1 vssd1 vccd1 vccd1 _2130_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_7_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2796_ _2795_/B _2795_/C _2795_/A vssd1 vssd1 vccd1 vccd1 _2797_/C sky130_fd_sc_hd__a21o_1
X_1747_ _1720_/A _1720_/B _1723_/Y vssd1 vssd1 vccd1 vccd1 _1747_/X sky130_fd_sc_hd__a21bo_1
X_1678_ _1678_/A _1678_/B vssd1 vssd1 vccd1 vccd1 _1679_/B sky130_fd_sc_hd__and2_1
XANTENNA__1681__A _1681_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_650 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_661 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_672 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_683 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_694 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2260__B1 _2258_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2650_ _2651_/A _2651_/B _2651_/C vssd1 vssd1 vccd1 vccd1 _2716_/A sky130_fd_sc_hd__o21ai_4
X_1601_ _1601_/A _1601_/B vssd1 vssd1 vccd1 vccd1 _1622_/A sky130_fd_sc_hd__nor2_1
XFILLER_8_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2581_ _2404_/X _2913_/B _2772_/A _2273_/X _2580_/X vssd1 vssd1 vccd1 vccd1 _2583_/C
+ sky130_fd_sc_hd__a221oi_4
X_1532_ _1532_/A _1532_/B vssd1 vssd1 vccd1 vccd1 _1533_/B sky130_fd_sc_hd__xnor2_4
XANTENNA__2597__A _2597_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2015_ _1968_/A _2071_/A _1968_/B vssd1 vssd1 vccd1 vccd1 _2015_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_63_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2917_ _2917_/A _2917_/B _2915_/Y vssd1 vssd1 vccd1 vccd1 _2918_/B sky130_fd_sc_hd__or3b_1
XFILLER_12_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2848_ _2857_/B _2848_/B vssd1 vssd1 vccd1 vccd1 _2896_/A sky130_fd_sc_hd__xnor2_2
X_2779_ _2808_/A _2779_/B _2779_/C vssd1 vssd1 vccd1 vccd1 _2808_/B sky130_fd_sc_hd__nor3_1
XTAP_480 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_491 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2954__B _2954_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2970__A _2970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2702_ _2919_/B _2702_/B _2702_/C _2702_/D vssd1 vssd1 vccd1 vccd1 _2703_/B sky130_fd_sc_hd__nand4_4
XFILLER_9_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2633_ _2629_/B _2316_/X _2698_/B _2692_/A vssd1 vssd1 vccd1 vccd1 _2633_/X sky130_fd_sc_hd__a22o_1
X_2564_ _2644_/A _2644_/B vssd1 vssd1 vccd1 vccd1 _2645_/A sky130_fd_sc_hd__xor2_2
X_1515_ _2740_/X vssd1 vssd1 vccd1 vccd1 _1515_/X sky130_fd_sc_hd__clkbuf_2
X_3072__166 vssd1 vssd1 vccd1 vccd1 _3072__166/HI io_out[32] sky130_fd_sc_hd__conb_1
X_2495_ input7/X _2647_/B vssd1 vssd1 vccd1 vccd1 _2496_/A sky130_fd_sc_hd__and2b_1
XFILLER_55_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2965__A _2965_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3207__301 vssd1 vssd1 vccd1 vccd1 _3207__301/HI wbs_dat_o[29] sky130_fd_sc_hd__conb_1
XFILLER_27_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1980__A2 _2775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2280_ _2273_/X _2347_/A _2403_/A _1899_/A _2279_/Y vssd1 vssd1 vccd1 vccd1 _2281_/B
+ sky130_fd_sc_hd__a221o_1
XANTENNA__2875__A _2911_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_144 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1799__A2 _1939_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1995_ _2052_/A _2052_/B vssd1 vssd1 vccd1 vccd1 _2053_/B sky130_fd_sc_hd__xnor2_1
XANTENNA__1971__A2 _2410_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2616_ _2758_/A _2820_/A _2615_/X vssd1 vssd1 vccd1 vccd1 _2616_/Y sky130_fd_sc_hd__a21oi_1
X_2547_ _2548_/B _2548_/C _2548_/A vssd1 vssd1 vccd1 vccd1 _2573_/A sky130_fd_sc_hd__o21ai_1
X_2478_ _2478_/A _2478_/B vssd1 vssd1 vccd1 vccd1 _2577_/A sky130_fd_sc_hd__xnor2_4
XFILLER_55_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input39_A la_data_in[44] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1780_ _2013_/B vssd1 vssd1 vccd1 vccd1 _2181_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_30_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2401_ _2528_/A _2400_/C _2400_/A vssd1 vssd1 vccd1 vccd1 _2425_/B sky130_fd_sc_hd__a21o_1
X_2332_ _2262_/A _2332_/B vssd1 vssd1 vccd1 vccd1 _2332_/X sky130_fd_sc_hd__and2b_1
XFILLER_34_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2263_ _2308_/A _2308_/B vssd1 vssd1 vccd1 vccd1 _2309_/A sky130_fd_sc_hd__xnor2_1
XFILLER_38_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2194_ _2194_/A vssd1 vssd1 vccd1 vccd1 _2539_/A sky130_fd_sc_hd__clkbuf_2
X_3184__278 vssd1 vssd1 vccd1 vccd1 _3184__278/HI wbs_dat_o[6] sky130_fd_sc_hd__conb_1
XANTENNA__2969__A1 _2970_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1949__A _2501_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1978_ _2337_/A _2028_/A _2142_/A _2020_/A vssd1 vssd1 vccd1 vccd1 _1978_/Y sky130_fd_sc_hd__a22oi_1
X_3078__172 vssd1 vssd1 vccd1 vccd1 _3078__172/HI irq[0] sky130_fd_sc_hd__conb_1
XFILLER_20_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_309 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2950_ _2950_/A _2950_/B vssd1 vssd1 vccd1 vccd1 _2951_/B sky130_fd_sc_hd__or2_1
XANTENNA__1488__B _1488_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1901_ _1953_/A _1901_/B _1901_/C vssd1 vssd1 vccd1 vccd1 _1953_/B sky130_fd_sc_hd__nand3_1
X_2881_ _2083_/X _2880_/X _2966_/A _2567_/X vssd1 vssd1 vccd1 vccd1 _2882_/B sky130_fd_sc_hd__a22o_1
X_1832_ _1832_/A vssd1 vssd1 vccd1 vccd1 _2142_/A sky130_fd_sc_hd__clkbuf_2
X_1763_ _1763_/A _1763_/B vssd1 vssd1 vccd1 vccd1 _1764_/B sky130_fd_sc_hd__xnor2_4
X_1694_ _1550_/X _1592_/X _1693_/X vssd1 vssd1 vccd1 vccd1 _1694_/X sky130_fd_sc_hd__a21o_1
XFILLER_7_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_810 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_843 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_832 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_821 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3112__206 vssd1 vssd1 vccd1 vccd1 _3112__206/HI la_data_out[31] sky130_fd_sc_hd__conb_1
XTAP_865 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_854 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2315_ _2454_/A _2530_/A _2391_/A _2314_/Y vssd1 vssd1 vccd1 vccd1 _2330_/A sky130_fd_sc_hd__a31o_1
X_2246_ _2281_/A vssd1 vssd1 vccd1 vccd1 _2623_/A sky130_fd_sc_hd__buf_2
X_2177_ _2177_/A _2177_/B vssd1 vssd1 vccd1 vccd1 _2177_/X sky130_fd_sc_hd__or2_1
XFILLER_25_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3006__100 vssd1 vssd1 vccd1 vccd1 _3006__100/HI io_oeb[3] sky130_fd_sc_hd__conb_1
XFILLER_15_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_25_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xoutput69 _1875_/Y vssd1 vssd1 vccd1 vccd1 la_data_out[68] sky130_fd_sc_hd__buf_2
XFILLER_17_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_320 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2030__A1 _2568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_139 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2100_ _2206_/A _2206_/B vssd1 vssd1 vccd1 vccd1 _2335_/A sky130_fd_sc_hd__nand2_1
XFILLER_39_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2031_ _2254_/A _2031_/B vssd1 vssd1 vccd1 vccd1 _2032_/B sky130_fd_sc_hd__xnor2_2
XFILLER_47_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_0 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_62_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2933_ _2933_/A vssd1 vssd1 vccd1 vccd1 _2933_/X sky130_fd_sc_hd__clkbuf_2
X_2864_ _2936_/A _2934_/A _2935_/A _2863_/X vssd1 vssd1 vccd1 vccd1 _2864_/X sky130_fd_sc_hd__a22o_1
X_1815_ _1815_/A vssd1 vssd1 vccd1 vccd1 _1815_/X sky130_fd_sc_hd__clkbuf_1
X_2795_ _2795_/A _2795_/B _2795_/C vssd1 vssd1 vccd1 vccd1 _2797_/B sky130_fd_sc_hd__nand3_1
X_1746_ _1746_/A _1746_/B vssd1 vssd1 vccd1 vccd1 _1750_/A sky130_fd_sc_hd__nand2_1
X_1677_ _1678_/A _1678_/B vssd1 vssd1 vccd1 vccd1 _1711_/A sky130_fd_sc_hd__nor2_2
XTAP_640 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_651 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_695 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_662 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_673 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_684 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2229_ _2289_/B _2228_/B _2228_/C vssd1 vssd1 vccd1 vccd1 _2230_/C sky130_fd_sc_hd__a21oi_1
XFILLER_53_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2017__B _2088_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input21_A la_data_in[28] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_17_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1600_ _1599_/B _1600_/B vssd1 vssd1 vccd1 vccd1 _1601_/B sky130_fd_sc_hd__and2b_1
XFILLER_8_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2580_ _1859_/Y _2964_/A _2774_/A _2434_/A vssd1 vssd1 vccd1 vccd1 _2580_/X sky130_fd_sc_hd__a2bb2o_1
X_1531_ _1576_/A _1577_/A vssd1 vssd1 vccd1 vccd1 _1532_/B sky130_fd_sc_hd__or2b_2
XFILLER_4_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2014_ _2189_/A vssd1 vssd1 vccd1 vccd1 _2071_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_35_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2916_ _2917_/A _2917_/B _2915_/Y vssd1 vssd1 vccd1 vccd1 _2992_/A sky130_fd_sc_hd__o21ba_1
XFILLER_31_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2847_ _2847_/A _2847_/B vssd1 vssd1 vccd1 vccd1 _2848_/B sky130_fd_sc_hd__xnor2_2
X_3118__212 vssd1 vssd1 vccd1 vccd1 _3118__212/HI la_data_out[37] sky130_fd_sc_hd__conb_1
X_2778_ _2807_/A _2807_/B vssd1 vssd1 vccd1 vccd1 _2779_/C sky130_fd_sc_hd__xnor2_1
X_1729_ _2880_/X _2871_/Y _1728_/X vssd1 vssd1 vccd1 vccd1 _1730_/B sky130_fd_sc_hd__a21oi_1
XTAP_470 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_481 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_492 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_562 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2861__B1_N _2812_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2701_ _2702_/B _2702_/C _2702_/D _2919_/B vssd1 vssd1 vccd1 vccd1 _2703_/A sky130_fd_sc_hd__a31o_2
XFILLER_9_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2632_ _2973_/A _2973_/B _2538_/A vssd1 vssd1 vccd1 vccd1 _2636_/B sky130_fd_sc_hd__a21o_2
X_2563_ _2824_/A _2563_/B vssd1 vssd1 vccd1 vccd1 _2644_/B sky130_fd_sc_hd__xnor2_1
X_1514_ _2814_/X vssd1 vssd1 vccd1 vccd1 _1514_/X sky130_fd_sc_hd__clkbuf_2
X_2494_ _2494_/A _2494_/B vssd1 vssd1 vccd1 vccd1 _2504_/B sky130_fd_sc_hd__nor2_1
XFILLER_55_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2311__A _2464_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1597__A _1597_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3095__189 vssd1 vssd1 vccd1 vccd1 _3095__189/HI la_data_out[14] sky130_fd_sc_hd__conb_1
XFILLER_37_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1994_ _1952_/A _1952_/B _1993_/X vssd1 vssd1 vccd1 vccd1 _2052_/B sky130_fd_sc_hd__a21oi_1
XFILLER_9_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2615_ _2552_/A _2748_/A _2749_/A _2829_/A vssd1 vssd1 vccd1 vccd1 _2615_/X sky130_fd_sc_hd__a22o_1
X_2546_ _2546_/A _2474_/B vssd1 vssd1 vccd1 vccd1 _2548_/A sky130_fd_sc_hd__or2b_1
X_2477_ _2559_/A _2609_/A _2258_/Y _2037_/X _2476_/X vssd1 vssd1 vccd1 vccd1 _2478_/B
+ sky130_fd_sc_hd__a221o_2
XFILLER_56_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3023__117 vssd1 vssd1 vccd1 vccd1 _3023__117/HI io_oeb[20] sky130_fd_sc_hd__conb_1
XFILLER_6_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2400_ _2400_/A _2528_/A _2400_/C vssd1 vssd1 vccd1 vccd1 _2425_/A sky130_fd_sc_hd__nand3_1
X_2331_ _2330_/B _2330_/C _2330_/A vssd1 vssd1 vccd1 vccd1 _2333_/B sky130_fd_sc_hd__a21oi_4
X_2262_ _2262_/A _2332_/B vssd1 vssd1 vccd1 vccd1 _2308_/B sky130_fd_sc_hd__xor2_1
XFILLER_27_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2193_ _2377_/A _2418_/A _2418_/B vssd1 vssd1 vccd1 vccd1 _2197_/B sky130_fd_sc_hd__or3_2
XFILLER_37_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_392 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1977_ _1977_/A _1977_/B vssd1 vssd1 vccd1 vccd1 _2775_/A sky130_fd_sc_hd__xnor2_4
XANTENNA__1965__A _1965_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2529_ _2529_/A _2529_/B vssd1 vssd1 vccd1 vccd1 _2529_/X sky130_fd_sc_hd__and2_1
XFILLER_56_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input51_A la_data_in[55] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2648__A1 _1888_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1900_ _2612_/A _1900_/B vssd1 vssd1 vccd1 vccd1 _1901_/C sky130_fd_sc_hd__xnor2_1
XFILLER_15_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2880_ _2880_/A vssd1 vssd1 vccd1 vccd1 _2880_/X sky130_fd_sc_hd__clkbuf_2
X_1831_ _1831_/A _1861_/C vssd1 vssd1 vccd1 vccd1 _1832_/A sky130_fd_sc_hd__nor2_1
XFILLER_30_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1762_ _1762_/A _1762_/B vssd1 vssd1 vccd1 vccd1 _1763_/B sky130_fd_sc_hd__xnor2_4
XFILLER_11_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1693_ _1761_/A _1502_/X _1761_/B _1514_/X vssd1 vssd1 vccd1 vccd1 _1693_/X sky130_fd_sc_hd__a22o_1
XFILLER_7_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_800 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_844 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_833 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_822 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_811 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3151__245 vssd1 vssd1 vccd1 vccd1 _3151__245/HI la_data_out[102] sky130_fd_sc_hd__conb_1
XTAP_866 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_855 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2314_ _2530_/A _2314_/B vssd1 vssd1 vccd1 vccd1 _2314_/Y sky130_fd_sc_hd__nor2_1
X_2245_ _2220_/B _2220_/C _2220_/A vssd1 vssd1 vccd1 vccd1 _2361_/A sky130_fd_sc_hd__a21bo_1
XFILLER_38_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2176_ _2176_/A _2176_/B vssd1 vssd1 vccd1 vccd1 _2230_/A sky130_fd_sc_hd__nand2_1
XFILLER_21_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3135__229 vssd1 vssd1 vccd1 vccd1 _3135__229/HI la_data_out[54] sky130_fd_sc_hd__conb_1
XFILLER_21_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2869__A1 _2819_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2030_ _2568_/A _2194_/A _2026_/Y _2027_/X _2029_/X vssd1 vssd1 vccd1 vccd1 _2031_/B
+ sky130_fd_sc_hd__a221o_2
X_3029__123 vssd1 vssd1 vccd1 vccd1 _3029__123/HI io_oeb[26] sky130_fd_sc_hd__conb_1
XFILLER_62_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_1 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2932_ _2932_/A _2932_/B vssd1 vssd1 vccd1 vccd1 _2932_/Y sky130_fd_sc_hd__nor2_1
X_2863_ _2863_/A vssd1 vssd1 vccd1 vccd1 _2863_/X sky130_fd_sc_hd__clkbuf_2
X_1814_ _1845_/B _1814_/B vssd1 vssd1 vccd1 vccd1 _1815_/A sky130_fd_sc_hd__and2b_1
X_2794_ _2523_/X _2518_/B _2603_/Y _2793_/X _2593_/X vssd1 vssd1 vccd1 vccd1 _2795_/C
+ sky130_fd_sc_hd__a311o_1
XFILLER_30_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1745_ _1745_/A _1745_/B vssd1 vssd1 vccd1 vccd1 _1746_/B sky130_fd_sc_hd__or2_1
XFILLER_7_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1676_ _1638_/A _1638_/B _1674_/B _1636_/B vssd1 vssd1 vccd1 vccd1 _1678_/B sky130_fd_sc_hd__o2bb2a_1
XTAP_630 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_641 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_652 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_663 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_674 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_685 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_696 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2228_ _2289_/B _2228_/B _2228_/C vssd1 vssd1 vccd1 vccd1 _2305_/A sky130_fd_sc_hd__and3_1
XFILLER_26_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2159_ _2159_/A _2159_/B vssd1 vssd1 vccd1 vccd1 _2160_/B sky130_fd_sc_hd__or2_1
XFILLER_41_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input14_A la_data_in[21] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1530_ _2996_/A _1530_/B vssd1 vssd1 vccd1 vccd1 _1577_/A sky130_fd_sc_hd__nand2_1
XFILLER_4_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2711__B1 _2712_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2013_ _2013_/A _2013_/B _2189_/A vssd1 vssd1 vccd1 vccd1 _2013_/X sky130_fd_sc_hd__and3_1
XFILLER_48_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2915_ _2141_/Y _2880_/X _2914_/X vssd1 vssd1 vccd1 vccd1 _2915_/Y sky130_fd_sc_hd__a21oi_1
X_2846_ _2846_/A _2846_/B vssd1 vssd1 vccd1 vccd1 _2847_/B sky130_fd_sc_hd__xor2_2
X_3157__251 vssd1 vssd1 vccd1 vccd1 _3157__251/HI la_data_out[108] sky130_fd_sc_hd__conb_1
X_2777_ _2568_/X _2772_/X _2776_/X vssd1 vssd1 vccd1 vccd1 _2807_/B sky130_fd_sc_hd__a21oi_4
X_1728_ _1761_/A _1592_/X _1761_/B _1550_/X vssd1 vssd1 vccd1 vccd1 _1728_/X sky130_fd_sc_hd__a22o_1
XFILLER_2_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1659_ _1659_/A _1716_/A vssd1 vssd1 vccd1 vccd1 _1659_/Y sky130_fd_sc_hd__nor2_1
XANTENNA_input6_A la_data_in[14] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_460 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_471 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_482 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_493 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2472__A2 _2468_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2700_ _2700_/A vssd1 vssd1 vccd1 vccd1 _2919_/B sky130_fd_sc_hd__buf_2
XFILLER_9_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2631_ _2630_/A _2630_/B _2630_/C _2630_/D vssd1 vssd1 vccd1 vccd1 _2973_/B sky130_fd_sc_hd__o31ai_2
XFILLER_57_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2562_ _2557_/X _2141_/Y _2820_/A _2686_/A _2561_/X vssd1 vssd1 vccd1 vccd1 _2563_/B
+ sky130_fd_sc_hd__a221o_1
X_1513_ _2932_/A _2468_/Y vssd1 vssd1 vccd1 vccd1 _1513_/Y sky130_fd_sc_hd__nor2_1
XFILLER_4_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2493_ _2493_/A vssd1 vssd1 vccd1 vccd1 _2494_/A sky130_fd_sc_hd__inv_2
XFILLER_55_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2129__A _2129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2829_ _2829_/A vssd1 vssd1 vccd1 vccd1 _2913_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_48_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_290 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2151__B2 _1939_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1878__A _2023_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1597__B _1597_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_6_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1993_ _1937_/A _1993_/B vssd1 vssd1 vccd1 vccd1 _1993_/X sky130_fd_sc_hd__and2b_1
XFILLER_9_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2614_ _2744_/A _2614_/B _2614_/C vssd1 vssd1 vccd1 vccd1 _2620_/B sky130_fd_sc_hd__nand3_2
X_2545_ _2544_/B _2544_/C _2544_/A vssd1 vssd1 vccd1 vccd1 _2548_/C sky130_fd_sc_hd__a21oi_1
X_2476_ _2134_/C _1943_/A _1947_/A _2131_/A vssd1 vssd1 vccd1 vccd1 _2476_/X sky130_fd_sc_hd__a22o_1
XFILLER_55_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2322__A _2322_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3062__156 vssd1 vssd1 vccd1 vccd1 _3062__156/HI io_out[22] sky130_fd_sc_hd__conb_1
XFILLER_15_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3103__197 vssd1 vssd1 vccd1 vccd1 _3103__197/HI la_data_out[22] sky130_fd_sc_hd__conb_1
X_2330_ _2330_/A _2330_/B _2330_/C vssd1 vssd1 vccd1 vccd1 _2400_/A sky130_fd_sc_hd__and3_2
XFILLER_2_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2261_ _2636_/A _2261_/B vssd1 vssd1 vccd1 vccd1 _2332_/B sky130_fd_sc_hd__xnor2_1
X_2192_ _2192_/A _2192_/B _2192_/C vssd1 vssd1 vccd1 vccd1 _2418_/B sky130_fd_sc_hd__and3_1
XFILLER_37_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1976_ _1976_/A _1976_/B vssd1 vssd1 vccd1 vccd1 _1977_/B sky130_fd_sc_hd__nor2_2
X_2528_ _2528_/A _2528_/B vssd1 vssd1 vccd1 vccd1 _2528_/Y sky130_fd_sc_hd__nor2_1
XFILLER_29_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2459_ _2461_/B vssd1 vssd1 vccd1 vccd1 _2459_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input44_A la_data_in[49] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1830_ _1830_/A _1830_/B vssd1 vssd1 vccd1 vccd1 _1861_/C sky130_fd_sc_hd__xnor2_1
XFILLER_42_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1761_ _1761_/A _1761_/B vssd1 vssd1 vccd1 vccd1 _1762_/B sky130_fd_sc_hd__nand2_2
XFILLER_51_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1692_ _1692_/A _1722_/A vssd1 vssd1 vccd1 vccd1 _1692_/Y sky130_fd_sc_hd__xnor2_1
XTAP_801 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3190__284 vssd1 vssd1 vccd1 vccd1 _3190__284/HI wbs_dat_o[12] sky130_fd_sc_hd__conb_1
XTAP_834 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_823 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_812 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2313_ _2464_/A _2534_/A _2313_/S vssd1 vssd1 vccd1 vccd1 _2314_/B sky130_fd_sc_hd__mux2_1
XTAP_856 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_845 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2244_ _2244_/A _2244_/B vssd1 vssd1 vccd1 vccd1 _2244_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_38_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2175_ _2175_/A _2175_/B vssd1 vssd1 vccd1 vccd1 _2175_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_26_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1959_ _1959_/A _1959_/B vssd1 vssd1 vccd1 vccd1 _1959_/X sky130_fd_sc_hd__or2_1
XFILLER_0_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3174__268 vssd1 vssd1 vccd1 vccd1 _3174__268/HI la_data_out[125] sky130_fd_sc_hd__conb_1
XFILLER_4_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2318__B2 _2608_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2869__A2 _2468_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3068__162 vssd1 vssd1 vccd1 vccd1 _3068__162/HI io_out[28] sky130_fd_sc_hd__conb_1
XFILLER_47_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_2 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_50_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2931_ _2931_/A _2931_/B vssd1 vssd1 vccd1 vccd1 _2932_/B sky130_fd_sc_hd__nand2_1
X_2862_ _2862_/A vssd1 vssd1 vccd1 vccd1 _2939_/A sky130_fd_sc_hd__clkbuf_8
XFILLER_30_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1813_ _1813_/A _1813_/B _1811_/X vssd1 vssd1 vccd1 vccd1 _1814_/B sky130_fd_sc_hd__or3b_1
X_2793_ _2793_/A _2793_/B vssd1 vssd1 vccd1 vccd1 _2793_/X sky130_fd_sc_hd__or2_1
XFILLER_30_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1744_ _1745_/A _1745_/B vssd1 vssd1 vccd1 vccd1 _1746_/A sky130_fd_sc_hd__nand2_1
X_1675_ _1675_/A _1675_/B vssd1 vssd1 vccd1 vccd1 _1678_/A sky130_fd_sc_hd__xnor2_1
XFILLER_58_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_620 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_631 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_642 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_653 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_664 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_675 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_686 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_697 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2227_ _2163_/A _2163_/B _2226_/X vssd1 vssd1 vccd1 vccd1 _2228_/C sky130_fd_sc_hd__a21o_1
X_2158_ _2159_/A _2159_/B vssd1 vssd1 vccd1 vccd1 _2160_/A sky130_fd_sc_hd__nand2_1
XFILLER_26_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2089_ _2032_/A _2032_/B _2088_/X vssd1 vssd1 vccd1 vccd1 _2090_/B sky130_fd_sc_hd__a21boi_4
XFILLER_26_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2012_ _2188_/A vssd1 vssd1 vccd1 vccd1 _2189_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_63_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2914_ _2758_/X _2772_/A _2966_/A _2686_/X _2913_/X vssd1 vssd1 vccd1 vccd1 _2914_/X
+ sky130_fd_sc_hd__a221o_1
X_2845_ _2845_/A _2845_/B vssd1 vssd1 vccd1 vccd1 _2846_/B sky130_fd_sc_hd__xor2_2
X_3196__290 vssd1 vssd1 vccd1 vccd1 _3196__290/HI wbs_dat_o[18] sky130_fd_sc_hd__conb_1
X_2776_ _2567_/X _2773_/X _2966_/A _2402_/X _2775_/Y vssd1 vssd1 vccd1 vccd1 _2776_/X
+ sky130_fd_sc_hd__a221o_1
X_1727_ _2983_/A _1699_/B _1697_/A vssd1 vssd1 vccd1 vccd1 _1730_/A sky130_fd_sc_hd__a21o_1
X_1658_ _1655_/X _1656_/X _1657_/Y _1618_/B vssd1 vssd1 vccd1 vccd1 _1692_/A sky130_fd_sc_hd__a22o_1
X_1589_ _1636_/B _1589_/B vssd1 vssd1 vccd1 vccd1 _1600_/B sky130_fd_sc_hd__xnor2_1
XTAP_450 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_461 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_472 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_483 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_494 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_37_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_39_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2630_ _2630_/A _2630_/B _2630_/C _2630_/D vssd1 vssd1 vccd1 vccd1 _2973_/A sky130_fd_sc_hd__or4_1
X_2561_ _2829_/A _2748_/A _2749_/A _2758_/A vssd1 vssd1 vccd1 vccd1 _2561_/X sky130_fd_sc_hd__a22o_1
X_1512_ _2818_/A _1538_/B vssd1 vssd1 vccd1 vccd1 _1539_/A sky130_fd_sc_hd__xnor2_4
X_2492_ _2492_/A _2492_/B vssd1 vssd1 vccd1 vccd1 _2504_/A sky130_fd_sc_hd__and2_1
XFILLER_4_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_534 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2828_ _2965_/A _2932_/A vssd1 vssd1 vccd1 vccd1 _2828_/Y sky130_fd_sc_hd__nor2_1
X_2759_ _2829_/A _2934_/A _2935_/A _2758_/X vssd1 vssd1 vccd1 vccd1 _2759_/X sky130_fd_sc_hd__a22o_1
XFILLER_2_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_280 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_291 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_9_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3108__202 vssd1 vssd1 vccd1 vccd1 _3108__202/HI la_data_out[27] sky130_fd_sc_hd__conb_1
XFILLER_52_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1992_ _1992_/A _1992_/B vssd1 vssd1 vccd1 vccd1 _2052_/A sky130_fd_sc_hd__xnor2_1
X_2613_ _2614_/B _2614_/C _2744_/A vssd1 vssd1 vccd1 vccd1 _2620_/A sky130_fd_sc_hd__a21o_1
X_2544_ _2544_/A _2544_/B _2544_/C vssd1 vssd1 vccd1 vccd1 _2548_/B sky130_fd_sc_hd__and3_1
X_2475_ _2528_/A _2528_/B vssd1 vssd1 vccd1 vccd1 _2529_/A sky130_fd_sc_hd__xor2_1
XFILLER_28_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1979__A _1979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_43_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2322__B _2322_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_504 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2260_ _2559_/A _2539_/A _2258_/Y _2027_/X _2259_/X vssd1 vssd1 vccd1 vccd1 _2261_/B
+ sky130_fd_sc_hd__a221o_2
XFILLER_1_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2191_ _2192_/B _2192_/C _2192_/A vssd1 vssd1 vccd1 vccd1 _2418_/A sky130_fd_sc_hd__a21oi_1
XFILLER_18_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1975_ _1975_/A _1975_/B vssd1 vssd1 vccd1 vccd1 _1976_/B sky130_fd_sc_hd__nor2_1
XFILLER_21_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2527_ _2527_/A _2527_/B vssd1 vssd1 vccd1 vccd1 _2527_/Y sky130_fd_sc_hd__nand2_1
X_2458_ _2458_/A _2462_/B _2458_/C vssd1 vssd1 vccd1 vccd1 _2461_/B sky130_fd_sc_hd__and3_1
XFILLER_29_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2389_ _2390_/B _2390_/C _2700_/A vssd1 vssd1 vccd1 vccd1 _2399_/B sky130_fd_sc_hd__a21o_1
XFILLER_16_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3085__179 vssd1 vssd1 vccd1 vccd1 _3085__179/HI la_data_out[4] sky130_fd_sc_hd__conb_1
XFILLER_36_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2333__A _2400_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input37_A la_data_in[42] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2508__A _2525_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1760_ _1760_/A _1760_/B vssd1 vssd1 vccd1 vccd1 _1762_/A sky130_fd_sc_hd__xnor2_2
XFILLER_7_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1691_ _1723_/A _1723_/B vssd1 vssd1 vccd1 vccd1 _1722_/A sky130_fd_sc_hd__xnor2_1
XTAP_835 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_824 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_813 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_802 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2312_ _2534_/A vssd1 vssd1 vccd1 vccd1 _2391_/A sky130_fd_sc_hd__clkbuf_2
XTAP_857 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_846 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2243_ _2173_/B _2175_/B _2242_/Y vssd1 vssd1 vccd1 vccd1 _2244_/B sky130_fd_sc_hd__o21ai_1
X_2174_ _2120_/X _2123_/B _2121_/A vssd1 vssd1 vccd1 vccd1 _2175_/B sky130_fd_sc_hd__a21oi_1
XFILLER_26_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2137__B _2188_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1958_ _1959_/A _1959_/B vssd1 vssd1 vccd1 vccd1 _1960_/A sky130_fd_sc_hd__and2_1
X_1889_ _1979_/A _1829_/A _1832_/A _1924_/A vssd1 vssd1 vccd1 vccd1 _1892_/C sky130_fd_sc_hd__a22o_1
X_3013__107 vssd1 vssd1 vccd1 vccd1 _3013__107/HI io_oeb[10] sky130_fd_sc_hd__conb_1
XFILLER_56_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_8_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2930_ _2930_/A vssd1 vssd1 vccd1 vccd1 _2930_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_30_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2861_ _2988_/A _2836_/B _2812_/B vssd1 vssd1 vccd1 vccd1 _2909_/A sky130_fd_sc_hd__o21ba_1
X_1812_ _1813_/A _1813_/B _1811_/X vssd1 vssd1 vccd1 vccd1 _1845_/B sky130_fd_sc_hd__o21ba_1
XFILLER_30_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2792_ _2664_/B _2791_/Y _2719_/Y vssd1 vssd1 vccd1 vccd1 _2795_/B sky130_fd_sc_hd__a21oi_2
X_1743_ _1743_/A _1743_/B vssd1 vssd1 vccd1 vccd1 _1745_/B sky130_fd_sc_hd__xnor2_4
X_1674_ _1700_/B _1674_/B vssd1 vssd1 vccd1 vccd1 _1675_/B sky130_fd_sc_hd__xnor2_1
XFILLER_7_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_610 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_621 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_632 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_643 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_654 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_665 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_676 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_698 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2226_ _2162_/B _2226_/B vssd1 vssd1 vccd1 vccd1 _2226_/X sky130_fd_sc_hd__and2b_1
XTAP_687 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2157_ _2205_/A _2157_/B vssd1 vssd1 vccd1 vccd1 _2159_/B sky130_fd_sc_hd__xnor2_1
XFILLER_26_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2088_ _2209_/A _2088_/B vssd1 vssd1 vccd1 vccd1 _2088_/X sky130_fd_sc_hd__or2_1
XFILLER_21_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2484__A1 _2568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3141__235 vssd1 vssd1 vccd1 vccd1 _3141__235/HI la_data_out[60] sky130_fd_sc_hd__conb_1
XFILLER_12_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2011_ _2926_/A vssd1 vssd1 vccd1 vccd1 _2269_/A sky130_fd_sc_hd__inv_2
XFILLER_63_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_35_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2913_ _2913_/A _2913_/B vssd1 vssd1 vccd1 vccd1 _2913_/X sky130_fd_sc_hd__and2_1
X_2844_ _2888_/A _2844_/B vssd1 vssd1 vccd1 vccd1 _2845_/B sky130_fd_sc_hd__nor2_1
X_2775_ _2775_/A _2964_/A vssd1 vssd1 vccd1 vccd1 _2775_/Y sky130_fd_sc_hd__nor2_1
X_1726_ _1726_/A _1709_/B vssd1 vssd1 vccd1 vccd1 _1738_/B sky130_fd_sc_hd__or2b_1
X_1657_ _1657_/A _1657_/B vssd1 vssd1 vccd1 vccd1 _1657_/Y sky130_fd_sc_hd__nor2_1
X_1588_ _2988_/A _1588_/B vssd1 vssd1 vccd1 vccd1 _1589_/B sky130_fd_sc_hd__or2_2
XTAP_440 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_451 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_462 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_473 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_484 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_495 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2209_ _2209_/A _2209_/B vssd1 vssd1 vccd1 vccd1 _2210_/B sky130_fd_sc_hd__xnor2_1
XFILLER_39_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3125__219 vssd1 vssd1 vccd1 vccd1 _3125__219/HI la_data_out[44] sky130_fd_sc_hd__conb_1
XFILLER_14_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3019__113 vssd1 vssd1 vccd1 vccd1 _3019__113/HI io_oeb[16] sky130_fd_sc_hd__conb_1
XFILLER_1_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2560_ _2560_/A vssd1 vssd1 vccd1 vccd1 _2749_/A sky130_fd_sc_hd__clkbuf_2
X_1511_ _2926_/A _1511_/B vssd1 vssd1 vccd1 vccd1 _1538_/B sky130_fd_sc_hd__xnor2_4
X_2491_ _2526_/A _2491_/B vssd1 vssd1 vccd1 vccd1 _2527_/A sky130_fd_sc_hd__xnor2_1
XFILLER_4_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2332__A_N _2262_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2145__B _2145_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2827_ _2827_/A vssd1 vssd1 vccd1 vccd1 _2932_/A sky130_fd_sc_hd__clkbuf_2
X_2758_ _2758_/A vssd1 vssd1 vccd1 vccd1 _2758_/X sky130_fd_sc_hd__clkbuf_2
X_1709_ _1726_/A _1709_/B vssd1 vssd1 vccd1 vccd1 _1711_/C sky130_fd_sc_hd__xnor2_2
X_2689_ _2862_/A _2689_/B vssd1 vssd1 vccd1 vccd1 _2770_/B sky130_fd_sc_hd__xnor2_2
XFILLER_59_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_48_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_270 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_281 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_292 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_226 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2336__A _2775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2678__A1 _2739_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3147__241 vssd1 vssd1 vccd1 vccd1 _3147__241/HI la_data_out[98] sky130_fd_sc_hd__conb_1
XFILLER_45_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1653__A2 _1613_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1991_ _2478_/A _1991_/B vssd1 vssd1 vccd1 vccd1 _1992_/B sky130_fd_sc_hd__xnor2_2
XFILLER_9_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2612_ _2612_/A vssd1 vssd1 vccd1 vccd1 _2744_/A sky130_fd_sc_hd__buf_2
X_2543_ _2636_/A _2543_/B _2543_/C vssd1 vssd1 vccd1 vccd1 _2544_/C sky130_fd_sc_hd__nand3_1
X_2474_ _2546_/A _2474_/B vssd1 vssd1 vccd1 vccd1 _2528_/B sky130_fd_sc_hd__xor2_1
XFILLER_28_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2841__A1 _2843_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_516 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2190_ _2190_/A _2189_/X vssd1 vssd1 vccd1 vccd1 _2192_/A sky130_fd_sc_hd__or2b_1
XFILLER_49_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1974_ _1974_/A _1975_/B vssd1 vssd1 vccd1 vccd1 _1976_/A sky130_fd_sc_hd__and2_1
X_2526_ _2526_/A _2491_/B vssd1 vssd1 vccd1 vccd1 _2526_/X sky130_fd_sc_hd__or2b_1
X_2457_ _2130_/X _2394_/X _2454_/X _2456_/Y vssd1 vssd1 vccd1 vccd1 _2546_/A sky130_fd_sc_hd__a211o_2
XFILLER_29_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2388_ _2608_/A _2539_/A _2387_/X vssd1 vssd1 vccd1 vccd1 _2390_/C sky130_fd_sc_hd__a21oi_1
XFILLER_28_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2333__B _2333_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1690_ _1690_/A _1690_/B vssd1 vssd1 vccd1 vccd1 _1723_/B sky130_fd_sc_hd__xnor2_4
XTAP_825 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_814 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_803 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2311_ _2464_/B vssd1 vssd1 vccd1 vccd1 _2534_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_858 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_847 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_836 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2242_ _2242_/A _2242_/B vssd1 vssd1 vccd1 vccd1 _2242_/Y sky130_fd_sc_hd__nand2_1
XFILLER_25_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2173_ _2173_/A _2173_/B vssd1 vssd1 vccd1 vccd1 _2175_/A sky130_fd_sc_hd__nor2_1
XFILLER_53_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2434__A _2434_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1957_ _1963_/A _1963_/B vssd1 vssd1 vccd1 vccd1 _1959_/B sky130_fd_sc_hd__xor2_1
X_1888_ _2027_/A _1888_/B vssd1 vssd1 vccd1 vccd1 _1892_/B sky130_fd_sc_hd__and2_1
X_2509_ _2523_/A _2523_/B vssd1 vssd1 vccd1 vccd1 _2509_/Y sky130_fd_sc_hd__nor2_1
X_3052__146 vssd1 vssd1 vccd1 vccd1 _3052__146/HI io_out[12] sky130_fd_sc_hd__conb_1
XFILLER_56_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_4 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_140 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2860_ _2877_/A vssd1 vssd1 vccd1 vccd1 _2988_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_1811_ _1845_/A _1811_/B vssd1 vssd1 vccd1 vccd1 _1811_/X sky130_fd_sc_hd__or2_1
X_2791_ _2791_/A vssd1 vssd1 vccd1 vccd1 _2791_/Y sky130_fd_sc_hd__inv_2
X_1742_ _1689_/A _1714_/B _1741_/Y _1690_/A _1754_/B vssd1 vssd1 vccd1 vccd1 _1743_/B
+ sky130_fd_sc_hd__a221o_2
XANTENNA__1765__A1 _2393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1673_ _2988_/X _1673_/B vssd1 vssd1 vccd1 vccd1 _1674_/B sky130_fd_sc_hd__or2_1
XFILLER_7_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_600 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_611 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_622 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_633 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_644 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_655 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_666 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_677 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_699 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2225_ _2289_/A _2224_/C _2160_/A vssd1 vssd1 vccd1 vccd1 _2228_/B sky130_fd_sc_hd__a21bo_1
XTAP_688 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2156_ _2402_/A _1988_/A _2154_/Y _2155_/X vssd1 vssd1 vccd1 vccd1 _2157_/B sky130_fd_sc_hd__a211o_1
XFILLER_26_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2087_ _2129_/A _2087_/B vssd1 vssd1 vccd1 vccd1 _2090_/A sky130_fd_sc_hd__xor2_4
XFILLER_53_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2989_ _2989_/A _2942_/A vssd1 vssd1 vccd1 vccd1 _2989_/X sky130_fd_sc_hd__or2b_1
XFILLER_57_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3180__274 vssd1 vssd1 vccd1 vccd1 _3180__274/HI wbs_dat_o[2] sky130_fd_sc_hd__conb_1
XFILLER_9_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2010_ input2/X vssd1 vssd1 vccd1 vccd1 _2926_/A sky130_fd_sc_hd__buf_6
XFILLER_63_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2912_ _2912_/A _2912_/B vssd1 vssd1 vccd1 vccd1 _2917_/B sky130_fd_sc_hd__and2_1
XFILLER_31_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2843_ _2843_/A _2843_/B _2843_/C vssd1 vssd1 vccd1 vccd1 _2844_/B sky130_fd_sc_hd__and3_1
X_2774_ _2774_/A vssd1 vssd1 vccd1 vccd1 _2966_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_1725_ _1725_/A _1725_/B vssd1 vssd1 vccd1 vccd1 _1725_/Y sky130_fd_sc_hd__xnor2_1
X_1656_ _1613_/A _1613_/B _1655_/B _1655_/A vssd1 vssd1 vccd1 vccd1 _1656_/X sky130_fd_sc_hd__a22o_1
X_1587_ _1629_/B _1587_/B vssd1 vssd1 vccd1 vccd1 _1636_/B sky130_fd_sc_hd__or2_2
XTAP_430 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_441 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_452 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_463 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_474 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_485 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_496 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2208_ _1888_/B _2557_/A _2150_/A _1939_/A _2207_/X vssd1 vssd1 vccd1 vccd1 _2209_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_39_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3164__258 vssd1 vssd1 vccd1 vccd1 _3164__258/HI la_data_out[115] sky130_fd_sc_hd__conb_1
X_2139_ _2139_/A _2139_/B vssd1 vssd1 vccd1 vccd1 _2187_/C sky130_fd_sc_hd__nand2_2
XFILLER_26_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3205__299 vssd1 vssd1 vccd1 vccd1 _3205__299/HI wbs_dat_o[27] sky130_fd_sc_hd__conb_1
XFILLER_22_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3058__152 vssd1 vssd1 vccd1 vccd1 _3058__152/HI io_out[18] sky130_fd_sc_hd__conb_1
XFILLER_49_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input12_A la_data_in[1] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1510_ _2557_/X _2871_/Y _1509_/X vssd1 vssd1 vccd1 vccd1 _1511_/B sky130_fd_sc_hd__a21oi_2
X_2490_ _2529_/A _2529_/B vssd1 vssd1 vccd1 vccd1 _2491_/B sky130_fd_sc_hd__xor2_1
XFILLER_4_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1656__B1 _1655_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2826_ _2825_/A _2825_/B _2825_/C _2825_/D vssd1 vssd1 vccd1 vccd1 _2833_/B sky130_fd_sc_hd__o22ai_4
X_2757_ _2757_/A vssd1 vssd1 vccd1 vccd1 _2935_/A sky130_fd_sc_hd__clkbuf_2
X_1708_ _1738_/A _1708_/B vssd1 vssd1 vccd1 vccd1 _1709_/B sky130_fd_sc_hd__and2_1
X_2688_ _2083_/X _2684_/X _2756_/A _2567_/X _2687_/X vssd1 vssd1 vccd1 vccd1 _2689_/B
+ sky130_fd_sc_hd__a221o_1
X_1639_ _1588_/B _1637_/B _1601_/A vssd1 vssd1 vccd1 vccd1 _1640_/B sky130_fd_sc_hd__a21o_1
XFILLER_58_124 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input4_A la_data_in[12] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_260 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_271 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_282 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_293 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1521__A _1521_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2336__B _2819_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2678__A2 _2468_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1886__B1 input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_38_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3186__280 vssd1 vssd1 vccd1 vccd1 _3186__280/HI wbs_dat_o[8] sky130_fd_sc_hd__conb_1
XFILLER_18_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1990_ _2404_/A _2549_/A _2609_/A _1899_/A _1989_/X vssd1 vssd1 vccd1 vccd1 _1991_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_20_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2262__A _2262_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2611_ _2936_/A _2609_/X _2610_/X vssd1 vssd1 vccd1 vccd1 _2614_/C sky130_fd_sc_hd__a21oi_2
XFILLER_55_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2542_ _2543_/B _2543_/C _2636_/A vssd1 vssd1 vccd1 vccd1 _2544_/B sky130_fd_sc_hd__a21o_1
X_2473_ _2700_/A _2473_/B vssd1 vssd1 vccd1 vccd1 _2474_/B sky130_fd_sc_hd__xnor2_4
XFILLER_56_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2809_ _2738_/A _2737_/A _2768_/A vssd1 vssd1 vccd1 vccd1 _2858_/B sky130_fd_sc_hd__o21ai_2
XANTENNA__2900__A _2956_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_61_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1973_ _1923_/X _1887_/B _1972_/X _1928_/B _1924_/X vssd1 vssd1 vccd1 vccd1 _1977_/A
+ sky130_fd_sc_hd__a311o_4
X_2525_ _2525_/A _2525_/B vssd1 vssd1 vccd1 vccd1 _2525_/Y sky130_fd_sc_hd__nand2_1
X_2456_ _2393_/A _2697_/A _2454_/B vssd1 vssd1 vccd1 vccd1 _2456_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_29_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2387_ _2740_/A _2316_/X _2698_/B _2469_/A vssd1 vssd1 vccd1 vccd1 _2387_/X sky130_fd_sc_hd__a22o_1
XFILLER_45_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2495__A_N input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2502__B2 _2434_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_826 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_815 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_804 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2310_ _2310_/A vssd1 vssd1 vccd1 vccd1 _2530_/A sky130_fd_sc_hd__inv_2
XTAP_859 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_848 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_837 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2241_ _2241_/A _2240_/X vssd1 vssd1 vccd1 vccd1 _2244_/A sky130_fd_sc_hd__or2b_1
XFILLER_38_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2172_ _2242_/A _2242_/B vssd1 vssd1 vccd1 vccd1 _2173_/B sky130_fd_sc_hd__nor2_1
XFILLER_18_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1956_ _2008_/B _1956_/B vssd1 vssd1 vccd1 vccd1 _1963_/B sky130_fd_sc_hd__xor2_1
X_1887_ _1887_/A _1887_/B vssd1 vssd1 vccd1 vccd1 _1888_/B sky130_fd_sc_hd__xnor2_4
XFILLER_0_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3091__185 vssd1 vssd1 vccd1 vccd1 _3091__185/HI la_data_out[10] sky130_fd_sc_hd__conb_1
X_2508_ _2525_/A _2525_/B vssd1 vssd1 vccd1 vccd1 _2523_/B sky130_fd_sc_hd__xnor2_1
X_2439_ _2510_/A _2439_/B vssd1 vssd1 vccd1 vccd1 _2451_/B sky130_fd_sc_hd__xnor2_1
XFILLER_56_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1513__B _2468_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input42_A la_data_in[47] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_5 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1810_ _1810_/A _1810_/B vssd1 vssd1 vccd1 vccd1 _1811_/B sky130_fd_sc_hd__nor2_1
XFILLER_30_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2790_ _2790_/A _2790_/B vssd1 vssd1 vccd1 vccd1 _2795_/A sky130_fd_sc_hd__nand2_1
X_1741_ _1741_/A _1741_/B vssd1 vssd1 vccd1 vccd1 _1741_/Y sky130_fd_sc_hd__nor2_1
X_1672_ _1697_/B _1672_/B vssd1 vssd1 vccd1 vccd1 _1700_/B sky130_fd_sc_hd__nor2_2
XANTENNA__1765__A2 _2434_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2270__A _2271_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3075__169 vssd1 vssd1 vccd1 vccd1 _3075__169/HI io_out[35] sky130_fd_sc_hd__conb_1
XFILLER_7_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_601 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_612 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_623 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_634 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_645 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_656 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_667 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2224_ _2160_/A _2289_/A _2224_/C vssd1 vssd1 vccd1 vccd1 _2289_/B sky130_fd_sc_hd__nand3b_1
XTAP_678 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_689 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2155_ _1916_/X _1943_/A _1946_/A _2021_/A vssd1 vssd1 vccd1 vccd1 _2155_/X sky130_fd_sc_hd__a22o_1
XFILLER_38_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2086_ _2086_/A _2086_/B vssd1 vssd1 vccd1 vccd1 _2087_/B sky130_fd_sc_hd__xnor2_4
XFILLER_22_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2988_ _2988_/A vssd1 vssd1 vccd1 vccd1 _2988_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_21_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1939_ _1939_/A vssd1 vssd1 vccd1 vccd1 _2273_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__2180__A _2322_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1747__A2 _1720_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1683__A1 _1597_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2911_ _2911_/A _2911_/B vssd1 vssd1 vccd1 vccd1 _2917_/A sky130_fd_sc_hd__nor2_1
X_2842_ _2842_/A vssd1 vssd1 vccd1 vccd1 _2888_/A sky130_fd_sc_hd__inv_2
X_2773_ _2913_/B vssd1 vssd1 vccd1 vccd1 _2773_/X sky130_fd_sc_hd__clkbuf_2
X_1724_ _1692_/A _1722_/Y _1723_/Y vssd1 vssd1 vccd1 vccd1 _1725_/B sky130_fd_sc_hd__a21bo_1
X_1655_ _1655_/A _1655_/B vssd1 vssd1 vccd1 vccd1 _1655_/X sky130_fd_sc_hd__or2_1
X_1586_ _1663_/A _1586_/B vssd1 vssd1 vccd1 vccd1 _1587_/B sky130_fd_sc_hd__nor2_1
XFILLER_58_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_420 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_431 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_442 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_453 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_464 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_475 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2207_ _2034_/A _2096_/A _2099_/A _1984_/A vssd1 vssd1 vccd1 vccd1 _2207_/X sky130_fd_sc_hd__a22o_1
XTAP_486 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_497 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2138_ _2138_/A _2188_/A vssd1 vssd1 vccd1 vccd1 _2139_/B sky130_fd_sc_hd__or2_1
XFILLER_26_236 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2069_ _2069_/A vssd1 vssd1 vccd1 vccd1 _2070_/A sky130_fd_sc_hd__inv_2
XANTENNA__1729__A2 _2871_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3097__191 vssd1 vssd1 vccd1 vccd1 _3097__191/HI la_data_out[16] sky130_fd_sc_hd__conb_1
XFILLER_49_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2723__A _2723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2825_ _2825_/A _2825_/B _2825_/C _2825_/D vssd1 vssd1 vccd1 vccd1 _2884_/A sky130_fd_sc_hd__or4_4
XFILLER_8_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2756_ _2756_/A vssd1 vssd1 vccd1 vccd1 _2930_/A sky130_fd_sc_hd__clkbuf_2
X_1707_ _1707_/A _1707_/B vssd1 vssd1 vccd1 vccd1 _1708_/B sky130_fd_sc_hd__or2_1
X_2687_ _2758_/A _2934_/A _2757_/A _2686_/X vssd1 vssd1 vccd1 vccd1 _2687_/X sky130_fd_sc_hd__a22o_1
X_1638_ _1638_/A _1638_/B vssd1 vssd1 vccd1 vccd1 _1640_/A sky130_fd_sc_hd__xor2_2
X_3131__225 vssd1 vssd1 vccd1 vccd1 _3131__225/HI la_data_out[50] sky130_fd_sc_hd__conb_1
XFILLER_58_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1569_ _2999_/A _1576_/A vssd1 vssd1 vccd1 vccd1 _1569_/Y sky130_fd_sc_hd__nor2_1
XTAP_250 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_261 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_272 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_283 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_294 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_350 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_64_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_548 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1583__B1 _2973_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2610_ _2740_/A _2549_/X _2550_/X _2747_/A vssd1 vssd1 vccd1 vccd1 _2610_/X sky130_fd_sc_hd__a22o_1
X_2541_ _2740_/A _2811_/C _2540_/X vssd1 vssd1 vccd1 vccd1 _2543_/C sky130_fd_sc_hd__a21oi_2
X_3115__209 vssd1 vssd1 vccd1 vccd1 _3115__209/HI la_data_out[34] sky130_fd_sc_hd__conb_1
X_2472_ _2538_/A _2468_/Y _2471_/Y vssd1 vssd1 vccd1 vccd1 _2473_/B sky130_fd_sc_hd__o21a_1
XFILLER_48_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3009__103 vssd1 vssd1 vccd1 vccd1 _3009__103/HI io_oeb[6] sky130_fd_sc_hd__conb_1
XFILLER_51_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2808_ _2808_/A _2808_/B vssd1 vssd1 vccd1 vccd1 _2846_/A sky130_fd_sc_hd__or2_1
XANTENNA__2900__B _2958_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2739_ _2739_/A _2921_/A _2921_/B vssd1 vssd1 vccd1 vccd1 _2745_/B sky130_fd_sc_hd__or3_1
XFILLER_3_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_59_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2817__B1 _2818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1972_ _1972_/A _1974_/A vssd1 vssd1 vccd1 vccd1 _1972_/X sky130_fd_sc_hd__or2_1
XFILLER_14_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1547__A0 _2926_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2524_ _2524_/A _2524_/B vssd1 vssd1 vccd1 vccd1 _2524_/Y sky130_fd_sc_hd__nand2_1
X_2455_ _2629_/B vssd1 vssd1 vccd1 vccd1 _2697_/A sky130_fd_sc_hd__clkbuf_2
X_2386_ _2386_/A vssd1 vssd1 vccd1 vccd1 _2698_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_45_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2911__A _2911_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3137__231 vssd1 vssd1 vccd1 vccd1 _3137__231/HI la_data_out[56] sky130_fd_sc_hd__conb_1
XFILLER_59_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_42_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_816 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_805 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_849 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_838 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_827 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2240_ _2240_/A _2240_/B vssd1 vssd1 vccd1 vccd1 _2240_/X sky130_fd_sc_hd__or2_1
X_2171_ _2242_/A _2242_/B vssd1 vssd1 vccd1 vccd1 _2173_/A sky130_fd_sc_hd__and2_1
XFILLER_61_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1955_ _2008_/A _2006_/A vssd1 vssd1 vccd1 vccd1 _1956_/B sky130_fd_sc_hd__nand2_1
X_1886_ input8/X _1923_/A input9/X vssd1 vssd1 vccd1 vccd1 _1887_/B sky130_fd_sc_hd__o21a_2
XFILLER_0_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2507_ _2524_/A _2524_/B vssd1 vssd1 vccd1 vccd1 _2525_/B sky130_fd_sc_hd__xor2_1
X_2438_ _2438_/A _2438_/B vssd1 vssd1 vccd1 vccd1 _2439_/B sky130_fd_sc_hd__or2_1
X_2369_ _2369_/A _2369_/B vssd1 vssd1 vccd1 vccd1 _2369_/X sky130_fd_sc_hd__or2_1
XFILLER_44_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_24_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1931__B1 _1929_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input35_A la_data_in[40] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_35_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1740_ _1753_/A _1740_/B vssd1 vssd1 vccd1 vccd1 _1743_/A sky130_fd_sc_hd__xnor2_2
XFILLER_7_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1671_ _1699_/B _1671_/B vssd1 vssd1 vccd1 vccd1 _1672_/B sky130_fd_sc_hd__nor2_1
XFILLER_7_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_602 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_613 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_624 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_635 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_646 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_657 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_668 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2223_ _2220_/X _2221_/Y _2177_/X _2178_/Y vssd1 vssd1 vccd1 vccd1 _2224_/C sky130_fd_sc_hd__o211ai_1
XTAP_679 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2154_ _2417_/A _2775_/A vssd1 vssd1 vccd1 vccd1 _2154_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__1630__A _1681_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2085_ _1916_/X _2194_/A _2083_/X _2027_/X _2084_/X vssd1 vssd1 vccd1 vccd1 _2086_/B
+ sky130_fd_sc_hd__a221o_2
XFILLER_61_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2987_ _2987_/A _2987_/B vssd1 vssd1 vccd1 vccd1 _2991_/A sky130_fd_sc_hd__xnor2_1
XFILLER_21_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1938_ _2205_/A vssd1 vssd1 vccd1 vccd1 _2478_/A sky130_fd_sc_hd__buf_4
X_1869_ _1869_/A _1870_/B vssd1 vssd1 vccd1 vccd1 _1903_/A sky130_fd_sc_hd__and2_1
XFILLER_1_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1683__A2 _1597_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2546__A _2546_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2910_ _2886_/A _2886_/B _2909_/X vssd1 vssd1 vccd1 vccd1 _2943_/A sky130_fd_sc_hd__o21a_1
XFILLER_50_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3042__136 vssd1 vssd1 vccd1 vccd1 _3042__136/HI io_out[2] sky130_fd_sc_hd__conb_1
X_2841_ _2843_/A _2843_/B _2843_/C vssd1 vssd1 vccd1 vccd1 _2842_/A sky130_fd_sc_hd__a21o_1
XANTENNA__2712__C _2712_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2772_ _2772_/A vssd1 vssd1 vccd1 vccd1 _2772_/X sky130_fd_sc_hd__buf_2
X_1723_ _1723_/A _1723_/B vssd1 vssd1 vccd1 vccd1 _1723_/Y sky130_fd_sc_hd__nand2_1
XANTENNA__2396__B1 _2919_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1654_ _1657_/B _1654_/B vssd1 vssd1 vccd1 vccd1 _1654_/Y sky130_fd_sc_hd__xnor2_1
X_1585_ _1663_/A _1586_/B vssd1 vssd1 vccd1 vccd1 _1629_/B sky130_fd_sc_hd__and2_1
XTAP_410 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_421 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_432 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_443 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_454 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_465 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_476 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2206_ _2206_/A _2206_/B vssd1 vssd1 vccd1 vccd1 _2557_/A sky130_fd_sc_hd__and2_2
XTAP_487 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_498 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2137_ _2137_/A _2188_/A vssd1 vssd1 vccd1 vccd1 _2139_/A sky130_fd_sc_hd__nand2_1
XFILLER_26_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2068_ _2068_/A vssd1 vssd1 vccd1 vccd1 _2127_/A sky130_fd_sc_hd__inv_2
XFILLER_26_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1656__A2 _1613_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2081__A2 _2023_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2824_ _2824_/A _2824_/B _2824_/C vssd1 vssd1 vccd1 vccd1 _2825_/D sky130_fd_sc_hd__and3_1
X_2755_ _2755_/A _2755_/B _2755_/C vssd1 vssd1 vccd1 vccd1 _2762_/B sky130_fd_sc_hd__nand3_2
X_1706_ _1707_/A _1707_/B vssd1 vssd1 vccd1 vccd1 _1738_/A sky130_fd_sc_hd__nand2_1
X_2686_ _2686_/A vssd1 vssd1 vccd1 vccd1 _2686_/X sky130_fd_sc_hd__clkbuf_2
X_1637_ _1673_/B _1637_/B vssd1 vssd1 vccd1 vccd1 _1638_/B sky130_fd_sc_hd__xor2_1
XFILLER_59_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3170__264 vssd1 vssd1 vccd1 vccd1 _3170__264/HI la_data_out[121] sky130_fd_sc_hd__conb_1
X_1568_ _2996_/A _2999_/B vssd1 vssd1 vccd1 vccd1 _1568_/X sky130_fd_sc_hd__or2_1
XTAP_251 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_240 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1499_ _2985_/B _1520_/B _2987_/B _2987_/A vssd1 vssd1 vccd1 vccd1 _1523_/B sky130_fd_sc_hd__o2bb2a_1
XTAP_262 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_273 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_284 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_295 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_446 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1583__B2 _2684_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_2_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2824__A _2824_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2543__B _2543_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2540_ _2692_/A _2316_/X _2698_/B _2391_/A vssd1 vssd1 vccd1 vccd1 _2540_/X sky130_fd_sc_hd__a22o_1
XFILLER_5_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1574__A1 _1533_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3154__248 vssd1 vssd1 vccd1 vccd1 _3154__248/HI la_data_out[105] sky130_fd_sc_hd__conb_1
X_2471_ _2747_/A _2539_/A _2470_/X vssd1 vssd1 vccd1 vccd1 _2471_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_5_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3048__142 vssd1 vssd1 vccd1 vccd1 _3048__142/HI io_out[8] sky130_fd_sc_hd__conb_1
XFILLER_36_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2807_ _2807_/A _2807_/B vssd1 vssd1 vccd1 vccd1 _2847_/A sky130_fd_sc_hd__nor2_2
X_2738_ _2738_/A _2738_/B vssd1 vssd1 vccd1 vccd1 _2764_/A sky130_fd_sc_hd__xnor2_1
X_2669_ _2523_/X _2515_/A _2593_/X _2793_/A vssd1 vssd1 vccd1 vccd1 _2669_/X sky130_fd_sc_hd__a211o_1
XFILLER_46_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2819__A _2819_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_560 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1971_ _2130_/A _2410_/A _1968_/X _1970_/Y vssd1 vssd1 vccd1 vccd1 _2009_/A sky130_fd_sc_hd__a211o_2
XFILLER_60_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2523_ _2523_/A _2523_/B vssd1 vssd1 vccd1 vccd1 _2523_/X sky130_fd_sc_hd__or2_2
X_2454_ _2454_/A _2454_/B _2629_/B vssd1 vssd1 vccd1 vccd1 _2454_/X sky130_fd_sc_hd__and3_1
X_2385_ _2385_/A vssd1 vssd1 vccd1 vccd1 _2740_/A sky130_fd_sc_hd__buf_2
XFILLER_56_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput1 la_data_in[0] vssd1 vssd1 vccd1 vccd1 input1/X sky130_fd_sc_hd__clkbuf_2
XFILLER_64_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3176__270 vssd1 vssd1 vccd1 vccd1 _3176__270/HI la_data_out[127] sky130_fd_sc_hd__conb_1
XFILLER_10_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_817 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_806 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_839 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_828 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2170_ _2170_/A _2170_/B vssd1 vssd1 vccd1 vccd1 _2242_/B sky130_fd_sc_hd__xnor2_1
XFILLER_38_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_61_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1954_ _2053_/A _1954_/B vssd1 vssd1 vccd1 vccd1 _2008_/B sky130_fd_sc_hd__xor2_2
X_1885_ _1924_/A _1926_/A vssd1 vssd1 vccd1 vccd1 _1887_/A sky130_fd_sc_hd__xnor2_2
X_2506_ _2527_/A _2527_/B vssd1 vssd1 vccd1 vccd1 _2524_/B sky130_fd_sc_hd__xor2_1
X_2437_ _2437_/A _2437_/B vssd1 vssd1 vccd1 vccd1 _2510_/A sky130_fd_sc_hd__xnor2_1
XFILLER_56_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2368_ _2369_/A _2369_/B vssd1 vssd1 vccd1 vccd1 _2370_/A sky130_fd_sc_hd__and2_1
XFILLER_29_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2299_ _2299_/A _2299_/B vssd1 vssd1 vccd1 vccd1 _2299_/X sky130_fd_sc_hd__or2_1
XFILLER_29_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2369__A _2369_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2088__B _2088_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input28_A la_data_in[34] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1720__B _1720_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_7 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1670_ _1699_/B _1671_/B vssd1 vssd1 vccd1 vccd1 _1697_/B sky130_fd_sc_hd__and2_1
XFILLER_7_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_603 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_614 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_625 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2279__A _2501_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_636 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_647 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_658 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2222_ _2177_/X _2178_/Y _2220_/X _2221_/Y vssd1 vssd1 vccd1 vccd1 _2289_/A sky130_fd_sc_hd__a211o_1
XTAP_669 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2153_ _2209_/A _2153_/B vssd1 vssd1 vccd1 vccd1 _2159_/A sky130_fd_sc_hd__xnor2_1
XFILLER_26_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2084_ _1968_/C _2028_/A _2142_/A _1919_/C vssd1 vssd1 vccd1 vccd1 _2084_/X sky130_fd_sc_hd__a22o_1
XANTENNA__1989__B2 _1939_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_21_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2986_ _2986_/A _2986_/B vssd1 vssd1 vccd1 vccd1 _2987_/B sky130_fd_sc_hd__xnor2_1
X_1937_ _1937_/A _1993_/B vssd1 vssd1 vccd1 vccd1 _1952_/A sky130_fd_sc_hd__xnor2_2
X_1868_ _1869_/A _1870_/A _1870_/B vssd1 vssd1 vccd1 vccd1 _1871_/A sky130_fd_sc_hd__nor3_1
X_1799_ _1816_/A _1939_/A _1796_/X _1798_/Y vssd1 vssd1 vccd1 vccd1 _1839_/A sky130_fd_sc_hd__a211o_1
XFILLER_57_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2636__B _2636_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3081__175 vssd1 vssd1 vccd1 vccd1 _3081__175/HI la_data_out[0] sky130_fd_sc_hd__conb_1
X_2840_ _2840_/A _2840_/B vssd1 vssd1 vccd1 vccd1 _2843_/C sky130_fd_sc_hd__nor2_1
XANTENNA__2396__A1 _2393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2771_ _2683_/A _2683_/B _2770_/X vssd1 vssd1 vccd1 vccd1 _2807_/A sky130_fd_sc_hd__a21oi_2
XFILLER_7_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1722_ _1722_/A vssd1 vssd1 vccd1 vccd1 _1722_/Y sky130_fd_sc_hd__inv_2
X_1653_ _1613_/A _1613_/B _1620_/A vssd1 vssd1 vccd1 vccd1 _1654_/B sky130_fd_sc_hd__a21o_1
X_1584_ _2939_/A _1584_/B vssd1 vssd1 vccd1 vccd1 _1586_/B sky130_fd_sc_hd__xnor2_1
XTAP_400 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_411 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_422 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_433 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_444 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_455 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_466 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2205_ _2205_/A _2205_/B vssd1 vssd1 vccd1 vccd1 _2210_/A sky130_fd_sc_hd__xnor2_2
XTAP_477 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_488 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_499 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2737__A _2737_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2136_ _2130_/X _2552_/A _2134_/X _2135_/Y vssd1 vssd1 vccd1 vccd1 _2179_/A sky130_fd_sc_hd__a211o_2
X_2067_ _2051_/A _2067_/B vssd1 vssd1 vccd1 vccd1 _2068_/A sky130_fd_sc_hd__and2b_1
XFILLER_22_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2969_ _2970_/A _2970_/B _2970_/C vssd1 vssd1 vccd1 vccd1 _2971_/A sky130_fd_sc_hd__o21ai_4
XFILLER_1_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3065__159 vssd1 vssd1 vccd1 vccd1 _3065__159/HI io_out[25] sky130_fd_sc_hd__conb_1
XFILLER_60_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_591 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2276__B input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2823_ _2824_/B _2824_/C _2976_/A vssd1 vssd1 vccd1 vccd1 _2825_/C sky130_fd_sc_hd__a21oi_2
X_2754_ _2755_/B _2755_/C _2755_/A vssd1 vssd1 vccd1 vccd1 _2843_/A sky130_fd_sc_hd__a21o_2
X_1705_ _1675_/A _1675_/B _1701_/B _1673_/B vssd1 vssd1 vccd1 vccd1 _1707_/B sky130_fd_sc_hd__a22o_1
X_2685_ _2685_/A vssd1 vssd1 vccd1 vccd1 _2934_/A sky130_fd_sc_hd__clkbuf_2
X_1636_ _2920_/A _1636_/B vssd1 vssd1 vccd1 vccd1 _1637_/B sky130_fd_sc_hd__and2_1
X_1567_ _1649_/A _1567_/B vssd1 vssd1 vccd1 vccd1 _1571_/A sky130_fd_sc_hd__or2_2
XFILLER_59_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_241 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_230 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1498_ _2988_/A _2986_/A vssd1 vssd1 vccd1 vccd1 _1520_/B sky130_fd_sc_hd__nor2_1
XTAP_252 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_263 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_274 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_296 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_285 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2119_ _2120_/A _2120_/B vssd1 vssd1 vccd1 vccd1 _2121_/A sky130_fd_sc_hd__and2_1
XFILLER_27_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input10_A la_data_in[18] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2543__C _2543_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1574__A2 _1533_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3193__287 vssd1 vssd1 vccd1 vccd1 _3193__287/HI wbs_dat_o[15] sky130_fd_sc_hd__conb_1
X_2470_ _2391_/A _2316_/X _2698_/B _2385_/A vssd1 vssd1 vccd1 vccd1 _2470_/X sky130_fd_sc_hd__a22o_1
XFILLER_64_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3087__181 vssd1 vssd1 vccd1 vccd1 _3087__181/HI la_data_out[6] sky130_fd_sc_hd__conb_1
XFILLER_63_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2806_ _2783_/A _2783_/C _2783_/B vssd1 vssd1 vccd1 vccd1 _2857_/B sky130_fd_sc_hd__o21bai_2
X_2737_ _2737_/A _2877_/A vssd1 vssd1 vccd1 vccd1 _2738_/B sky130_fd_sc_hd__nor2_1
X_2668_ _2668_/A _2668_/B vssd1 vssd1 vccd1 vccd1 _2668_/Y sky130_fd_sc_hd__xnor2_2
X_1619_ _1618_/B _1657_/A vssd1 vssd1 vccd1 vccd1 _1620_/B sky130_fd_sc_hd__and2b_1
X_2599_ _2599_/A _2599_/B vssd1 vssd1 vccd1 vccd1 _2602_/A sky130_fd_sc_hd__nor2_2
XANTENNA_input2_A la_data_in[10] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input58_A la_data_in[61] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1723__B _1723_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_1_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1492__A1 _1488_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1970_ _2181_/A _2416_/A _2181_/B vssd1 vssd1 vccd1 vccd1 _1970_/Y sky130_fd_sc_hd__a21oi_1
X_3121__215 vssd1 vssd1 vccd1 vccd1 _3121__215/HI la_data_out[40] sky130_fd_sc_hd__conb_1
XFILLER_41_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2522_ _2522_/A _2522_/B vssd1 vssd1 vccd1 vccd1 _2522_/Y sky130_fd_sc_hd__xnor2_2
XFILLER_5_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2453_ _2425_/B _2425_/C _2425_/A vssd1 vssd1 vccd1 vccd1 _2526_/A sky130_fd_sc_hd__a21boi_1
X_2384_ _2538_/A _2979_/A _2979_/B vssd1 vssd1 vccd1 vccd1 _2390_/B sky130_fd_sc_hd__or3_1
Xinput2 la_data_in[10] vssd1 vssd1 vccd1 vccd1 input2/X sky130_fd_sc_hd__buf_2
XFILLER_28_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2464__B _2464_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2735__A1 _2919_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_524 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_535 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_807 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_829 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_818 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1953_ _1953_/A _1953_/B vssd1 vssd1 vccd1 vccd1 _1954_/B sky130_fd_sc_hd__nand2_1
X_3199__293 vssd1 vssd1 vccd1 vccd1 _3199__293/HI wbs_dat_o[21] sky130_fd_sc_hd__conb_1
X_1884_ _1884_/A _1884_/B vssd1 vssd1 vccd1 vccd1 _2027_/A sky130_fd_sc_hd__and2_1
X_2505_ _2589_/A _2505_/B vssd1 vssd1 vccd1 vccd1 _2527_/B sky130_fd_sc_hd__and2_1
X_2436_ _2525_/A _2436_/B vssd1 vssd1 vccd1 vccd1 _2437_/B sky130_fd_sc_hd__nor2_1
X_2367_ _2367_/A _2367_/B vssd1 vssd1 vccd1 vccd1 _2369_/B sky130_fd_sc_hd__xnor2_1
X_2298_ _2299_/A _2299_/B vssd1 vssd1 vccd1 vccd1 _2300_/A sky130_fd_sc_hd__and2_1
XANTENNA__2475__A _2528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_8 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_604 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_615 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2221_ _2220_/A _2220_/B _2220_/C vssd1 vssd1 vccd1 vccd1 _2221_/Y sky130_fd_sc_hd__a21oi_1
XTAP_626 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_637 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_648 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_659 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2152_ _1984_/A _2411_/A _2558_/A _1807_/A _2151_/X vssd1 vssd1 vccd1 vccd1 _2153_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_38_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2083_ _2083_/A _2083_/B vssd1 vssd1 vccd1 vccd1 _2083_/X sky130_fd_sc_hd__xor2_4
XFILLER_38_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3127__221 vssd1 vssd1 vccd1 vccd1 _3127__221/HI la_data_out[46] sky130_fd_sc_hd__conb_1
XFILLER_22_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2985_ _2988_/A _2985_/B vssd1 vssd1 vccd1 vccd1 _2986_/B sky130_fd_sc_hd__nor2_1
X_1936_ _2205_/A _1883_/B _1895_/B vssd1 vssd1 vccd1 vccd1 _1993_/B sky130_fd_sc_hd__o21ai_2
X_1867_ _1895_/A _1867_/B vssd1 vssd1 vccd1 vccd1 _1870_/B sky130_fd_sc_hd__nor2_1
Xinput60 la_data_in[63] vssd1 vssd1 vccd1 vccd1 _1759_/A sky130_fd_sc_hd__buf_2
X_1798_ _1821_/A _1817_/A _1968_/B vssd1 vssd1 vccd1 vccd1 _1798_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_29_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2419_ _2739_/A _2965_/A vssd1 vssd1 vccd1 vccd1 _2419_/Y sky130_fd_sc_hd__nor2_1
XFILLER_29_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2636__C _2636_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input40_A la_data_in[45] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2843__A _2843_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2770_ _2690_/A _2770_/B vssd1 vssd1 vccd1 vccd1 _2770_/X sky130_fd_sc_hd__and2b_1
X_1721_ _1721_/A _1749_/A vssd1 vssd1 vccd1 vccd1 _1725_/A sky130_fd_sc_hd__or2_1
X_1652_ _1655_/A _1655_/B vssd1 vssd1 vccd1 vccd1 _1657_/B sky130_fd_sc_hd__xnor2_1
XFILLER_7_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1583_ _1514_/X _2930_/X _2973_/Y _2684_/X _1582_/X vssd1 vssd1 vccd1 vccd1 _1584_/B
+ sky130_fd_sc_hd__a221o_1
XTAP_401 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_412 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_423 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_434 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_445 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_456 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_467 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2204_ _2568_/A _1987_/A _2026_/Y _2037_/A _2203_/X vssd1 vssd1 vccd1 vccd1 _2205_/B
+ sky130_fd_sc_hd__a221o_1
XTAP_478 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_489 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2135_ _2313_/S _2134_/C _2310_/A vssd1 vssd1 vccd1 vccd1 _2135_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_39_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2066_ _2112_/B _2066_/B vssd1 vssd1 vccd1 vccd1 _2125_/A sky130_fd_sc_hd__or2_1
XFILLER_22_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2968_ _2913_/A _2772_/X _2965_/Y _2967_/X vssd1 vssd1 vccd1 vccd1 _2970_/C sky130_fd_sc_hd__a211o_1
X_1919_ _1968_/A _2013_/B _1919_/C vssd1 vssd1 vccd1 vccd1 _1919_/X sky130_fd_sc_hd__and3_1
X_2899_ _2899_/A _2899_/B vssd1 vssd1 vccd1 vccd1 _2958_/B sky130_fd_sc_hd__xor2_4
XFILLER_57_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1889__A1 _1979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2822_ _2936_/A _2820_/X _2821_/X vssd1 vssd1 vccd1 vccd1 _2824_/C sky130_fd_sc_hd__a21oi_1
XFILLER_31_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2753_ _2976_/A _2753_/B vssd1 vssd1 vccd1 vccd1 _2755_/A sky130_fd_sc_hd__xnor2_1
X_1704_ _1704_/A _1704_/B vssd1 vssd1 vccd1 vccd1 _1707_/A sky130_fd_sc_hd__nor2_1
XANTENNA__1917__A _2023_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2684_ _2684_/A vssd1 vssd1 vccd1 vccd1 _2684_/X sky130_fd_sc_hd__clkbuf_2
X_1635_ _1663_/A _1635_/B vssd1 vssd1 vccd1 vccd1 _1673_/B sky130_fd_sc_hd__xor2_2
X_1566_ _1566_/A _1577_/B vssd1 vssd1 vccd1 vccd1 _1567_/B sky130_fd_sc_hd__nor2_1
XTAP_242 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_231 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_220 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1497_ _2992_/A _2992_/B vssd1 vssd1 vccd1 vccd1 _1527_/B sky130_fd_sc_hd__and2_1
XTAP_253 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_264 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_275 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_297 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_286 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2118_ _2118_/A _2118_/B vssd1 vssd1 vccd1 vccd1 _2120_/B sky130_fd_sc_hd__xnor2_1
XFILLER_27_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2049_ _2049_/A _2049_/B vssd1 vssd1 vccd1 vccd1 _2049_/Y sky130_fd_sc_hd__nor2_1
XFILLER_42_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_22_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3032__126 vssd1 vssd1 vccd1 vccd1 _3032__126/HI io_oeb[29] sky130_fd_sc_hd__conb_1
XFILLER_1_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_33_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2393__A _2393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2568__A _2568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2805_ _2805_/A _2805_/B vssd1 vssd1 vccd1 vccd1 _2850_/A sky130_fd_sc_hd__nor2_1
X_2736_ _2919_/A _2919_/B vssd1 vssd1 vccd1 vccd1 _2877_/A sky130_fd_sc_hd__nor2_2
X_2667_ _2602_/A _2602_/B _2599_/A vssd1 vssd1 vccd1 vccd1 _2668_/B sky130_fd_sc_hd__a21oi_1
X_1618_ _1657_/A _1618_/B vssd1 vssd1 vccd1 vccd1 _1620_/A sky130_fd_sc_hd__and2b_1
X_2598_ _2597_/B _2597_/C _2597_/A vssd1 vssd1 vccd1 vccd1 _2599_/B sky130_fd_sc_hd__a21oi_1
X_1549_ _2932_/A _2921_/X vssd1 vssd1 vccd1 vccd1 _1549_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__2197__B _2197_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1557__A _1557_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_40_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_37_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1492__A2 _1488_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3160__254 vssd1 vssd1 vccd1 vccd1 _3160__254/HI la_data_out[111] sky130_fd_sc_hd__conb_1
X_3201__295 vssd1 vssd1 vccd1 vccd1 _3201__295/HI wbs_dat_o[23] sky130_fd_sc_hd__conb_1
X_2521_ _2521_/A _2521_/B vssd1 vssd1 vccd1 vccd1 _2522_/B sky130_fd_sc_hd__nand2_1
X_2452_ _2429_/B _2437_/B _2427_/X vssd1 vssd1 vccd1 vccd1 _2524_/A sky130_fd_sc_hd__a21o_1
XFILLER_46_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2383_ _2462_/A _2931_/A _2383_/C vssd1 vssd1 vccd1 vccd1 _2979_/B sky130_fd_sc_hd__and3_1
XANTENNA__1499__A1_N _2985_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput3 la_data_in[11] vssd1 vssd1 vccd1 vccd1 input3/X sky130_fd_sc_hd__clkbuf_2
XFILLER_64_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2680__A1 _2608_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2719_ _2719_/A _2791_/A vssd1 vssd1 vccd1 vccd1 _2719_/Y sky130_fd_sc_hd__nor2_1
XANTENNA__2499__A1 input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3144__238 vssd1 vssd1 vccd1 vccd1 _3144__238/HI la_data_out[63] sky130_fd_sc_hd__conb_1
XFILLER_15_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3038__132 vssd1 vssd1 vccd1 vccd1 _3038__132/HI io_oeb[35] sky130_fd_sc_hd__conb_1
XTAP_808 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_819 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1952_ _1952_/A _1952_/B vssd1 vssd1 vccd1 vccd1 _2053_/A sky130_fd_sc_hd__xnor2_2
X_1883_ _2612_/A _1883_/B vssd1 vssd1 vccd1 vccd1 _1893_/A sky130_fd_sc_hd__xnor2_1
X_2504_ _2504_/A _2504_/B _2504_/C vssd1 vssd1 vccd1 vccd1 _2505_/B sky130_fd_sc_hd__or3_1
X_2435_ _2434_/A _2647_/B _2434_/B vssd1 vssd1 vccd1 vccd1 _2436_/B sky130_fd_sc_hd__a21oi_1
X_2366_ _2306_/Y _2364_/X _2444_/A vssd1 vssd1 vccd1 vccd1 _2367_/B sky130_fd_sc_hd__o21a_1
XFILLER_29_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2297_ _2294_/A _2294_/Y _2297_/S vssd1 vssd1 vccd1 vccd1 _2299_/B sky130_fd_sc_hd__mux2_1
XFILLER_37_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1695__A2 _2973_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2666__A _2725_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_605 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_616 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2220_ _2220_/A _2220_/B _2220_/C vssd1 vssd1 vccd1 vccd1 _2220_/X sky130_fd_sc_hd__and3_1
XTAP_627 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_638 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_649 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2883__A1 _2884_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2151_ _1859_/Y _2335_/A _2099_/A _1939_/A vssd1 vssd1 vccd1 vccd1 _2151_/X sky130_fd_sc_hd__a2bb2o_1
XFILLER_38_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2082_ _1977_/A _1977_/B _2026_/A _2081_/X vssd1 vssd1 vccd1 vccd1 _2083_/B sky130_fd_sc_hd__a31o_2
XFILLER_19_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3166__260 vssd1 vssd1 vccd1 vccd1 _3166__260/HI la_data_out[117] sky130_fd_sc_hd__conb_1
XFILLER_19_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2635__A1 _2636_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2984_ _2984_/A _2984_/B vssd1 vssd1 vccd1 vccd1 _2986_/A sky130_fd_sc_hd__xnor2_4
XFILLER_21_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1935_ _2266_/A vssd1 vssd1 vccd1 vccd1 _2205_/A sky130_fd_sc_hd__buf_2
XFILLER_21_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1866_ _1865_/B _1865_/C _1865_/A vssd1 vssd1 vccd1 vccd1 _1867_/B sky130_fd_sc_hd__a21oi_1
Xinput61 la_data_in[6] vssd1 vssd1 vccd1 vccd1 _1944_/B sky130_fd_sc_hd__buf_2
Xinput50 la_data_in[54] vssd1 vssd1 vccd1 vccd1 _2954_/A sky130_fd_sc_hd__buf_2
X_1797_ _1879_/B vssd1 vssd1 vccd1 vccd1 _1968_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_1_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2418_ _2418_/A _2418_/B vssd1 vssd1 vccd1 vccd1 _2965_/A sky130_fd_sc_hd__or2_4
X_2349_ _2406_/B _2349_/B vssd1 vssd1 vccd1 vccd1 _2483_/A sky130_fd_sc_hd__and2_1
XFILLER_29_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_476 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3002__304 vssd1 vssd1 vccd1 vccd1 io_out[0] _3002__304/LO sky130_fd_sc_hd__conb_1
XANTENNA__1549__B _2921_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input33_A la_data_in[39] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2865__A1 _2258_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_63_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2617__A1 _2819_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1720_ _1720_/A _1720_/B vssd1 vssd1 vccd1 vccd1 _1749_/A sky130_fd_sc_hd__nor2_1
X_1651_ _1651_/A _1651_/B vssd1 vssd1 vccd1 vccd1 _1655_/B sky130_fd_sc_hd__xor2_4
X_1582_ _2927_/A _2934_/X _2935_/X _2922_/X vssd1 vssd1 vccd1 vccd1 _1582_/X sky130_fd_sc_hd__a22o_1
XTAP_402 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_413 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_424 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_435 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_446 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_457 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2203_ _1919_/C _1942_/A _1946_/A _1916_/X vssd1 vssd1 vccd1 vccd1 _2203_/X sky130_fd_sc_hd__a22o_1
XTAP_468 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_479 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2134_ _2313_/S _2134_/B _2134_/C vssd1 vssd1 vccd1 vccd1 _2134_/X sky130_fd_sc_hd__and3_1
XFILLER_54_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2065_ _2057_/A _2063_/Y _2064_/X vssd1 vssd1 vccd1 vccd1 _2118_/A sky130_fd_sc_hd__a21bo_1
XFILLER_19_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2967_ _2863_/X _2773_/X _2966_/X _2758_/X vssd1 vssd1 vccd1 vccd1 _2967_/X sky130_fd_sc_hd__a22o_1
X_1918_ _2079_/A vssd1 vssd1 vccd1 vccd1 _1919_/C sky130_fd_sc_hd__clkbuf_2
X_2898_ _2898_/A _3001_/A vssd1 vssd1 vccd1 vccd1 _2899_/B sky130_fd_sc_hd__nand2_1
X_1849_ _1837_/A _1849_/B vssd1 vssd1 vccd1 vccd1 _1869_/A sky130_fd_sc_hd__and2b_1
XFILLER_1_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1510__A1 _2557_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2821_ _2740_/A _2748_/X _2749_/A _2933_/A vssd1 vssd1 vccd1 vccd1 _2821_/X sky130_fd_sc_hd__a22o_1
X_2752_ _2752_/A _2752_/B vssd1 vssd1 vccd1 vccd1 _2753_/B sky130_fd_sc_hd__nor2_1
X_1703_ _1703_/A _1703_/B vssd1 vssd1 vccd1 vccd1 _1704_/B sky130_fd_sc_hd__and2_1
XFILLER_8_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2683_ _2683_/A _2683_/B vssd1 vssd1 vccd1 vccd1 _2690_/A sky130_fd_sc_hd__xnor2_1
X_1634_ _2983_/A _1634_/B vssd1 vssd1 vccd1 vccd1 _1635_/B sky130_fd_sc_hd__xnor2_2
X_1565_ _1566_/A _1577_/B vssd1 vssd1 vccd1 vccd1 _1649_/A sky130_fd_sc_hd__and2_1
XTAP_232 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_221 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_210 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1933__A _1965_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1496_ _2991_/A _2991_/B vssd1 vssd1 vccd1 vccd1 _1527_/A sky130_fd_sc_hd__nor2_1
XTAP_254 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1652__B _1655_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_243 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_265 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_276 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_298 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_287 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2117_ _2125_/A _2125_/B vssd1 vssd1 vccd1 vccd1 _2118_/B sky130_fd_sc_hd__xnor2_1
XFILLER_54_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2048_ _2048_/A _2048_/B vssd1 vssd1 vccd1 vccd1 _2051_/A sky130_fd_sc_hd__xnor2_1
XFILLER_50_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2517__B1 _2518_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2939__A _2939_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3071__165 vssd1 vssd1 vccd1 vccd1 _3071__165/HI io_out[31] sky130_fd_sc_hd__conb_1
XFILLER_49_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3206__300 vssd1 vssd1 vccd1 vccd1 _3206__300/HI wbs_dat_o[28] sky130_fd_sc_hd__conb_1
XFILLER_51_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2804_ _2804_/A _2905_/A vssd1 vssd1 vccd1 vccd1 _2852_/A sky130_fd_sc_hd__nand2_2
X_2735_ _2919_/A _2919_/B _2810_/A _2811_/C vssd1 vssd1 vccd1 vccd1 _2737_/A sky130_fd_sc_hd__a22o_2
X_2666_ _2725_/A _2725_/B vssd1 vssd1 vccd1 vccd1 _2668_/A sky130_fd_sc_hd__xor2_2
X_3055__149 vssd1 vssd1 vccd1 vccd1 _3055__149/HI io_out[15] sky130_fd_sc_hd__conb_1
X_1617_ _1573_/B _1614_/Y _1615_/X _1616_/X vssd1 vssd1 vccd1 vccd1 _1618_/B sky130_fd_sc_hd__a22o_1
X_2597_ _2597_/A _2597_/B _2597_/C vssd1 vssd1 vccd1 vccd1 _2599_/A sky130_fd_sc_hd__and3_1
X_1548_ _2977_/A _1548_/B vssd1 vssd1 vccd1 vccd1 _1554_/A sky130_fd_sc_hd__xnor2_2
XFILLER_59_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2941__B _2985_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_45_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2520_ _2371_/A _2369_/X _2446_/X _2370_/A vssd1 vssd1 vccd1 vccd1 _2521_/B sky130_fd_sc_hd__a211o_1
X_2451_ _2451_/A _2451_/B vssd1 vssd1 vccd1 vccd1 _2523_/A sky130_fd_sc_hd__nand2_1
XANTENNA__2579__A _2978_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2382_ _2462_/A _2931_/A _2383_/C vssd1 vssd1 vccd1 vccd1 _2979_/A sky130_fd_sc_hd__a21oi_2
XFILLER_39_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput4 la_data_in[12] vssd1 vssd1 vccd1 vccd1 input4/X sky130_fd_sc_hd__clkbuf_4
XFILLER_37_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_452 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_51_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2196__A1 _2416_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2718_ _2718_/A _2791_/A vssd1 vssd1 vccd1 vccd1 _2793_/B sky130_fd_sc_hd__and2_1
XFILLER_10_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2649_ _2649_/A _2649_/B vssd1 vssd1 vccd1 vccd1 _2651_/C sky130_fd_sc_hd__or2_1
XFILLER_59_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3183__277 vssd1 vssd1 vccd1 vccd1 _3183__277/HI wbs_dat_o[5] sky130_fd_sc_hd__conb_1
XFILLER_35_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3077__171 vssd1 vssd1 vccd1 vccd1 _3077__171/HI io_out[37] sky130_fd_sc_hd__conb_1
XANTENNA_input63_A la_data_in[8] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_809 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1951_ _2478_/A _1951_/B vssd1 vssd1 vccd1 vccd1 _1952_/B sky130_fd_sc_hd__xnor2_2
X_1882_ _1816_/A _2020_/A _1879_/X _1881_/Y vssd1 vssd1 vccd1 vccd1 _1883_/B sky130_fd_sc_hd__a211o_2
X_2503_ _2504_/A _2504_/B _2504_/C vssd1 vssd1 vccd1 vccd1 _2589_/A sky130_fd_sc_hd__o21ai_4
X_2434_ _2434_/A _2434_/B _2647_/B vssd1 vssd1 vccd1 vccd1 _2525_/A sky130_fd_sc_hd__and3_2
X_2365_ _2365_/A _2450_/B vssd1 vssd1 vccd1 vccd1 _2444_/A sky130_fd_sc_hd__or2_1
XFILLER_56_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2296_ _2296_/A _2296_/B vssd1 vssd1 vccd1 vccd1 _2297_/S sky130_fd_sc_hd__nor2_1
XFILLER_52_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_21_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__2012__A _2188_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3111__205 vssd1 vssd1 vccd1 vccd1 _3111__205/HI la_data_out[30] sky130_fd_sc_hd__conb_1
XANTENNA__1851__A _1974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2341__B2 _2416_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_62_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2682__A _2824_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_31_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1745__B _1745_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2580__B2 _2434_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_606 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_617 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_628 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_639 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2150_ _2150_/A vssd1 vssd1 vccd1 vccd1 _2558_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_38_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2081_ _1975_/A _2023_/B _1975_/B vssd1 vssd1 vccd1 vccd1 _2081_/X sky130_fd_sc_hd__o21a_1
XFILLER_19_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2635__A2 _2636_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2983_ _2983_/A _2983_/B vssd1 vssd1 vccd1 vccd1 _2984_/B sky130_fd_sc_hd__xnor2_2
X_1934_ _2043_/A vssd1 vssd1 vccd1 vccd1 _2266_/A sky130_fd_sc_hd__inv_2
X_1865_ _1865_/A _1865_/B _1865_/C vssd1 vssd1 vccd1 vccd1 _1895_/A sky130_fd_sc_hd__and3_1
Xinput40 la_data_in[45] vssd1 vssd1 vccd1 vccd1 _2369_/A sky130_fd_sc_hd__clkbuf_2
Xinput51 la_data_in[55] vssd1 vssd1 vccd1 vccd1 _1488_/A sky130_fd_sc_hd__buf_2
Xinput62 la_data_in[7] vssd1 vssd1 vccd1 vccd1 _2043_/A sky130_fd_sc_hd__buf_2
X_1796_ _1968_/A _2013_/B _1817_/A vssd1 vssd1 vccd1 vccd1 _1796_/X sky130_fd_sc_hd__and3_1
XANTENNA__1655__B _1655_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2417_ _2417_/A vssd1 vssd1 vccd1 vccd1 _2739_/A sky130_fd_sc_hd__buf_2
X_2348_ _2214_/A _2348_/B vssd1 vssd1 vccd1 vccd1 _2349_/B sky130_fd_sc_hd__and2b_1
XFILLER_57_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2279_ _2501_/A _2827_/A vssd1 vssd1 vccd1 vccd1 _2279_/Y sky130_fd_sc_hd__nor2_1
XFILLER_52_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_488 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2151__A1_N _1859_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2562__A1 _2557_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2865__A2 _2684_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input26_A la_data_in[32] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3189__283 vssd1 vssd1 vccd1 vccd1 _3189__283/HI wbs_dat_o[11] sky130_fd_sc_hd__conb_1
XFILLER_35_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2617__A2 _2965_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_16_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1650_ _1567_/B _1610_/B _1649_/Y _1571_/B _1611_/A vssd1 vssd1 vccd1 vccd1 _1651_/B
+ sky130_fd_sc_hd__a221o_4
XFILLER_7_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1581_ _1623_/A _1581_/B vssd1 vssd1 vccd1 vccd1 _1663_/A sky130_fd_sc_hd__nor2_2
XTAP_403 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_414 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_425 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_436 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_447 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_458 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_21_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2202_ _2201_/B _2201_/C _2201_/A vssd1 vssd1 vccd1 vccd1 _2220_/B sky130_fd_sc_hd__o21ai_1
XTAP_469 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2133_ _2321_/A vssd1 vssd1 vccd1 vccd1 _2134_/C sky130_fd_sc_hd__dlymetal6s2s_1
X_2064_ _2064_/A _2064_/B vssd1 vssd1 vccd1 vccd1 _2064_/X sky130_fd_sc_hd__or2_1
XFILLER_19_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2966_ _2966_/A vssd1 vssd1 vccd1 vccd1 _2966_/X sky130_fd_sc_hd__clkbuf_2
X_1917_ _2023_/B vssd1 vssd1 vccd1 vccd1 _2079_/A sky130_fd_sc_hd__clkbuf_2
X_2897_ _2790_/B _2896_/Y _2851_/B vssd1 vssd1 vccd1 vccd1 _3001_/A sky130_fd_sc_hd__o21ba_1
X_1848_ _1848_/A _1848_/B vssd1 vssd1 vccd1 vccd1 _1876_/A sky130_fd_sc_hd__or2_1
X_1779_ _1879_/B vssd1 vssd1 vccd1 vccd1 _2013_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__2497__A input7/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3117__211 vssd1 vssd1 vccd1 vccd1 _3117__211/HI la_data_out[36] sky130_fd_sc_hd__conb_1
XANTENNA__1510__A2 _2871_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_314 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2820_ _2820_/A vssd1 vssd1 vccd1 vccd1 _2820_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2751_ _2557_/X _2931_/A _2931_/B _2820_/A _2863_/A vssd1 vssd1 vccd1 vccd1 _2752_/B
+ sky130_fd_sc_hd__a32o_1
X_1702_ _1703_/A _1703_/B vssd1 vssd1 vccd1 vccd1 _1704_/A sky130_fd_sc_hd__nor2_1
X_2682_ _2824_/A _2682_/B vssd1 vssd1 vccd1 vccd1 _2683_/B sky130_fd_sc_hd__xnor2_1
X_1633_ _2684_/X _2871_/Y _1632_/X vssd1 vssd1 vccd1 vccd1 _1634_/B sky130_fd_sc_hd__a21oi_1
XFILLER_8_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1564_ _1610_/A _1564_/B vssd1 vssd1 vccd1 vccd1 _1577_/B sky130_fd_sc_hd__or2_1
XTAP_233 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_222 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_211 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_200 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1495_ _2952_/A _3000_/B _2999_/A _1494_/X vssd1 vssd1 vccd1 vccd1 _1532_/A sky130_fd_sc_hd__o31ai_4
XTAP_255 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_244 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_266 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_277 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_299 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_288 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2116_ _2116_/A _2116_/B vssd1 vssd1 vccd1 vccd1 _2125_/B sky130_fd_sc_hd__or2_1
XFILLER_39_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2047_ _2069_/A _2070_/B vssd1 vssd1 vccd1 vccd1 _2048_/B sky130_fd_sc_hd__xnor2_1
XFILLER_35_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2949_ _2949_/A vssd1 vssd1 vccd1 vccd1 _2950_/A sky130_fd_sc_hd__inv_2
XFILLER_1_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_32_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2803_ _2719_/A _2791_/A _2789_/B _2790_/B vssd1 vssd1 vccd1 vccd1 _2905_/A sky130_fd_sc_hd__o31a_1
X_2734_ _2703_/A _2703_/B _2766_/A vssd1 vssd1 vccd1 vccd1 _2738_/A sky130_fd_sc_hd__a21o_1
XFILLER_8_292 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2665_ _2665_/A _2665_/B vssd1 vssd1 vccd1 vccd1 _2725_/B sky130_fd_sc_hd__xnor2_2
X_1616_ _1616_/A _1616_/B vssd1 vssd1 vccd1 vccd1 _1616_/X sky130_fd_sc_hd__or2_1
X_3094__188 vssd1 vssd1 vccd1 vccd1 _3094__188/HI la_data_out[13] sky130_fd_sc_hd__conb_1
X_2596_ _2593_/X _2603_/A _2523_/X _2518_/B vssd1 vssd1 vccd1 vccd1 _2597_/C sky130_fd_sc_hd__o211ai_1
XANTENNA__1970__A2 _2416_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1547_ _2926_/A _2097_/B _1547_/S vssd1 vssd1 vccd1 vccd1 _1548_/B sky130_fd_sc_hd__mux2_2
XANTENNA__2775__A _2775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_27_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_24_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_623 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_61_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_575 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2450_ _2450_/A _2450_/B _2451_/B vssd1 vssd1 vccd1 vccd1 _2450_/X sky130_fd_sc_hd__or3b_1
XANTENNA__2579__B input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2381_ _2462_/B _2458_/C vssd1 vssd1 vccd1 vccd1 _2383_/C sky130_fd_sc_hd__nand2_1
Xinput5 la_data_in[13] vssd1 vssd1 vccd1 vccd1 input5/X sky130_fd_sc_hd__clkbuf_4
XFILLER_36_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1939__A _1939_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3022__116 vssd1 vssd1 vccd1 vccd1 _3022__116/HI io_oeb[19] sky130_fd_sc_hd__conb_1
XFILLER_20_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2717_ _2731_/A _2731_/B vssd1 vssd1 vccd1 vccd1 _2791_/A sky130_fd_sc_hd__xnor2_2
X_2648_ _1888_/B _2880_/A _2496_/A _2402_/X vssd1 vssd1 vccd1 vccd1 _2649_/B sky130_fd_sc_hd__a22o_1
X_2579_ _2978_/A input6/X _2647_/A vssd1 vssd1 vccd1 vccd1 _2774_/A sky130_fd_sc_hd__and3_1
XFILLER_59_214 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_59_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1584__A _2939_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input56_A la_data_in[5] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1759__A _1759_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1950_ _2273_/A _2549_/A _2550_/A _1807_/A _1949_/Y vssd1 vssd1 vccd1 vccd1 _1951_/B
+ sky130_fd_sc_hd__a221o_1
X_1881_ _2013_/A _2337_/A _2013_/B vssd1 vssd1 vccd1 vccd1 _1881_/Y sky130_fd_sc_hd__a21oi_1
X_2502_ _2273_/X _2913_/B _2578_/A _2434_/A _2501_/Y vssd1 vssd1 vccd1 vccd1 _2504_/C
+ sky130_fd_sc_hd__a221o_2
XFILLER_51_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2433_ _2433_/A vssd1 vssd1 vccd1 vccd1 _2647_/B sky130_fd_sc_hd__clkbuf_2
X_2364_ _2450_/A _2450_/B vssd1 vssd1 vccd1 vccd1 _2364_/X sky130_fd_sc_hd__xor2_2
X_2295_ _2170_/A _2235_/X _2234_/A _2236_/X vssd1 vssd1 vccd1 vccd1 _2296_/B sky130_fd_sc_hd__a211oi_2
XFILLER_56_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_431 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2638__B1 _2766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_52_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3150__244 vssd1 vssd1 vccd1 vccd1 _3150__244/HI la_data_out[101] sky130_fd_sc_hd__conb_1
XFILLER_46_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1579__A _2818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_607 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_618 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_629 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2080_ _2187_/A _2187_/B vssd1 vssd1 vccd1 vccd1 _2083_/A sky130_fd_sc_hd__nor2_2
XFILLER_34_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2982_ _2932_/A _2979_/X _2981_/Y vssd1 vssd1 vccd1 vccd1 _2983_/B sky130_fd_sc_hd__o21a_1
XFILLER_21_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1933_ _1965_/A _1933_/B vssd1 vssd1 vccd1 vccd1 _1937_/A sky130_fd_sc_hd__xor2_2
X_1864_ _1981_/A _1864_/B _1864_/C vssd1 vssd1 vccd1 vccd1 _1865_/C sky130_fd_sc_hd__or3_1
Xinput30 la_data_in[36] vssd1 vssd1 vccd1 vccd1 _1873_/A sky130_fd_sc_hd__clkbuf_1
X_1795_ _1924_/A vssd1 vssd1 vccd1 vccd1 _1817_/A sky130_fd_sc_hd__clkbuf_2
Xinput52 la_data_in[56] vssd1 vssd1 vccd1 vccd1 _1533_/A sky130_fd_sc_hd__buf_2
Xinput41 la_data_in[46] vssd1 vssd1 vccd1 vccd1 _2447_/A sky130_fd_sc_hd__clkbuf_2
Xinput63 la_data_in[8] vssd1 vssd1 vccd1 vccd1 _2097_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3134__228 vssd1 vssd1 vccd1 vccd1 _3134__228/HI la_data_out[53] sky130_fd_sc_hd__conb_1
X_2416_ _2416_/A vssd1 vssd1 vccd1 vccd1 _2758_/A sky130_fd_sc_hd__clkbuf_2
X_2347_ _2347_/A vssd1 vssd1 vccd1 vccd1 _2685_/A sky130_fd_sc_hd__clkbuf_2
X_2278_ _2406_/A _2406_/B vssd1 vssd1 vccd1 vccd1 _2827_/A sky130_fd_sc_hd__nand2_2
X_3028__122 vssd1 vssd1 vccd1 vccd1 _3028__122/HI io_oeb[25] sky130_fd_sc_hd__conb_1
XFILLER_40_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2023__A _2023_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2562__A2 _2141_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input19_A la_data_in[26] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1580_ _2972_/A _2926_/A vssd1 vssd1 vccd1 vccd1 _1581_/B sky130_fd_sc_hd__nor2_1
XFILLER_7_187 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2553__A2 _2931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_404 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_415 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_426 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_437 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_448 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2201_ _2201_/A _2201_/B _2201_/C vssd1 vssd1 vccd1 vccd1 _2220_/A sky130_fd_sc_hd__or3_1
XTAP_459 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2132_ _2322_/A vssd1 vssd1 vccd1 vccd1 _2321_/A sky130_fd_sc_hd__buf_2
XFILLER_54_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2063_ _2064_/A _2064_/B vssd1 vssd1 vccd1 vccd1 _2063_/Y sky130_fd_sc_hd__nand2_1
XFILLER_34_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2965_ _2965_/A _2965_/B vssd1 vssd1 vccd1 vccd1 _2965_/Y sky130_fd_sc_hd__nor2_1
X_1916_ _2337_/A vssd1 vssd1 vccd1 vccd1 _1916_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_30_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2896_ _2896_/A vssd1 vssd1 vccd1 vccd1 _2896_/Y sky130_fd_sc_hd__inv_2
XFILLER_8_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1847_ _1847_/A vssd1 vssd1 vccd1 vccd1 _1847_/X sky130_fd_sc_hd__clkbuf_1
X_1778_ _1801_/A vssd1 vssd1 vccd1 vccd1 _1879_/B sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_57_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_53_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2480__A1 _2083_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2480__B2 _2567_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3156__250 vssd1 vssd1 vccd1 vccd1 _3156__250/HI la_data_out[107] sky130_fd_sc_hd__conb_1
XFILLER_4_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2750_ _2933_/A _2748_/X _2749_/X _2936_/A vssd1 vssd1 vccd1 vccd1 _2752_/A sky130_fd_sc_hd__a22o_1
X_1701_ _1731_/B _1701_/B vssd1 vssd1 vccd1 vccd1 _1703_/B sky130_fd_sc_hd__xnor2_1
X_2681_ _2829_/A _2820_/A _2258_/Y _2557_/X _2680_/X vssd1 vssd1 vccd1 vccd1 _2682_/B
+ sky130_fd_sc_hd__a221o_1
X_1632_ _1761_/A _2935_/X _2930_/X _1550_/X vssd1 vssd1 vccd1 vccd1 _1632_/X sky130_fd_sc_hd__a22o_1
X_1563_ _1562_/B _1563_/B vssd1 vssd1 vccd1 vccd1 _1564_/B sky130_fd_sc_hd__and2b_1
XTAP_223 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_212 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_201 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1494_ _2998_/A _2951_/B _2998_/B vssd1 vssd1 vccd1 vccd1 _1494_/X sky130_fd_sc_hd__a21o_1
XTAP_256 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_245 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_234 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_267 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_278 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_289 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2115_ _2127_/A _2235_/B _2235_/A vssd1 vssd1 vccd1 vccd1 _2116_/B sky130_fd_sc_hd__a21oi_1
X_2046_ _2556_/A _2046_/B vssd1 vssd1 vccd1 vccd1 _2070_/B sky130_fd_sc_hd__xnor2_1
XFILLER_35_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2948_ _2949_/A _2950_/B vssd1 vssd1 vccd1 vccd1 _3000_/B sky130_fd_sc_hd__and2b_1
X_2879_ _2758_/X _2773_/X _2772_/A _2686_/X vssd1 vssd1 vccd1 vccd1 _2882_/A sky130_fd_sc_hd__a22o_1
XFILLER_1_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_790 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2211__A input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2802_ _2669_/X _2670_/Y _2789_/A _2789_/B _2793_/B vssd1 vssd1 vccd1 vccd1 _2804_/A
+ sky130_fd_sc_hd__a221o_1
X_2733_ _2733_/A _2733_/B vssd1 vssd1 vccd1 vccd1 _2733_/Y sky130_fd_sc_hd__nand2_1
XFILLER_8_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2664_ _2793_/A _2664_/B vssd1 vssd1 vccd1 vccd1 _2665_/B sky130_fd_sc_hd__nor2_1
XANTENNA__1944__B _1944_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1615_ _1533_/A _1533_/B _1616_/B _1616_/A vssd1 vssd1 vccd1 vccd1 _1615_/X sky130_fd_sc_hd__a22o_1
X_2595_ _2595_/A _2663_/A _2595_/C vssd1 vssd1 vccd1 vccd1 _2603_/A sky130_fd_sc_hd__nor3_2
X_1546_ _2927_/A _2149_/B vssd1 vssd1 vccd1 vccd1 _1547_/S sky130_fd_sc_hd__and2_1
XFILLER_59_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_39_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2029_ _1919_/C _2316_/A _2142_/A _2337_/A vssd1 vssd1 vccd1 vccd1 _2029_/X sky130_fd_sc_hd__a22o_1
XANTENNA__2435__A1 _2434_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_58_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_60_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1764__B _1764_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2380_ _2380_/A _2380_/B vssd1 vssd1 vccd1 vccd1 _2458_/C sky130_fd_sc_hd__or2_1
Xinput6 la_data_in[14] vssd1 vssd1 vccd1 vccd1 input6/X sky130_fd_sc_hd__buf_2
X_3001_ _3001_/A _3001_/B vssd1 vssd1 vccd1 vccd1 _3001_/X sky130_fd_sc_hd__or2_1
XFILLER_49_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3061__155 vssd1 vssd1 vccd1 vccd1 _3061__155/HI io_out[21] sky130_fd_sc_hd__conb_1
XFILLER_20_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3102__196 vssd1 vssd1 vccd1 vccd1 _3102__196/HI la_data_out[21] sky130_fd_sc_hd__conb_1
X_2716_ _2716_/A _2716_/B vssd1 vssd1 vccd1 vccd1 _2731_/B sky130_fd_sc_hd__xor2_2
X_2647_ _2647_/A _2647_/B vssd1 vssd1 vccd1 vccd1 _2880_/A sky130_fd_sc_hd__and2_1
X_2578_ _2578_/A vssd1 vssd1 vccd1 vccd1 _2772_/A sky130_fd_sc_hd__clkbuf_2
X_1529_ _2996_/A _1530_/B vssd1 vssd1 vccd1 vccd1 _1576_/A sky130_fd_sc_hd__nor2_1
XFILLER_19_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input49_A la_data_in[53] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3045__139 vssd1 vssd1 vccd1 vccd1 _3045__139/HI io_out[5] sky130_fd_sc_hd__conb_1
XFILLER_61_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_362 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1880_ _1975_/B vssd1 vssd1 vccd1 vccd1 _2337_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_41_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1775__A _2393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2501_ _2501_/A _2964_/A vssd1 vssd1 vccd1 vccd1 _2501_/Y sky130_fd_sc_hd__nor2_1
X_2432_ _2978_/A input6/X vssd1 vssd1 vccd1 vccd1 _2433_/A sky130_fd_sc_hd__xor2_1
XFILLER_44_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2363_ _2363_/A _2440_/B vssd1 vssd1 vccd1 vccd1 _2450_/B sky130_fd_sc_hd__xor2_2
X_2294_ _2294_/A _2294_/B vssd1 vssd1 vccd1 vccd1 _2294_/Y sky130_fd_sc_hd__nor2_1
XFILLER_2_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2638__A1 _2544_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_20_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_3_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_608 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_619 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2981_ _2936_/X _2930_/A _2980_/X vssd1 vssd1 vccd1 vccd1 _2981_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_14_170 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1932_ _2086_/A _1932_/B vssd1 vssd1 vccd1 vccd1 _1933_/B sky130_fd_sc_hd__xnor2_1
XFILLER_21_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1863_ _1864_/B _1864_/C _2329_/A vssd1 vssd1 vccd1 vccd1 _1865_/B sky130_fd_sc_hd__o21ai_1
Xinput31 la_data_in[37] vssd1 vssd1 vccd1 vccd1 _1910_/A sky130_fd_sc_hd__clkbuf_1
Xinput20 la_data_in[27] vssd1 vssd1 vccd1 vccd1 _2322_/B sky130_fd_sc_hd__clkbuf_2
X_1794_ _1923_/A vssd1 vssd1 vccd1 vccd1 _1924_/A sky130_fd_sc_hd__clkbuf_4
Xinput53 la_data_in[57] vssd1 vssd1 vccd1 vccd1 _1616_/A sky130_fd_sc_hd__buf_2
Xinput42 la_data_in[47] vssd1 vssd1 vccd1 vccd1 _2518_/A sky130_fd_sc_hd__clkbuf_2
Xinput64 la_data_in[9] vssd1 vssd1 vccd1 vccd1 _2097_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_6_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3173__267 vssd1 vssd1 vccd1 vccd1 _3173__267/HI la_data_out[124] sky130_fd_sc_hd__conb_1
X_2415_ _2478_/A vssd1 vssd1 vccd1 vccd1 _2818_/A sky130_fd_sc_hd__buf_6
XFILLER_57_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2346_ _2346_/A _2346_/B vssd1 vssd1 vccd1 vccd1 _2353_/A sky130_fd_sc_hd__nor2_1
XFILLER_57_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2277_ _2406_/A _2348_/B vssd1 vssd1 vccd1 vccd1 _2403_/A sky130_fd_sc_hd__nor2_1
X_3067__161 vssd1 vssd1 vccd1 vccd1 _3067__161/HI io_out[27] sky130_fd_sc_hd__conb_1
XFILLER_16_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_12_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2023__B _2023_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2958__B _2958_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_57_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_57_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2553__A3 _2931_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_405 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_416 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_427 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_438 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2200_ _2199_/B _2199_/C _2199_/A vssd1 vssd1 vccd1 vccd1 _2201_/C sky130_fd_sc_hd__a21oi_1
XTAP_449 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2884__A _2884_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2131_ _2131_/A vssd1 vssd1 vccd1 vccd1 _2552_/A sky130_fd_sc_hd__clkbuf_2
X_2062_ _2062_/A _2062_/B vssd1 vssd1 vccd1 vccd1 _2062_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_34_221 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2964_ _2964_/A vssd1 vssd1 vccd1 vccd1 _2965_/B sky130_fd_sc_hd__clkbuf_2
X_1915_ _1915_/A _1915_/B vssd1 vssd1 vccd1 vccd1 _1915_/Y sky130_fd_sc_hd__xnor2_1
X_2895_ _2795_/B _2795_/C _2894_/Y vssd1 vssd1 vccd1 vccd1 _2898_/A sky130_fd_sc_hd__a21o_1
XFILLER_8_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1846_ _1844_/X _1846_/B vssd1 vssd1 vccd1 vccd1 _1847_/A sky130_fd_sc_hd__and2b_1
X_1777_ _1821_/A _1890_/A vssd1 vssd1 vccd1 vccd1 _1805_/B sky130_fd_sc_hd__nand2_1
XFILLER_1_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2778__B _2807_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1504__A1 _2258_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2329_ _2329_/A _2329_/B _2329_/C vssd1 vssd1 vccd1 vccd1 _2330_/C sky130_fd_sc_hd__or3_1
XFILLER_27_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_43_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input31_A la_data_in[37] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1700_ _2988_/X _1700_/B vssd1 vssd1 vccd1 vccd1 _1701_/B sky130_fd_sc_hd__nor2_1
X_2680_ _2608_/A _2748_/A _2749_/A _2863_/A vssd1 vssd1 vccd1 vccd1 _2680_/X sky130_fd_sc_hd__a22o_1
X_1631_ _2927_/A vssd1 vssd1 vccd1 vccd1 _1761_/A sky130_fd_sc_hd__clkbuf_2
X_1562_ _1563_/B _1562_/B vssd1 vssd1 vccd1 vccd1 _1610_/A sky130_fd_sc_hd__and2b_1
X_1493_ _2960_/A _2960_/B _1490_/A _1492_/X vssd1 vssd1 vccd1 vccd1 _1573_/B sky130_fd_sc_hd__a31o_1
XTAP_224 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_213 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_202 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_257 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_246 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_235 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_268 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_279 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2114_ _2114_/A vssd1 vssd1 vccd1 vccd1 _2235_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_54_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2045_ _2430_/A _2206_/A vssd1 vssd1 vccd1 vccd1 _2046_/B sky130_fd_sc_hd__nand2_1
XFILLER_50_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2947_ _2947_/A _2961_/A vssd1 vssd1 vccd1 vccd1 _2950_/B sky130_fd_sc_hd__xor2_1
X_3179__273 vssd1 vssd1 vccd1 vccd1 _3179__273/HI wbs_dat_o[1] sky130_fd_sc_hd__conb_1
X_2878_ _2909_/A _2909_/B vssd1 vssd1 vccd1 vccd1 _2886_/A sky130_fd_sc_hd__xnor2_1
X_1829_ _1829_/A vssd1 vssd1 vccd1 vccd1 _2028_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_38_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_791 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_780 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2801_ _2801_/A _2801_/B vssd1 vssd1 vccd1 vccd1 _2801_/Y sky130_fd_sc_hd__xnor2_2
X_2732_ _2732_/A _2706_/B vssd1 vssd1 vccd1 vccd1 _2732_/X sky130_fd_sc_hd__or2b_1
XFILLER_8_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2663_ _2663_/A _2719_/A _2663_/C vssd1 vssd1 vccd1 vccd1 _2664_/B sky130_fd_sc_hd__and3_1
X_1614_ _1614_/A _1614_/B vssd1 vssd1 vccd1 vccd1 _1614_/Y sky130_fd_sc_hd__nor2_1
X_2594_ _2523_/X _2518_/B _2593_/X vssd1 vssd1 vccd1 vccd1 _2597_/B sky130_fd_sc_hd__a21o_1
X_1545_ _1605_/A _1545_/B vssd1 vssd1 vccd1 vccd1 _1557_/A sky130_fd_sc_hd__nand2_4
XFILLER_59_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3107__201 vssd1 vssd1 vccd1 vccd1 _3107__201/HI la_data_out[26] sky130_fd_sc_hd__conb_1
X_2028_ _2028_/A vssd1 vssd1 vccd1 vccd1 _2316_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_42_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput7 la_data_in[15] vssd1 vssd1 vccd1 vccd1 input7/X sky130_fd_sc_hd__clkbuf_2
XFILLER_37_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3000_ _3000_/A _3000_/B vssd1 vssd1 vccd1 vccd1 _3001_/B sky130_fd_sc_hd__or2_1
XFILLER_49_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2715_ _2715_/A _2715_/B vssd1 vssd1 vccd1 vccd1 _2716_/B sky130_fd_sc_hd__xnor2_2
XANTENNA__2132__A _2322_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2646_ _2404_/X _2578_/A _2774_/A _2273_/X vssd1 vssd1 vccd1 vccd1 _2649_/A sky130_fd_sc_hd__a22o_1
XFILLER_10_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2577_ _2577_/A _2577_/B vssd1 vssd1 vccd1 vccd1 _2583_/A sky130_fd_sc_hd__nand2_1
X_1528_ _1566_/A _1528_/B vssd1 vssd1 vccd1 vccd1 _1530_/B sky130_fd_sc_hd__and2_1
XFILLER_19_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_168 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3084__178 vssd1 vssd1 vccd1 vccd1 _3084__178/HI la_data_out[3] sky130_fd_sc_hd__conb_1
XPHY_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_540 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2500_ _2647_/A _2647_/B vssd1 vssd1 vccd1 vccd1 _2964_/A sky130_fd_sc_hd__nand2_2
XFILLER_6_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2431_ _2353_/A _2353_/B _2346_/A vssd1 vssd1 vccd1 vccd1 _2434_/B sky130_fd_sc_hd__a21o_1
X_2362_ _2288_/A _2288_/B _2361_/Y vssd1 vssd1 vccd1 vccd1 _2440_/B sky130_fd_sc_hd__o21ai_2
XFILLER_37_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2293_ _2374_/A _2305_/B vssd1 vssd1 vccd1 vccd1 _2294_/B sky130_fd_sc_hd__and2b_1
XFILLER_64_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_52_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1966__A _2138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_32_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2797__A _2797_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2629_ _2629_/A _2629_/B vssd1 vssd1 vccd1 vccd1 _2630_/D sky130_fd_sc_hd__xnor2_4
XFILLER_47_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input61_A la_data_in[6] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_609 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3012__106 vssd1 vssd1 vccd1 vccd1 _3012__106/HI io_oeb[9] sky130_fd_sc_hd__conb_1
XFILLER_3_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2980_ _2740_/X _2934_/X _2935_/A _2933_/A vssd1 vssd1 vccd1 vccd1 _2980_/X sky130_fd_sc_hd__a22o_1
X_1931_ _1817_/A _2022_/A _1929_/Y _2027_/A _1930_/X vssd1 vssd1 vccd1 vccd1 _1932_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_14_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1862_ _1817_/A _2028_/A _2022_/A _1800_/A vssd1 vssd1 vccd1 vccd1 _1864_/C sky130_fd_sc_hd__a22o_1
Xinput21 la_data_in[28] vssd1 vssd1 vccd1 vccd1 _2380_/B sky130_fd_sc_hd__buf_2
Xinput10 la_data_in[18] vssd1 vssd1 vccd1 vccd1 _1923_/A sky130_fd_sc_hd__clkbuf_2
Xinput32 la_data_in[38] vssd1 vssd1 vccd1 vccd1 _1959_/A sky130_fd_sc_hd__clkbuf_1
Xinput54 la_data_in[58] vssd1 vssd1 vccd1 vccd1 _1613_/A sky130_fd_sc_hd__clkbuf_2
Xinput43 la_data_in[48] vssd1 vssd1 vccd1 vccd1 _2597_/A sky130_fd_sc_hd__buf_2
X_1793_ _2013_/A vssd1 vssd1 vccd1 vccd1 _1968_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__2410__A _2410_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2414_ _2556_/A _2414_/B vssd1 vssd1 vccd1 vccd1 _2492_/A sky130_fd_sc_hd__xnor2_1
XFILLER_57_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2345_ _2345_/A _2345_/B vssd1 vssd1 vccd1 vccd1 _2346_/B sky130_fd_sc_hd__nor2_1
XFILLER_29_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2276_ input3/X input4/X vssd1 vssd1 vccd1 vccd1 _2348_/B sky130_fd_sc_hd__xnor2_1
XFILLER_37_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_156 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_406 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_417 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_428 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_439 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2130_ _2130_/A vssd1 vssd1 vccd1 vccd1 _2130_/X sky130_fd_sc_hd__clkbuf_2
X_2061_ _2002_/X _2005_/B _2003_/A vssd1 vssd1 vccd1 vccd1 _2062_/B sky130_fd_sc_hd__a21o_1
XFILLER_47_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2963_ _2963_/A _2963_/B vssd1 vssd1 vccd1 vccd1 _2970_/B sky130_fd_sc_hd__and2_2
XFILLER_34_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3140__234 vssd1 vssd1 vccd1 vccd1 _3140__234/HI la_data_out[59] sky130_fd_sc_hd__conb_1
X_1914_ _1873_/A _1873_/B _1913_/X vssd1 vssd1 vccd1 vccd1 _1915_/B sky130_fd_sc_hd__a21o_1
X_2894_ _2850_/A _2896_/A _2790_/A vssd1 vssd1 vccd1 vccd1 _2894_/Y sky130_fd_sc_hd__o21ai_1
X_1845_ _1845_/A _1845_/B _1843_/Y vssd1 vssd1 vccd1 vccd1 _1846_/B sky130_fd_sc_hd__or3b_1
X_1776_ input9/X vssd1 vssd1 vccd1 vccd1 _1890_/A sky130_fd_sc_hd__clkbuf_2
X_2328_ _2329_/B _2329_/C _2700_/A vssd1 vssd1 vccd1 vccd1 _2330_/B sky130_fd_sc_hd__o21ai_2
XFILLER_27_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2259_ _2134_/C _2316_/A _2386_/A _2131_/A vssd1 vssd1 vccd1 vccd1 _2259_/X sky130_fd_sc_hd__a22o_1
XFILLER_25_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_4_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input24_A la_data_in[30] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_369 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_550 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3124__218 vssd1 vssd1 vccd1 vccd1 _3124__218/HI la_data_out[43] sky130_fd_sc_hd__conb_1
XFILLER_16_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1630_ _1681_/A _1630_/B vssd1 vssd1 vccd1 vccd1 _1638_/A sky130_fd_sc_hd__and2_1
XFILLER_8_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3018__112 vssd1 vssd1 vccd1 vccd1 _3018__112/HI io_oeb[15] sky130_fd_sc_hd__conb_1
X_1561_ _1561_/A _1561_/B vssd1 vssd1 vccd1 vccd1 _1562_/B sky130_fd_sc_hd__xor2_1
X_1492_ _1488_/A _1488_/B _1491_/X vssd1 vssd1 vccd1 vccd1 _1492_/X sky130_fd_sc_hd__o21a_1
XTAP_214 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_203 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_247 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_236 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_225 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_258 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_269 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2113_ _2127_/A _2114_/A _2235_/B vssd1 vssd1 vccd1 vccd1 _2116_/A sky130_fd_sc_hd__and3_1
X_2044_ _2044_/A vssd1 vssd1 vccd1 vccd1 _2206_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_47_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2946_ _2888_/A _2888_/B _2945_/X vssd1 vssd1 vccd1 vccd1 _2961_/A sky130_fd_sc_hd__a21oi_1
X_2877_ _2877_/A _2920_/B vssd1 vssd1 vccd1 vccd1 _2909_/B sky130_fd_sc_hd__xnor2_1
X_1828_ _1884_/B _1831_/A vssd1 vssd1 vccd1 vccd1 _1829_/A sky130_fd_sc_hd__and2b_1
XANTENNA__1974__A _1974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1759_ _1759_/A _1759_/B vssd1 vssd1 vccd1 vccd1 _1760_/B sky130_fd_sc_hd__xor2_1
XFILLER_2_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_770 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_792 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_781 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_63_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2800_ _2723_/A _2723_/B _2729_/A vssd1 vssd1 vccd1 vccd1 _2801_/B sky130_fd_sc_hd__a21boi_1
X_2731_ _2731_/A _2731_/B vssd1 vssd1 vccd1 vccd1 _2789_/A sky130_fd_sc_hd__nand2_1
X_2662_ _2719_/A _2663_/C _2663_/A vssd1 vssd1 vccd1 vccd1 _2793_/A sky130_fd_sc_hd__a21oi_1
X_1613_ _1613_/A _1613_/B vssd1 vssd1 vccd1 vccd1 _1657_/A sky130_fd_sc_hd__xnor2_1
X_2593_ _2663_/A _2595_/C _2595_/A vssd1 vssd1 vccd1 vccd1 _2593_/X sky130_fd_sc_hd__o21a_1
X_1544_ _1544_/A _1544_/B _1544_/C vssd1 vssd1 vccd1 vccd1 _1545_/B sky130_fd_sc_hd__or3_1
XFILLER_27_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_39_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3146__240 vssd1 vssd1 vccd1 vccd1 _3146__240/HI la_data_out[97] sky130_fd_sc_hd__conb_1
X_2027_ _2027_/A vssd1 vssd1 vccd1 vccd1 _2027_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_42_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2929_ _2962_/A _2962_/B vssd1 vssd1 vccd1 vccd1 _2963_/A sky130_fd_sc_hd__xor2_4
XFILLER_10_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_49_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput8 la_data_in[16] vssd1 vssd1 vccd1 vccd1 input8/X sky130_fd_sc_hd__buf_2
XFILLER_37_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_32_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2714_ _2733_/A _2733_/B vssd1 vssd1 vccd1 vccd1 _2715_/B sky130_fd_sc_hd__xnor2_2
X_2645_ _2645_/A _2645_/B vssd1 vssd1 vccd1 vccd1 _2651_/B sky130_fd_sc_hd__and2_1
X_2576_ _2573_/Y _2574_/X _2528_/Y _2529_/X vssd1 vssd1 vccd1 vccd1 _2585_/B sky130_fd_sc_hd__a211o_1
X_1527_ _1527_/A _1527_/B _1527_/C vssd1 vssd1 vccd1 vccd1 _1528_/B sky130_fd_sc_hd__or3_1
XFILLER_19_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2813__B1 _2739_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_103 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1607__A1 _1561_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_10_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2430_ _2430_/A vssd1 vssd1 vccd1 vccd1 _2434_/A sky130_fd_sc_hd__buf_2
XFILLER_6_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2361_ _2361_/A _2361_/B vssd1 vssd1 vccd1 vccd1 _2361_/Y sky130_fd_sc_hd__nand2_1
X_2292_ _2374_/A _2374_/B vssd1 vssd1 vccd1 vccd1 _2294_/A sky130_fd_sc_hd__and2_1
XFILLER_2_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_434 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1982__A _2009_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2628_ _2467_/A _2467_/B _2467_/C _2536_/C vssd1 vssd1 vccd1 vccd1 _2630_/C sky130_fd_sc_hd__a211oi_1
X_2559_ _2559_/A vssd1 vssd1 vccd1 vccd1 _2829_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_46_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_23_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input54_A la_data_in[58] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3051__145 vssd1 vssd1 vccd1 vccd1 _3051__145/HI io_out[11] sky130_fd_sc_hd__conb_1
XFILLER_59_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_19_478 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1930_ _2020_/A _1829_/A _1832_/A _1926_/A vssd1 vssd1 vccd1 vccd1 _1930_/X sky130_fd_sc_hd__a22o_1
X_1861_ _1884_/A _1884_/B _1861_/C vssd1 vssd1 vccd1 vccd1 _2022_/A sky130_fd_sc_hd__and3b_1
XFILLER_14_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput22 la_data_in[29] vssd1 vssd1 vccd1 vccd1 _2464_/B sky130_fd_sc_hd__buf_2
Xinput11 la_data_in[19] vssd1 vssd1 vccd1 vccd1 _1972_/A sky130_fd_sc_hd__clkbuf_2
Xinput33 la_data_in[39] vssd1 vssd1 vccd1 vccd1 _2002_/A sky130_fd_sc_hd__clkbuf_1
Xinput44 la_data_in[49] vssd1 vssd1 vccd1 vccd1 _2725_/A sky130_fd_sc_hd__clkbuf_4
Xinput55 la_data_in[59] vssd1 vssd1 vccd1 vccd1 _1655_/A sky130_fd_sc_hd__clkbuf_2
X_1792_ _1890_/A vssd1 vssd1 vccd1 vccd1 _1939_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_6_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2413_ _2026_/Y _2557_/A _2558_/A _2568_/A _2412_/X vssd1 vssd1 vccd1 vccd1 _2414_/B
+ sky130_fd_sc_hd__a221o_1
X_2344_ _2345_/A _2345_/B vssd1 vssd1 vccd1 vccd1 _2346_/A sky130_fd_sc_hd__and2_1
XFILLER_57_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2275_ _2406_/B _2406_/A vssd1 vssd1 vccd1 vccd1 _2347_/A sky130_fd_sc_hd__and2b_1
XANTENNA__2138__A _2138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3035__129 vssd1 vssd1 vccd1 vccd1 _3035__129/HI io_oeb[32] sky130_fd_sc_hd__conb_1
XFILLER_0_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_0_536 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_407 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_418 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_429 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2060_ _2060_/A _2059_/X vssd1 vssd1 vccd1 vccd1 _2062_/A sky130_fd_sc_hd__or2b_1
XFILLER_47_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_267 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2962_ _2962_/A _2962_/B vssd1 vssd1 vccd1 vccd1 _2970_/A sky130_fd_sc_hd__and2_2
X_1913_ _1875_/A _1913_/B vssd1 vssd1 vccd1 vccd1 _1913_/X sky130_fd_sc_hd__and2b_1
X_2893_ _3000_/A _2892_/Y vssd1 vssd1 vccd1 vccd1 _2899_/A sky130_fd_sc_hd__or2b_2
X_1844_ _1845_/A _1845_/B _1843_/Y vssd1 vssd1 vccd1 vccd1 _1844_/X sky130_fd_sc_hd__o21ba_1
X_1775_ _2393_/A _2430_/A _1775_/C vssd1 vssd1 vccd1 vccd1 _1788_/A sky130_fd_sc_hd__and3_1
XFILLER_8_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2327_ _2329_/A vssd1 vssd1 vccd1 vccd1 _2700_/A sky130_fd_sc_hd__clkbuf_4
X_2258_ _2258_/A _2258_/B vssd1 vssd1 vccd1 vccd1 _2258_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_27_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_551 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2189_ _2189_/A _2255_/A vssd1 vssd1 vccd1 vccd1 _2189_/X sky130_fd_sc_hd__or2_1
XFILLER_53_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_21_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2985__B _2985_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input17_A la_data_in[24] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2456__A1 _2393_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3163__257 vssd1 vssd1 vccd1 vccd1 _3163__257/HI la_data_out[114] sky130_fd_sc_hd__conb_1
XFILLER_16_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2208__B2 _1939_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2208__A1 _1888_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3204__298 vssd1 vssd1 vccd1 vccd1 _3204__298/HI wbs_dat_o[26] sky130_fd_sc_hd__conb_1
XFILLER_8_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3057__151 vssd1 vssd1 vccd1 vccd1 _3057__151/HI io_out[17] sky130_fd_sc_hd__conb_1
X_1560_ _1560_/A _1560_/B vssd1 vssd1 vccd1 vccd1 _1561_/B sky130_fd_sc_hd__nor2_1
X_1491_ _2954_/A _2954_/B _1488_/B _1488_/A vssd1 vssd1 vccd1 vccd1 _1491_/X sky130_fd_sc_hd__a22o_1
XTAP_215 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_204 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_248 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_237 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_226 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2144__B1 _2141_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_259 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2112_ _2112_/A _2112_/B vssd1 vssd1 vccd1 vccd1 _2235_/B sky130_fd_sc_hd__or2_2
XFILLER_54_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2043_ _2043_/A _2097_/A vssd1 vssd1 vccd1 vccd1 _2044_/A sky130_fd_sc_hd__xor2_1
XANTENNA__2416__A _2416_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2945_ _2887_/B _2945_/B vssd1 vssd1 vccd1 vccd1 _2945_/X sky130_fd_sc_hd__and2b_1
X_2876_ _2912_/A _2912_/B vssd1 vssd1 vccd1 vccd1 _2920_/B sky130_fd_sc_hd__xnor2_2
XFILLER_30_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1827_ _1897_/A _1830_/B vssd1 vssd1 vccd1 vccd1 _1884_/B sky130_fd_sc_hd__xor2_2
X_1758_ _1730_/A _1730_/B _1733_/A vssd1 vssd1 vccd1 vccd1 _1759_/B sky130_fd_sc_hd__o21bai_1
X_1689_ _1689_/A _1741_/A vssd1 vssd1 vccd1 vccd1 _1690_/B sky130_fd_sc_hd__or2_2
XFILLER_1_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_760 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_input9_A la_data_in[17] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_793 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_782 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_771 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_54_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2730_ _2730_/A vssd1 vssd1 vccd1 vccd1 _2730_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_8_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2661_ _2657_/Y _2658_/X _2589_/B _2589_/Y vssd1 vssd1 vccd1 vccd1 _2663_/C sky130_fd_sc_hd__a211o_1
XFILLER_60_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1612_ _1612_/A _1612_/B vssd1 vssd1 vccd1 vccd1 _1613_/B sky130_fd_sc_hd__xnor2_4
XFILLER_8_296 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3005__99 vssd1 vssd1 vccd1 vccd1 _3005__99/HI io_oeb[2] sky130_fd_sc_hd__conb_1
X_2592_ _2589_/Y _2590_/X _2524_/Y _2525_/Y vssd1 vssd1 vccd1 vccd1 _2595_/C sky130_fd_sc_hd__o211a_1
X_1543_ _1544_/A _1544_/B _1544_/C vssd1 vssd1 vccd1 vccd1 _1605_/A sky130_fd_sc_hd__o21ai_4
XFILLER_5_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_54_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2026_ _2026_/A _2026_/B vssd1 vssd1 vccd1 vccd1 _2026_/Y sky130_fd_sc_hd__xnor2_4
XANTENNA__2146__A _2179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2928_ _1944_/B _2972_/A _2928_/S vssd1 vssd1 vccd1 vccd1 _2962_/B sky130_fd_sc_hd__mux2_2
X_2859_ _2845_/A _2845_/B _2858_/X vssd1 vssd1 vccd1 vccd1 _2945_/B sky130_fd_sc_hd__a21o_1
XFILLER_40_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_590 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_129 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_53_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3169__263 vssd1 vssd1 vccd1 vccd1 _3169__263/HI la_data_out[120] sky130_fd_sc_hd__conb_1
XFILLER_39_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput9 la_data_in[17] vssd1 vssd1 vccd1 vccd1 input9/X sky130_fd_sc_hd__clkbuf_4
XFILLER_36_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_498 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2713_ _2783_/A _2713_/B vssd1 vssd1 vccd1 vccd1 _2733_/B sky130_fd_sc_hd__and2_1
X_2644_ _2644_/A _2644_/B vssd1 vssd1 vccd1 vccd1 _2651_/A sky130_fd_sc_hd__and2_1
X_2575_ _2528_/Y _2529_/X _2573_/Y _2574_/X vssd1 vssd1 vccd1 vccd1 _2585_/A sky130_fd_sc_hd__o211ai_2
X_1526_ _1527_/A _1527_/B _1527_/C vssd1 vssd1 vccd1 vccd1 _1566_/A sky130_fd_sc_hd__o21ai_2
XFILLER_35_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2009_ _2009_/A _1982_/B vssd1 vssd1 vccd1 vccd1 _2108_/A sky130_fd_sc_hd__or2b_1
XFILLER_23_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1855__A2 _1979_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_61_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_354 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2360_ _2438_/B _2360_/B vssd1 vssd1 vccd1 vccd1 _2363_/A sky130_fd_sc_hd__or2_1
X_2291_ _2305_/A _2305_/B vssd1 vssd1 vccd1 vccd1 _2374_/B sky130_fd_sc_hd__xnor2_1
XFILLER_1_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_37_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2627_ _2694_/B vssd1 vssd1 vccd1 vccd1 _2630_/B sky130_fd_sc_hd__inv_2
XANTENNA__2326__A3 _2931_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2558_ _2558_/A vssd1 vssd1 vccd1 vccd1 _2820_/A sky130_fd_sc_hd__clkbuf_2
X_1509_ _2810_/A _2749_/X _2820_/X _2922_/X vssd1 vssd1 vccd1 vccd1 _1509_/X sky130_fd_sc_hd__a22o_1
X_2489_ _2583_/B _2489_/B vssd1 vssd1 vccd1 vccd1 _2529_/B sky130_fd_sc_hd__and2_1
XFILLER_46_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2798__B1 _2797_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_11_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_339 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input47_A la_data_in[51] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3090__184 vssd1 vssd1 vccd1 vccd1 _3090__184/HI la_data_out[9] sky130_fd_sc_hd__conb_1
XFILLER_19_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_59_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1860_ _2377_/A _1859_/Y _1832_/A _1890_/A vssd1 vssd1 vccd1 vccd1 _1864_/B sky130_fd_sc_hd__a2bb2o_1
XFILLER_42_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
Xinput12 la_data_in[1] vssd1 vssd1 vccd1 vccd1 _1801_/A sky130_fd_sc_hd__clkbuf_1
X_1791_ _1791_/A vssd1 vssd1 vccd1 vccd1 _1816_/A sky130_fd_sc_hd__clkbuf_2
Xinput45 la_data_in[4] vssd1 vssd1 vccd1 vccd1 _1897_/A sky130_fd_sc_hd__clkbuf_2
Xinput23 la_data_in[2] vssd1 vssd1 vccd1 vccd1 _1830_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput34 la_data_in[3] vssd1 vssd1 vccd1 vccd1 _1830_/B sky130_fd_sc_hd__dlymetal6s2s_1
Xinput56 la_data_in[5] vssd1 vssd1 vccd1 vccd1 _1944_/A sky130_fd_sc_hd__clkbuf_1
X_2412_ _2686_/A _2748_/A _2560_/A _2567_/A vssd1 vssd1 vccd1 vccd1 _2412_/X sky130_fd_sc_hd__a22o_1
XFILLER_42_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2343_ _2478_/A _2343_/B vssd1 vssd1 vccd1 vccd1 _2345_/B sky130_fd_sc_hd__xnor2_1
X_2274_ input5/X input4/X vssd1 vssd1 vccd1 vccd1 _2406_/B sky130_fd_sc_hd__xor2_2
XANTENNA__2419__A _2739_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2138__B _2188_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_427 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_20_132 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1989_ _1859_/Y _2417_/A _1947_/A _1939_/A vssd1 vssd1 vccd1 vccd1 _1989_/X sky130_fd_sc_hd__a2bb2o_1
X_3074__168 vssd1 vssd1 vccd1 vccd1 _3074__168/HI io_out[34] sky130_fd_sc_hd__conb_1
XFILLER_57_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_28_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_342 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_408 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_419 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3209__303 vssd1 vssd1 vccd1 vccd1 _3209__303/HI wbs_dat_o[31] sky130_fd_sc_hd__conb_1
XFILLER_47_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2961_ _2961_/A _2947_/A vssd1 vssd1 vccd1 vccd1 _2998_/A sky130_fd_sc_hd__or2b_1
XFILLER_15_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1912_ _1912_/A _1911_/X vssd1 vssd1 vccd1 vccd1 _1915_/A sky130_fd_sc_hd__or2b_1
XFILLER_30_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2892_ _2892_/A _2892_/B vssd1 vssd1 vccd1 vccd1 _2892_/Y sky130_fd_sc_hd__nand2_1
XFILLER_8_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1843_ _1843_/A _1843_/B vssd1 vssd1 vccd1 vccd1 _1843_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_30_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1774_ _1899_/A vssd1 vssd1 vccd1 vccd1 _2430_/A sky130_fd_sc_hd__clkbuf_2
X_2326_ _2027_/X _2378_/A _2931_/B _2194_/A _2552_/A vssd1 vssd1 vccd1 vccd1 _2329_/C
+ sky130_fd_sc_hd__a32o_1
X_2257_ _2139_/B _2189_/X _2256_/X _2190_/A vssd1 vssd1 vccd1 vccd1 _2258_/B sky130_fd_sc_hd__a31o_1
XFILLER_38_530 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_53_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2188_ _2188_/A _2188_/B vssd1 vssd1 vccd1 vccd1 _2190_/A sky130_fd_sc_hd__and2_1
XFILLER_25_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3096__190 vssd1 vssd1 vccd1 vccd1 _3096__190/HI la_data_out[15] sky130_fd_sc_hd__conb_1
X_1490_ _1490_/A _1490_/B vssd1 vssd1 vccd1 vccd1 _1490_/X sky130_fd_sc_hd__xor2_1
XTAP_205 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_238 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_227 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_216 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2144__A1 _2410_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_249 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_90 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2111_ _2111_/A _2111_/B vssd1 vssd1 vccd1 vccd1 _2114_/A sky130_fd_sc_hd__xnor2_1
X_2042_ _2209_/A vssd1 vssd1 vccd1 vccd1 _2556_/A sky130_fd_sc_hd__buf_2
XFILLER_47_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_62_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2944_ _2944_/A _2944_/B vssd1 vssd1 vccd1 vccd1 _2947_/A sky130_fd_sc_hd__xor2_1
X_2875_ _2911_/A _2911_/B vssd1 vssd1 vccd1 vccd1 _2912_/B sky130_fd_sc_hd__xor2_2
XFILLER_30_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1826_ _1981_/A vssd1 vssd1 vccd1 vccd1 _2086_/A sky130_fd_sc_hd__clkinv_4
XANTENNA__2432__A _2978_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1757_ _1736_/A _1736_/B _1739_/A _1756_/X vssd1 vssd1 vccd1 vccd1 _1760_/A sky130_fd_sc_hd__a211o_1
X_1688_ _1688_/A _1688_/B vssd1 vssd1 vccd1 vccd1 _1741_/A sky130_fd_sc_hd__nor2_1
XTAP_761 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_750 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_794 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_783 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_772 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2309_ _2309_/A _2285_/B vssd1 vssd1 vccd1 vccd1 _2309_/X sky130_fd_sc_hd__or2b_1
XFILLER_38_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1511__A _2926_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_54_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_26_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2607__A _2739_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3130__224 vssd1 vssd1 vccd1 vccd1 _3130__224/HI la_data_out[49] sky130_fd_sc_hd__conb_1
XFILLER_0_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2660_ _2718_/A vssd1 vssd1 vccd1 vccd1 _2719_/A sky130_fd_sc_hd__clkbuf_2
X_1611_ _1611_/A _1659_/A vssd1 vssd1 vccd1 vccd1 _1612_/B sky130_fd_sc_hd__or2_2
X_2591_ _2524_/Y _2525_/Y _2589_/Y _2590_/X vssd1 vssd1 vccd1 vccd1 _2663_/A sky130_fd_sc_hd__a211oi_4
X_1542_ _2936_/X _2772_/X _1540_/Y _1541_/X vssd1 vssd1 vccd1 vccd1 _1544_/C sky130_fd_sc_hd__a211o_1
XFILLER_5_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2025_ _1977_/A _1977_/B _1976_/A vssd1 vssd1 vccd1 vccd1 _2026_/B sky130_fd_sc_hd__a21oi_2
XFILLER_62_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2927_ _2927_/A _2927_/B vssd1 vssd1 vccd1 vccd1 _2928_/S sky130_fd_sc_hd__nand2_1
X_2858_ _2837_/B _2858_/B vssd1 vssd1 vccd1 vccd1 _2858_/X sky130_fd_sc_hd__and2b_1
X_1809_ _1810_/A _1810_/B vssd1 vssd1 vccd1 vccd1 _1845_/A sky130_fd_sc_hd__and2_1
X_2789_ _2789_/A _2789_/B vssd1 vssd1 vccd1 vccd1 _2790_/B sky130_fd_sc_hd__or2_1
X_3114__208 vssd1 vssd1 vccd1 vccd1 _3114__208/HI la_data_out[33] sky130_fd_sc_hd__conb_1
XFILLER_49_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_591 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_580 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_61_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_26_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3008__102 vssd1 vssd1 vccd1 vccd1 _3008__102/HI io_oeb[5] sky130_fd_sc_hd__conb_1
XFILLER_53_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_26_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2072__A _2188_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_403 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_64_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_458 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_17_352 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_32_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2712_ _2712_/A _2712_/B _2712_/C vssd1 vssd1 vccd1 vccd1 _2713_/B sky130_fd_sc_hd__or3_1
XANTENNA__2338__A1 _2567_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2643_ _2642_/B _2642_/C _2642_/A vssd1 vssd1 vccd1 vccd1 _2653_/B sky130_fd_sc_hd__a21oi_1
X_2574_ _2573_/A _2573_/B _2573_/C vssd1 vssd1 vccd1 vccd1 _2574_/X sky130_fd_sc_hd__a21o_1
X_1525_ _2971_/A _1525_/B vssd1 vssd1 vccd1 vccd1 _1527_/C sky130_fd_sc_hd__xnor2_1
XFILLER_28_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2008_ _2008_/A _2008_/B _2053_/B vssd1 vssd1 vccd1 vccd1 _2064_/A sky130_fd_sc_hd__or3_1
XFILLER_23_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_58_274 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_19_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2265__B1 _2083_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3136__230 vssd1 vssd1 vccd1 vccd1 _3136__230/HI la_data_out[55] sky130_fd_sc_hd__conb_1
X_2290_ _2307_/A _2307_/B vssd1 vssd1 vccd1 vccd1 _2305_/B sky130_fd_sc_hd__xor2_1
XFILLER_2_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2626_ _2694_/A vssd1 vssd1 vccd1 vccd1 _2630_/A sky130_fd_sc_hd__inv_2
X_2557_ _2557_/A vssd1 vssd1 vccd1 vccd1 _2557_/X sky130_fd_sc_hd__buf_2
X_1508_ _1561_/A _1508_/B vssd1 vssd1 vccd1 vccd1 _1521_/A sky130_fd_sc_hd__and2b_2
X_2488_ _2488_/A _2488_/B vssd1 vssd1 vccd1 vccd1 _2489_/B sky130_fd_sc_hd__or2_1
XFILLER_55_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_7_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2525__A _2525_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1790_ input1/X vssd1 vssd1 vccd1 vccd1 _1791_/A sky130_fd_sc_hd__inv_2
Xinput13 la_data_in[20] vssd1 vssd1 vccd1 vccd1 _1974_/A sky130_fd_sc_hd__clkbuf_2
Xinput35 la_data_in[40] vssd1 vssd1 vccd1 vccd1 _2059_/A sky130_fd_sc_hd__clkbuf_1
Xinput24 la_data_in[30] vssd1 vssd1 vccd1 vccd1 _2629_/A sky130_fd_sc_hd__buf_4
Xinput46 la_data_in[50] vssd1 vssd1 vccd1 vccd1 _2723_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_6_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput57 la_data_in[60] vssd1 vssd1 vccd1 vccd1 _1723_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_2411_ _2411_/A vssd1 vssd1 vccd1 vccd1 _2748_/A sky130_fd_sc_hd__clkbuf_2
X_2342_ _2410_/A _1988_/A _2141_/Y _2037_/X _2341_/X vssd1 vssd1 vccd1 vccd1 _2343_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_35_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1604__A _1605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2273_ _2273_/A vssd1 vssd1 vccd1 vccd1 _2273_/X sky130_fd_sc_hd__clkbuf_2
XANTENNA__2477__B1 _2258_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2419__B _2965_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_200 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_37_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2154__B _2775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_33_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_20_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1988_ _1988_/A vssd1 vssd1 vccd1 vccd1 _2609_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__2401__B1 _2400_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2609_ _2609_/A vssd1 vssd1 vccd1 vccd1 _2609_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_57_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_16_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_409 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2960_ _2960_/A _2960_/B vssd1 vssd1 vccd1 vccd1 _2960_/X sky130_fd_sc_hd__xor2_2
X_1911_ _1963_/A _1910_/C _1910_/A vssd1 vssd1 vccd1 vccd1 _1911_/X sky130_fd_sc_hd__a21o_1
XFILLER_15_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2891_ _2892_/A _2892_/B vssd1 vssd1 vccd1 vccd1 _3000_/A sky130_fd_sc_hd__nor2_1
X_1842_ _1848_/A _1848_/B vssd1 vssd1 vccd1 vccd1 _1843_/B sky130_fd_sc_hd__xor2_1
XFILLER_30_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1773_ _1800_/A vssd1 vssd1 vccd1 vccd1 _1899_/A sky130_fd_sc_hd__buf_2
X_2325_ _2458_/A _2325_/B _2461_/A vssd1 vssd1 vccd1 vccd1 _2931_/B sky130_fd_sc_hd__or3_4
X_2256_ _2083_/A _2083_/B _2192_/B vssd1 vssd1 vccd1 vccd1 _2256_/X sky130_fd_sc_hd__a21bo_1
X_2187_ _2187_/A _2187_/B _2187_/C _2083_/B vssd1 vssd1 vccd1 vccd1 _2192_/C sky130_fd_sc_hd__or4b_2
XFILLER_38_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3041__135 vssd1 vssd1 vccd1 vccd1 _3041__135/HI io_out[1] sky130_fd_sc_hd__conb_1
XANTENNA__2925__A1 _2819_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_206 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_239 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_228 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_217 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2110_ _2164_/B _2110_/B vssd1 vssd1 vccd1 vccd1 _2111_/B sky130_fd_sc_hd__xnor2_1
XFILLER_54_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2041_ _2269_/A vssd1 vssd1 vccd1 vccd1 _2209_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_35_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3025__119 vssd1 vssd1 vccd1 vccd1 _3025__119/HI io_oeb[22] sky130_fd_sc_hd__conb_1
XFILLER_35_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2943_ _2943_/A _2943_/B vssd1 vssd1 vccd1 vccd1 _2944_/B sky130_fd_sc_hd__xor2_1
XFILLER_30_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2874_ _2972_/A _2874_/B vssd1 vssd1 vccd1 vccd1 _2911_/B sky130_fd_sc_hd__xnor2_2
X_1825_ _1897_/A vssd1 vssd1 vccd1 vccd1 _1981_/A sky130_fd_sc_hd__buf_2
XANTENNA__2432__B input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1756_ _1756_/A _1756_/B vssd1 vssd1 vccd1 vccd1 _1756_/X sky130_fd_sc_hd__and2_1
X_1687_ _1688_/A _1688_/B vssd1 vssd1 vccd1 vccd1 _1689_/A sky130_fd_sc_hd__and2_1
XTAP_751 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_740 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_795 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_784 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_773 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_762 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2308_ _2308_/A _2308_/B vssd1 vssd1 vccd1 vccd1 _2308_/X sky130_fd_sc_hd__or2_1
X_2239_ _2240_/A _2240_/B vssd1 vssd1 vccd1 vccd1 _2241_/A sky130_fd_sc_hd__and2_1
XFILLER_26_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input22_A la_data_in[29] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_48_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1860__A2_N _1859_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_250 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1610_ _1610_/A _1610_/B vssd1 vssd1 vccd1 vccd1 _1659_/A sky130_fd_sc_hd__nor2_1
XFILLER_8_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2590_ _2589_/B _2589_/C _2589_/A vssd1 vssd1 vccd1 vccd1 _2590_/X sky130_fd_sc_hd__o21a_1
X_1541_ _2933_/X _2773_/X _2966_/X _2863_/X vssd1 vssd1 vccd1 vccd1 _1541_/X sky130_fd_sc_hd__a22o_1
XFILLER_4_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2024_ _2024_/A vssd1 vssd1 vccd1 vccd1 _2026_/A sky130_fd_sc_hd__clkinv_2
XFILLER_62_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2926_ _2926_/A _2926_/B vssd1 vssd1 vccd1 vccd1 _2962_/A sky130_fd_sc_hd__xnor2_2
XFILLER_50_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2857_ _2848_/B _2857_/B vssd1 vssd1 vccd1 vccd1 _2892_/A sky130_fd_sc_hd__and2b_1
X_1808_ _1839_/A _1839_/B _1806_/Y _1848_/A vssd1 vssd1 vccd1 vccd1 _1810_/B sky130_fd_sc_hd__o211a_1
X_2788_ _2789_/A _2789_/B vssd1 vssd1 vccd1 vccd1 _2790_/A sky130_fd_sc_hd__nand2_1
X_1739_ _1739_/A _1739_/B vssd1 vssd1 vccd1 vccd1 _1740_/B sky130_fd_sc_hd__or2_2
X_3153__247 vssd1 vssd1 vccd1 vccd1 _3153__247/HI la_data_out[104] sky130_fd_sc_hd__conb_1
XTAP_570 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_581 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_592 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_18_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2618__A _2824_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3047__141 vssd1 vssd1 vccd1 vccd1 _3047__141/HI io_out[7] sky130_fd_sc_hd__conb_1
XFILLER_26_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2528__A _2528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_20_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2711_ _2712_/A _2712_/B _2712_/C vssd1 vssd1 vccd1 vccd1 _2783_/A sky130_fd_sc_hd__o21ai_2
XFILLER_9_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2642_ _2642_/A _2642_/B _2642_/C vssd1 vssd1 vccd1 vccd1 _2653_/A sky130_fd_sc_hd__and3_1
X_2573_ _2573_/A _2573_/B _2573_/C vssd1 vssd1 vccd1 vccd1 _2573_/Y sky130_fd_sc_hd__nand3_1
X_1524_ _1524_/A _1524_/B vssd1 vssd1 vccd1 vccd1 _1525_/B sky130_fd_sc_hd__nor2_1
XFILLER_28_618 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_55_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2007_ _2000_/A _2000_/B _2006_/X vssd1 vssd1 vccd1 vccd1 _2057_/A sky130_fd_sc_hd__a21bo_1
XFILLER_63_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_50_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2909_ _2909_/A _2909_/B vssd1 vssd1 vccd1 vccd1 _2909_/X sky130_fd_sc_hd__or2_1
XANTENNA__2901__A _2901_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_40 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_84 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2811__A _2919_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_64_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_212 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2625_ _2624_/A _2624_/B _2624_/C vssd1 vssd1 vccd1 vccd1 _2640_/B sky130_fd_sc_hd__a21oi_2
X_2556_ _2556_/A vssd1 vssd1 vccd1 vccd1 _2824_/A sky130_fd_sc_hd__clkbuf_4
X_1507_ _1507_/A _1507_/B _1505_/Y vssd1 vssd1 vccd1 vccd1 _1508_/B sky130_fd_sc_hd__or3b_1
X_2487_ _2488_/A _2488_/B vssd1 vssd1 vccd1 vccd1 _2583_/B sky130_fd_sc_hd__nand2_1
XFILLER_55_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3159__253 vssd1 vssd1 vccd1 vccd1 _3159__253/HI la_data_out[110] sky130_fd_sc_hd__conb_1
XFILLER_11_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_46_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput36 la_data_in[41] vssd1 vssd1 vccd1 vccd1 _2120_/A sky130_fd_sc_hd__clkbuf_1
Xinput14 la_data_in[21] vssd1 vssd1 vccd1 vccd1 _2023_/A sky130_fd_sc_hd__clkbuf_2
Xinput25 la_data_in[31] vssd1 vssd1 vccd1 vccd1 _2629_/B sky130_fd_sc_hd__buf_4
Xinput47 la_data_in[51] vssd1 vssd1 vccd1 vccd1 _2797_/A sky130_fd_sc_hd__buf_2
Xinput58 la_data_in[61] vssd1 vssd1 vccd1 vccd1 _1720_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2410_ _2410_/A vssd1 vssd1 vccd1 vccd1 _2686_/A sky130_fd_sc_hd__clkbuf_2
X_2341_ _2071_/A _1943_/A _1947_/A _2416_/A vssd1 vssd1 vccd1 vccd1 _2341_/X sky130_fd_sc_hd__a22o_1
X_2272_ _2272_/A _2272_/B vssd1 vssd1 vccd1 vccd1 _2283_/A sky130_fd_sc_hd__and2_1
XFILLER_28_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_440 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1987_ _1987_/A vssd1 vssd1 vccd1 vccd1 _1988_/A sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__2401__A1 _2528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2608_ _2608_/A vssd1 vssd1 vccd1 vccd1 _2936_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_0_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2539_ _2539_/A vssd1 vssd1 vccd1 vccd1 _2811_/C sky130_fd_sc_hd__clkbuf_2
XFILLER_57_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_418 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_484 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2957__A2_N _2958_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input52_A la_data_in[56] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_3_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_34_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1910_ _1910_/A _1963_/A _1910_/C vssd1 vssd1 vccd1 vccd1 _1912_/A sky130_fd_sc_hd__and3_1
X_2890_ _2908_/A _2908_/B vssd1 vssd1 vccd1 vccd1 _2892_/B sky130_fd_sc_hd__xor2_1
X_1841_ _1841_/A _1850_/B vssd1 vssd1 vccd1 vccd1 _1848_/B sky130_fd_sc_hd__xor2_1
XFILLER_30_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2271__A _2271_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1772_ input8/X vssd1 vssd1 vccd1 vccd1 _1800_/A sky130_fd_sc_hd__clkbuf_2
X_2324_ _2325_/B _2461_/A _2458_/A vssd1 vssd1 vccd1 vccd1 _2378_/A sky130_fd_sc_hd__o21ai_1
X_2255_ _2255_/A _2321_/A vssd1 vssd1 vccd1 vccd1 _2258_/A sky130_fd_sc_hd__xnor2_4
X_2186_ _2079_/A _2189_/A _2137_/A vssd1 vssd1 vccd1 vccd1 _2192_/B sky130_fd_sc_hd__o21ai_2
XFILLER_38_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2446__A _2447_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_53_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_53_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3080__174 vssd1 vssd1 vccd1 vccd1 _3080__174/HI irq[2] sky130_fd_sc_hd__conb_1
XANTENNA__2622__A1 _2026_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2925__A2 _2921_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_130 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_229 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_218 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_207 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2040_ _2612_/A _2040_/B vssd1 vssd1 vccd1 vccd1 _2069_/A sky130_fd_sc_hd__xnor2_2
X_3064__158 vssd1 vssd1 vccd1 vccd1 _3064__158/HI io_out[24] sky130_fd_sc_hd__conb_1
XFILLER_62_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2942_ _2942_/A _2989_/A vssd1 vssd1 vccd1 vccd1 _2943_/B sky130_fd_sc_hd__xor2_2
XFILLER_15_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3105__199 vssd1 vssd1 vccd1 vccd1 _3105__199/HI la_data_out[24] sky130_fd_sc_hd__conb_1
X_2873_ _2037_/X _2871_/Y _2872_/X vssd1 vssd1 vccd1 vccd1 _2874_/B sky130_fd_sc_hd__a21o_1
X_1824_ _2130_/A _1984_/A _1821_/X _1823_/Y vssd1 vssd1 vccd1 vccd1 _1837_/A sky130_fd_sc_hd__a211o_1
X_1755_ _1718_/B _1752_/X _1754_/Y _1740_/B vssd1 vssd1 vccd1 vccd1 _1763_/A sky130_fd_sc_hd__o22a_2
X_1686_ _1714_/A _1686_/B vssd1 vssd1 vccd1 vccd1 _1688_/B sky130_fd_sc_hd__and2b_1
XTAP_752 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_741 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_730 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_785 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_774 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_763 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2307_ _2307_/A _2307_/B vssd1 vssd1 vccd1 vccd1 _2450_/A sky130_fd_sc_hd__or2_2
XTAP_796 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2238_ _2238_/A _2238_/B vssd1 vssd1 vccd1 vccd1 _2240_/B sky130_fd_sc_hd__xnor2_1
XFILLER_26_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_310 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2169_ _2235_/C _2169_/B vssd1 vssd1 vccd1 vccd1 _2170_/B sky130_fd_sc_hd__xnor2_1
XFILLER_41_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2531__B1 _2766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_input15_A la_data_in[22] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2086__A _2086_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2834__A1 _2884_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2598__B1 _2597_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2533__B _2629_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_1540_ _2932_/B _2965_/B vssd1 vssd1 vccd1 vccd1 _1540_/Y sky130_fd_sc_hd__nor2_1
XFILLER_5_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA_output83_A _2730_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2023_ _2023_/A _2023_/B vssd1 vssd1 vccd1 vccd1 _2024_/A sky130_fd_sc_hd__xnor2_1
XFILLER_23_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2925_ _2819_/A _2921_/X _2924_/Y vssd1 vssd1 vccd1 vccd1 _2926_/B sky130_fd_sc_hd__o21a_1
X_2856_ _2856_/A _2856_/B vssd1 vssd1 vccd1 vccd1 _2856_/X sky130_fd_sc_hd__xor2_2
X_1807_ _1807_/A _1839_/A _1807_/C vssd1 vssd1 vccd1 vccd1 _1848_/A sky130_fd_sc_hd__or3_1
X_2787_ _2805_/A _2805_/B vssd1 vssd1 vccd1 vccd1 _2789_/B sky130_fd_sc_hd__xnor2_2
X_1738_ _1738_/A _1738_/B _1738_/C vssd1 vssd1 vccd1 vccd1 _1739_/B sky130_fd_sc_hd__and3_1
X_3192__286 vssd1 vssd1 vccd1 vccd1 _3192__286/HI wbs_dat_o[14] sky130_fd_sc_hd__conb_1
X_1669_ input4/X _2983_/A _1669_/S vssd1 vssd1 vccd1 vccd1 _1671_/B sky130_fd_sc_hd__mux2_1
XFILLER_49_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input7_A la_data_in[15] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_560 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_582 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_571 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_593 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3086__180 vssd1 vssd1 vccd1 vccd1 _3086__180/HI la_data_out[5] sky130_fd_sc_hd__conb_1
XFILLER_26_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_302 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_5_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_57_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_118 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1491__B1 _1488_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2544__A _2544_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2710_ _2710_/A _2710_/B vssd1 vssd1 vccd1 vccd1 _2712_/C sky130_fd_sc_hd__or2_2
X_2641_ _2712_/B _2640_/B _2640_/C vssd1 vssd1 vccd1 vccd1 _2642_/C sky130_fd_sc_hd__o21ai_1
XFILLER_58_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2572_ _2645_/A _2645_/B vssd1 vssd1 vccd1 vccd1 _2573_/C sky130_fd_sc_hd__xor2_2
X_1523_ _1522_/B _1523_/B vssd1 vssd1 vccd1 vccd1 _1524_/B sky130_fd_sc_hd__and2b_1
XFILLER_4_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2006_ _2006_/A _2008_/B _2006_/C vssd1 vssd1 vccd1 vccd1 _2006_/X sky130_fd_sc_hd__or3_1
XFILLER_63_460 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3120__214 vssd1 vssd1 vccd1 vccd1 _3120__214/HI la_data_out[39] sky130_fd_sc_hd__conb_1
X_2908_ _2908_/A _2908_/B vssd1 vssd1 vccd1 vccd1 _2949_/A sky130_fd_sc_hd__nor2_1
X_2839_ _2026_/Y _2880_/A _2966_/A _2568_/X vssd1 vssd1 vccd1 vccd1 _2840_/B sky130_fd_sc_hd__a22o_1
XANTENNA__1537__A1 _1521_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2734__B1 _2766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1533__A _1533_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2629__A _2629_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_390 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_25_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_41_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_176 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_482 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2274__A input5/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2624_ _2624_/A _2624_/B _2624_/C vssd1 vssd1 vccd1 vccd1 _2712_/B sky130_fd_sc_hd__and3_2
X_2555_ _2612_/A _2555_/B vssd1 vssd1 vccd1 vccd1 _2644_/A sky130_fd_sc_hd__xnor2_2
X_1506_ _1507_/A _1507_/B _1505_/Y vssd1 vssd1 vccd1 vccd1 _1561_/A sky130_fd_sc_hd__o21ba_4
X_2486_ _2623_/A _2486_/B vssd1 vssd1 vccd1 vccd1 _2488_/B sky130_fd_sc_hd__xnor2_1
XFILLER_28_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2247__A2 _2185_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_51_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3198__292 vssd1 vssd1 vccd1 vccd1 _3198__292/HI wbs_dat_o[20] sky130_fd_sc_hd__conb_1
XFILLER_11_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_19_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2078__B _2138_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_46_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_246 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_42_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput26 la_data_in[32] vssd1 vssd1 vccd1 vccd1 _1775_/C sky130_fd_sc_hd__clkbuf_1
Xinput15 la_data_in[22] vssd1 vssd1 vccd1 vccd1 _2023_/B sky130_fd_sc_hd__buf_2
Xinput37 la_data_in[42] vssd1 vssd1 vccd1 vccd1 _2242_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput48 la_data_in[52] vssd1 vssd1 vccd1 vccd1 _2901_/A sky130_fd_sc_hd__clkbuf_4
Xinput59 la_data_in[62] vssd1 vssd1 vccd1 vccd1 _1745_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_2340_ _2556_/A _2340_/B vssd1 vssd1 vccd1 vccd1 _2345_/A sky130_fd_sc_hd__xnor2_1
XFILLER_2_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2271_ _2271_/A _2271_/B vssd1 vssd1 vccd1 vccd1 _2272_/B sky130_fd_sc_hd__or2_1
XFILLER_52_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_282 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1986_ _2036_/B _2927_/B vssd1 vssd1 vccd1 vccd1 _1987_/A sky130_fd_sc_hd__and2_1
XANTENNA__2401__A2 _2400_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2607_ _2739_/A _2979_/A _2979_/B vssd1 vssd1 vccd1 vccd1 _2614_/B sky130_fd_sc_hd__or3_2
X_2538_ _2538_/A _2921_/A _2921_/B vssd1 vssd1 vccd1 vccd1 _2543_/B sky130_fd_sc_hd__or3_4
XANTENNA__2179__A _2179_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2469_ _2469_/A vssd1 vssd1 vccd1 vccd1 _2747_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_28_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3126__220 vssd1 vssd1 vccd1 vccd1 _3126__220/HI la_data_out[45] sky130_fd_sc_hd__conb_1
XFILLER_24_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_496 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2928__A0 _1944_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_3_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input45_A la_data_in[4] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1840_ _2329_/A _1839_/B _1839_/Y vssd1 vssd1 vccd1 vccd1 _1850_/B sky130_fd_sc_hd__a21o_1
XFILLER_30_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_30_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1771_ _2454_/A vssd1 vssd1 vccd1 vccd1 _2393_/A sky130_fd_sc_hd__buf_2
XFILLER_6_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2323_ _2462_/A _2323_/B vssd1 vssd1 vccd1 vccd1 _2458_/A sky130_fd_sc_hd__and2_1
X_2254_ _2254_/A vssd1 vssd1 vccd1 vccd1 _2636_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_38_522 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2185_ input5/X _2185_/B vssd1 vssd1 vccd1 vccd1 _2199_/A sky130_fd_sc_hd__xnor2_1
XFILLER_38_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_455 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1969_ _2137_/A vssd1 vssd1 vccd1 vccd1 _2416_/A sky130_fd_sc_hd__buf_2
XFILLER_4_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_219 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_208 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_514 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2941_ _2941_/A _2985_/B vssd1 vssd1 vccd1 vccd1 _2989_/A sky130_fd_sc_hd__xor2_2
XFILLER_50_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2872_ _2697_/A _2550_/X _2609_/X _2922_/A vssd1 vssd1 vccd1 vccd1 _2872_/X sky130_fd_sc_hd__a22o_1
X_1823_ _2181_/A _2034_/A _2134_/B vssd1 vssd1 vccd1 vccd1 _1823_/Y sky130_fd_sc_hd__a21oi_1
X_1754_ _1754_/A _1754_/B vssd1 vssd1 vccd1 vccd1 _1754_/Y sky130_fd_sc_hd__nor2_1
XFILLER_7_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_7_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1591__A2 _1548_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1685_ _1685_/A _1685_/B vssd1 vssd1 vccd1 vccd1 _1686_/B sky130_fd_sc_hd__or2_1
XTAP_742 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_731 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_720 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_786 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_775 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_764 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_753 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2306_ _2365_/A vssd1 vssd1 vccd1 vccd1 _2306_/Y sky130_fd_sc_hd__inv_2
XTAP_797 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_57_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2237_ _2170_/A _2235_/X _2236_/X vssd1 vssd1 vccd1 vccd1 _2238_/B sky130_fd_sc_hd__a21o_1
XFILLER_54_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2168_ _2235_/A _2235_/B vssd1 vssd1 vccd1 vccd1 _2169_/B sky130_fd_sc_hd__nor2_1
XFILLER_26_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2099_ _2099_/A vssd1 vssd1 vccd1 vccd1 _2560_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_21_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2834__A2 _2833_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3031__125 vssd1 vssd1 vccd1 vccd1 _3031__125/HI io_oeb[28] sky130_fd_sc_hd__conb_1
XFILLER_39_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2022_ _2022_/A vssd1 vssd1 vccd1 vccd1 _2194_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_35_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2924_ _2740_/X _2820_/X _2923_/X vssd1 vssd1 vccd1 vccd1 _2924_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_31_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2855_ _2728_/A _2728_/B _2801_/A _2854_/X vssd1 vssd1 vccd1 vccd1 _2856_/B sky130_fd_sc_hd__a31o_1
X_1806_ _1899_/A _1807_/C _1839_/B _1839_/A vssd1 vssd1 vccd1 vccd1 _1806_/Y sky130_fd_sc_hd__o211ai_1
X_2786_ _2715_/A _2715_/B _2716_/B _2716_/A vssd1 vssd1 vccd1 vccd1 _2805_/B sky130_fd_sc_hd__o22a_1
X_1737_ _1738_/A _1738_/B _1738_/C vssd1 vssd1 vccd1 vccd1 _1739_/A sky130_fd_sc_hd__a21oi_1
X_1668_ _1761_/A _2349_/B vssd1 vssd1 vccd1 vccd1 _1669_/S sky130_fd_sc_hd__nand2_1
X_1599_ _1600_/B _1599_/B vssd1 vssd1 vccd1 vccd1 _1601_/A sky130_fd_sc_hd__and2b_1
XTAP_550 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_561 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_583 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_572 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_594 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3015__109 vssd1 vssd1 vccd1 vccd1 _3015__109/HI io_oeb[12] sky130_fd_sc_hd__conb_1
XFILLER_1_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_487 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_49_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_94 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1491__B2 _1488_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1491__A1 _2954_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_13_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2640_ _2712_/B _2640_/B _2640_/C vssd1 vssd1 vccd1 vccd1 _2642_/B sky130_fd_sc_hd__or3_1
X_2571_ _2862_/A _2571_/B vssd1 vssd1 vccd1 vccd1 _2645_/B sky130_fd_sc_hd__xnor2_2
X_1522_ _1523_/B _1522_/B vssd1 vssd1 vccd1 vccd1 _1524_/A sky130_fd_sc_hd__and2b_1
XFILLER_4_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2005_ _2005_/A _2005_/B vssd1 vssd1 vccd1 vccd1 _2005_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_51_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2907_ _2804_/A _2905_/B _2905_/X _2906_/Y vssd1 vssd1 vccd1 vccd1 _2952_/A sky130_fd_sc_hd__o211a_2
X_3200__294 vssd1 vssd1 vccd1 vccd1 _3200__294/HI wbs_dat_o[22] sky130_fd_sc_hd__conb_1
X_2838_ _2686_/X _2913_/B _2772_/A _2567_/X vssd1 vssd1 vccd1 vccd1 _2840_/A sky130_fd_sc_hd__a22o_1
X_2769_ _2768_/A _2768_/B _2768_/C vssd1 vssd1 vccd1 vccd1 _2779_/B sky130_fd_sc_hd__a21oi_1
XFILLER_2_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2734__A1 _2703_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_4_9 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1533__B _1533_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2629__B _2629_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_380 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_391 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_480 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_75 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_1_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_49_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_49_266 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3143__237 vssd1 vssd1 vccd1 vccd1 _3143__237/HI la_data_out[62] sky130_fd_sc_hd__conb_1
XFILLER_17_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2274__B input4/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2623_ _2623_/A _2623_/B vssd1 vssd1 vccd1 vccd1 _2624_/C sky130_fd_sc_hd__xnor2_1
X_3037__131 vssd1 vssd1 vccd1 vccd1 _3037__131/HI io_oeb[34] sky130_fd_sc_hd__conb_1
X_2554_ _2554_/A _2554_/B vssd1 vssd1 vccd1 vccd1 _2555_/B sky130_fd_sc_hd__nor2_1
X_1505_ _1505_/A _1505_/B vssd1 vssd1 vccd1 vccd1 _1505_/Y sky130_fd_sc_hd__nor2_1
X_2485_ _1929_/Y _2684_/A _2756_/A _2404_/X _2484_/X vssd1 vssd1 vccd1 vccd1 _2486_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_28_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_450 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_51_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_199 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_3_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_269 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_483 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_27_494 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
Xinput27 la_data_in[33] vssd1 vssd1 vccd1 vccd1 _1784_/A sky130_fd_sc_hd__clkbuf_1
Xinput16 la_data_in[23] vssd1 vssd1 vccd1 vccd1 _2138_/A sky130_fd_sc_hd__buf_2
Xinput38 la_data_in[43] vssd1 vssd1 vccd1 vccd1 _2240_/A sky130_fd_sc_hd__dlymetal6s2s_1
Xinput49 la_data_in[53] vssd1 vssd1 vccd1 vccd1 _2956_/A sky130_fd_sc_hd__buf_2
XFILLER_6_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1921__A2 _2410_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2270_ _2271_/A _2271_/B vssd1 vssd1 vccd1 vccd1 _2272_/A sky130_fd_sc_hd__nand2_1
XFILLER_37_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1985_ _1898_/A _1985_/B vssd1 vssd1 vccd1 vccd1 _2927_/B sky130_fd_sc_hd__and2b_1
XFILLER_20_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2606_ _2573_/A _2573_/C _2573_/B vssd1 vssd1 vccd1 vccd1 _2642_/A sky130_fd_sc_hd__a21bo_1
X_2537_ _2694_/A _2536_/B _2536_/C vssd1 vssd1 vccd1 vccd1 _2921_/B sky130_fd_sc_hd__a21oi_1
X_2468_ _2536_/B _2468_/B vssd1 vssd1 vccd1 vccd1 _2468_/Y sky130_fd_sc_hd__nand2_4
X_2399_ _2399_/A _2399_/B _2399_/C vssd1 vssd1 vccd1 vccd1 _2400_/C sky130_fd_sc_hd__nand3_4
XFILLER_24_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_11_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input38_A la_data_in[43] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_420 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2092__A1 _1929_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2833__A _2884_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_423 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_283 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1770_ _2313_/S vssd1 vssd1 vccd1 vccd1 _2454_/A sky130_fd_sc_hd__clkbuf_1
XFILLER_6_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2322_ _2322_/A _2322_/B vssd1 vssd1 vccd1 vccd1 _2323_/B sky130_fd_sc_hd__or2_1
XFILLER_33_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2253_ _2130_/X _2469_/A _2250_/X _2252_/Y vssd1 vssd1 vccd1 vccd1 _2262_/A sky130_fd_sc_hd__a211o_2
XFILLER_38_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3149__243 vssd1 vssd1 vccd1 vccd1 _3149__243/HI la_data_out[100] sky130_fd_sc_hd__conb_1
X_2184_ _2130_/A _2134_/C _2181_/X _2183_/Y vssd1 vssd1 vccd1 vccd1 _2185_/B sky130_fd_sc_hd__a211o_2
XFILLER_38_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_38_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_467 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1968_ _1968_/A _1968_/B _1968_/C vssd1 vssd1 vccd1 vccd1 _1968_/X sky130_fd_sc_hd__and3_1
X_1899_ _1899_/A _2036_/A vssd1 vssd1 vccd1 vccd1 _1900_/B sky130_fd_sc_hd__nand2_1
XFILLER_48_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_272 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_209 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2828__A _2965_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_35_526 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_62_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2940_ _2963_/A _2963_/B vssd1 vssd1 vccd1 vccd1 _2985_/B sky130_fd_sc_hd__xor2_4
XFILLER_50_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2563__A _2824_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2871_ _2922_/A _2694_/X _2630_/D _2695_/Y vssd1 vssd1 vccd1 vccd1 _2871_/Y sky130_fd_sc_hd__a211oi_4
XFILLER_43_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1822_ _1968_/A vssd1 vssd1 vccd1 vccd1 _2181_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_1753_ _1753_/A vssd1 vssd1 vccd1 vccd1 _1754_/A sky130_fd_sc_hd__inv_2
X_1684_ _1685_/A _1685_/B vssd1 vssd1 vccd1 vccd1 _1714_/A sky130_fd_sc_hd__and2_1
XTAP_710 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_743 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_732 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_721 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_776 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_765 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_754 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2305_ _2305_/A _2305_/B vssd1 vssd1 vccd1 vccd1 _2365_/A sky130_fd_sc_hd__nand2_1
XTAP_798 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_787 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2236_ _2235_/A _2235_/B _2235_/C vssd1 vssd1 vccd1 vccd1 _2236_/X sky130_fd_sc_hd__o21a_1
X_2167_ _2233_/C _2233_/D vssd1 vssd1 vccd1 vccd1 _2235_/C sky130_fd_sc_hd__xnor2_1
X_2098_ _2206_/A _2148_/B vssd1 vssd1 vccd1 vccd1 _2099_/A sky130_fd_sc_hd__nor2_1
XFILLER_13_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__1536__B _2986_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_179 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_331 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_375 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_44_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_8_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_286 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3070__164 vssd1 vssd1 vccd1 vccd1 _3070__164/HI io_out[30] sky130_fd_sc_hd__conb_1
XFILLER_39_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2021_ _2021_/A vssd1 vssd1 vccd1 vccd1 _2568_/A sky130_fd_sc_hd__buf_2
XFILLER_63_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_120 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2038__A1 _1888_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_50_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2923_ _2922_/X _2748_/X _2749_/X _2814_/X vssd1 vssd1 vccd1 vccd1 _2923_/X sky130_fd_sc_hd__a22o_1
X_2854_ _2723_/A _2723_/B _2799_/B _2797_/X vssd1 vssd1 vccd1 vccd1 _2854_/X sky130_fd_sc_hd__a31o_1
XFILLER_31_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1805_ _2134_/B _1805_/B vssd1 vssd1 vccd1 vccd1 _1807_/C sky130_fd_sc_hd__nand2_1
X_2785_ _2785_/A _2785_/B vssd1 vssd1 vccd1 vccd1 _2805_/A sky130_fd_sc_hd__nand2_1
X_1736_ _1736_/A _1736_/B vssd1 vssd1 vccd1 vccd1 _1738_/C sky130_fd_sc_hd__xnor2_1
X_1667_ _1726_/A _1667_/B vssd1 vssd1 vccd1 vccd1 _1675_/A sky130_fd_sc_hd__and2_1
X_1598_ _1641_/A _1598_/B vssd1 vssd1 vccd1 vccd1 _1599_/B sky130_fd_sc_hd__and2_1
XTAP_540 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_551 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_426 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_562 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_584 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_573 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_595 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2219_ _2219_/A _2219_/B vssd1 vssd1 vccd1 vccd1 _2220_/C sky130_fd_sc_hd__nor2_1
XFILLER_53_142 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2931__A _2931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_30_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3054__148 vssd1 vssd1 vccd1 vccd1 _3054__148/HI io_out[14] sky130_fd_sc_hd__conb_1
XFILLER_1_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_52 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input20_A la_data_in[27] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2268__A1 _1929_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_29_150 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1491__A2 _2954_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_370 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_599 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2570_ _2402_/X _2756_/A _2566_/Y _2569_/X vssd1 vssd1 vccd1 vccd1 _2571_/B sky130_fd_sc_hd__a211o_1
X_1521_ _1521_/A _1521_/B vssd1 vssd1 vccd1 vccd1 _1522_/B sky130_fd_sc_hd__xor2_1
XFILLER_36_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2004_ _1959_/X _1962_/B _1960_/A vssd1 vssd1 vccd1 vccd1 _2005_/B sky130_fd_sc_hd__a21o_1
XFILLER_23_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2454__C _2629_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2906_ _2892_/A _2851_/B _2892_/B vssd1 vssd1 vccd1 vccd1 _2906_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_50_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2837_ _2858_/B _2837_/B vssd1 vssd1 vccd1 vccd1 _2845_/A sky130_fd_sc_hd__xnor2_2
X_2768_ _2768_/A _2768_/B _2768_/C vssd1 vssd1 vccd1 vccd1 _2808_/A sky130_fd_sc_hd__and3_1
X_1719_ _1720_/A _1720_/B vssd1 vssd1 vccd1 vccd1 _1721_/A sky130_fd_sc_hd__and2_1
X_2699_ _2922_/A _2811_/C vssd1 vssd1 vccd1 vccd1 _2702_/D sky130_fd_sc_hd__nand2_1
XANTENNA__2734__A2 _2703_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2498__A1 input6/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_370 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_381 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_392 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2926__A _2926_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_18_109 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_492 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_10 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_495 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_10_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2380__B _2380_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_64 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_6_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3182__276 vssd1 vssd1 vccd1 vccd1 _3182__276/HI wbs_dat_o[4] sky130_fd_sc_hd__conb_1
XFILLER_32_112 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2413__A1 _2026_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2413__B2 _2568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2622_ _2026_/Y _2684_/A _2756_/A _2568_/X _2621_/X vssd1 vssd1 vccd1 vccd1 _2623_/B
+ sky130_fd_sc_hd__a221o_1
X_3076__170 vssd1 vssd1 vccd1 vccd1 _3076__170/HI io_out[36] sky130_fd_sc_hd__conb_1
X_2553_ _2037_/X _2931_/A _2931_/B _2609_/A _2863_/A vssd1 vssd1 vccd1 vccd1 _2554_/B
+ sky130_fd_sc_hd__a32o_1
X_1504_ _2258_/Y _2880_/X _2966_/X _2913_/A vssd1 vssd1 vccd1 vccd1 _1505_/B sky130_fd_sc_hd__a22o_1
X_2484_ _2568_/A _2347_/A _2403_/A _2402_/A vssd1 vssd1 vccd1 vccd1 _2484_/X sky130_fd_sc_hd__a22o_1
XANTENNA__2746__A _2824_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_602 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_23_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_454 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xinput28 la_data_in[34] vssd1 vssd1 vccd1 vccd1 _1810_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__1719__B _1720_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xinput17 la_data_in[24] vssd1 vssd1 vccd1 vccd1 _2188_/A sky130_fd_sc_hd__buf_2
Xinput39 la_data_in[44] vssd1 vssd1 vccd1 vccd1 _2299_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_3110__204 vssd1 vssd1 vccd1 vccd1 _3110__204/HI la_data_out[29] sky130_fd_sc_hd__conb_1
XFILLER_37_204 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2566__A _2775_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_60_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1984_ _1984_/A vssd1 vssd1 vccd1 vccd1 _2404_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_9_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2605_ _2528_/Y _2529_/X _2573_/Y _2574_/X vssd1 vssd1 vccd1 vccd1 _2605_/X sky130_fd_sc_hd__o211a_1
XFILLER_0_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2536_ _2694_/A _2536_/B _2536_/C vssd1 vssd1 vccd1 vccd1 _2921_/A sky130_fd_sc_hd__and3_1
X_2467_ _2467_/A _2467_/B _2467_/C vssd1 vssd1 vccd1 vccd1 _2468_/B sky130_fd_sc_hd__nand3_1
X_2398_ _2399_/B _2399_/C _2399_/A vssd1 vssd1 vccd1 vccd1 _2528_/A sky130_fd_sc_hd__a21o_2
XFILLER_28_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_47_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2833__B _2833_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_295 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2321_ _2321_/A _2380_/A vssd1 vssd1 vccd1 vccd1 _2462_/A sky130_fd_sc_hd__nand2_1
X_2252_ _2454_/A _2385_/A _2454_/B vssd1 vssd1 vccd1 vccd1 _2252_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_26_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3188__282 vssd1 vssd1 vccd1 vccd1 _3188__282/HI wbs_dat_o[10] sky130_fd_sc_hd__conb_1
X_2183_ _2181_/A _2469_/A _2134_/B vssd1 vssd1 vccd1 vccd1 _2183_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_53_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_549 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1967_ _2137_/A vssd1 vssd1 vccd1 vccd1 _1968_/C sky130_fd_sc_hd__clkbuf_2
X_1898_ _1898_/A vssd1 vssd1 vccd1 vccd1 _2036_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_2519_ _2600_/A _2519_/B vssd1 vssd1 vccd1 vccd1 _2522_/A sky130_fd_sc_hd__nor2_1
XFILLER_56_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_56_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_590 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input50_A la_data_in[54] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_35_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2870_ _2976_/A _2870_/B vssd1 vssd1 vccd1 vccd1 _2911_/A sky130_fd_sc_hd__xnor2_4
X_1821_ _1821_/A _1968_/B _2034_/A vssd1 vssd1 vccd1 vccd1 _1821_/X sky130_fd_sc_hd__and3_1
XFILLER_30_232 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_30_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1752_ _1753_/A _1740_/B _1741_/B vssd1 vssd1 vccd1 vccd1 _1752_/X sky130_fd_sc_hd__a21o_1
X_1683_ _1597_/A _1597_/B _1641_/B _1640_/B _1640_/A vssd1 vssd1 vccd1 vccd1 _1685_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_7_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3116__210 vssd1 vssd1 vccd1 vccd1 _3116__210/HI la_data_out[35] sky130_fd_sc_hd__conb_1
XTAP_700 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_733 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_722 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_711 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_777 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_766 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_755 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_744 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2304_ _2297_/S _2294_/A _2294_/B vssd1 vssd1 vccd1 vccd1 _2367_/A sky130_fd_sc_hd__o21ba_1
XTAP_799 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_788 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2235_ _2235_/A _2235_/B _2235_/C vssd1 vssd1 vccd1 vccd1 _2235_/X sky130_fd_sc_hd__or3_1
X_2166_ _2176_/A _2176_/B vssd1 vssd1 vccd1 vccd1 _2233_/D sky130_fd_sc_hd__xor2_2
XFILLER_53_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2097_ _2097_/A _2097_/B vssd1 vssd1 vccd1 vccd1 _2148_/B sky130_fd_sc_hd__xnor2_1
XFILLER_21_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2999_ _2999_/A _2999_/B vssd1 vssd1 vccd1 vccd1 _2999_/X sky130_fd_sc_hd__or2_2
XANTENNA__1536__C _1555_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1833__A input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_387 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2383__B _2931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_44_97 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_8_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2020_ _2020_/A vssd1 vssd1 vccd1 vccd1 _2021_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_35_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2922_ _2922_/A vssd1 vssd1 vccd1 vccd1 _2922_/X sky130_fd_sc_hd__clkbuf_2
XFILLER_31_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2853_ _2901_/A _2901_/B vssd1 vssd1 vccd1 vccd1 _2856_/A sky130_fd_sc_hd__xor2_2
XFILLER_31_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1804_ _1968_/B vssd1 vssd1 vccd1 vccd1 _2134_/B sky130_fd_sc_hd__clkbuf_2
X_2784_ _2783_/B _2783_/C _2783_/A vssd1 vssd1 vccd1 vccd1 _2785_/B sky130_fd_sc_hd__o21ai_1
X_1735_ _1756_/A _1756_/B vssd1 vssd1 vccd1 vccd1 _1736_/B sky130_fd_sc_hd__xor2_1
X_1666_ _1666_/A _1666_/B _1666_/C vssd1 vssd1 vccd1 vccd1 _1667_/B sky130_fd_sc_hd__or3_1
X_1597_ _1597_/A _1597_/B vssd1 vssd1 vccd1 vccd1 _1598_/B sky130_fd_sc_hd__or2_1
XTAP_530 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_541 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_552 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_563 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_585 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_574 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_596 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2218_ _2217_/B _2218_/B vssd1 vssd1 vccd1 vccd1 _2219_/B sky130_fd_sc_hd__and2b_1
X_2149_ _2206_/B _2149_/B vssd1 vssd1 vccd1 vccd1 _2150_/A sky130_fd_sc_hd__and2_1
XFILLER_53_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_41_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2931__B _2931_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_5_206 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3093__187 vssd1 vssd1 vccd1 vccd1 _3093__187/HI la_data_out[12] sky130_fd_sc_hd__conb_1
XFILLER_1_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_471 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_162 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_45_611 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input13_A la_data_in[20] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_154 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_32_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_382 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1520_ _1555_/B _1520_/B vssd1 vssd1 vccd1 vccd1 _1521_/B sky130_fd_sc_hd__xnor2_1
XFILLER_4_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2003_ _2003_/A _2002_/X vssd1 vssd1 vccd1 vccd1 _2005_/A sky130_fd_sc_hd__or2b_1
XFILLER_63_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_23_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2905_ _2905_/A _2905_/B vssd1 vssd1 vccd1 vccd1 _2905_/X sky130_fd_sc_hd__or2_1
X_2836_ _2836_/A _2836_/B vssd1 vssd1 vccd1 vccd1 _2837_/B sky130_fd_sc_hd__xor2_2
X_2767_ _2705_/A _2705_/B _2766_/Y _2674_/A vssd1 vssd1 vccd1 vccd1 _2768_/C sky130_fd_sc_hd__a22o_1
X_1718_ _1718_/A _1718_/B vssd1 vssd1 vccd1 vccd1 _1720_/B sky130_fd_sc_hd__xnor2_4
X_2698_ _2810_/A _2698_/B vssd1 vssd1 vccd1 vccd1 _2702_/C sky130_fd_sc_hd__nand2_1
X_1649_ _1649_/A _1659_/A vssd1 vssd1 vccd1 vccd1 _1649_/Y sky130_fd_sc_hd__nor2_1
XFILLER_58_224 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input5_A la_data_in[13] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_360 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_371 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_382 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_393 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XPHY_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_22 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_54_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3021__115 vssd1 vssd1 vccd1 vccd1 _3021__115/HI io_oeb[18] sky130_fd_sc_hd__conb_1
XFILLER_10_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2621_ _2686_/A _2685_/A _2757_/A _2567_/A vssd1 vssd1 vccd1 vccd1 _2621_/X sky130_fd_sc_hd__a22o_1
XFILLER_56_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2552_ _2552_/A vssd1 vssd1 vccd1 vccd1 _2863_/A sky130_fd_sc_hd__clkbuf_2
X_1503_ _2936_/X _1502_/X _2772_/X _2863_/X vssd1 vssd1 vccd1 vccd1 _1505_/A sky130_fd_sc_hd__a22o_1
X_2483_ _2483_/A vssd1 vssd1 vccd1 vccd1 _2756_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_55_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_24_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2762__A _2843_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_23_157 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2819_ _2819_/A _2979_/A _2979_/B vssd1 vssd1 vccd1 vccd1 _2824_/B sky130_fd_sc_hd__or3_1
XFILLER_11_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_190 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_21 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_36_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_400 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_42_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_53 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xinput18 la_data_in[25] vssd1 vssd1 vccd1 vccd1 _2188_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_6_323 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3099__193 vssd1 vssd1 vccd1 vccd1 _3099__193/HI la_data_out[18] sky130_fd_sc_hd__conb_1
Xinput29 la_data_in[35] vssd1 vssd1 vccd1 vccd1 _1843_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_6_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_208 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_260 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_422 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1983_ _2049_/A _2049_/B vssd1 vssd1 vccd1 vccd1 _1992_/A sky130_fd_sc_hd__xor2_1
X_2604_ _2523_/X _2515_/A _2603_/Y _2593_/X vssd1 vssd1 vccd1 vccd1 _2665_/A sky130_fd_sc_hd__a31o_1
X_2535_ _2694_/B _2535_/B vssd1 vssd1 vccd1 vccd1 _2536_/C sky130_fd_sc_hd__nand2_1
X_2466_ _2467_/A _2467_/B _2467_/C vssd1 vssd1 vccd1 vccd1 _2536_/B sky130_fd_sc_hd__a21o_1
X_2397_ _2130_/X _2814_/A _2393_/X _2396_/Y vssd1 vssd1 vccd1 vccd1 _2399_/A sky130_fd_sc_hd__a211o_1
XANTENNA__2873__A2 _2871_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1836__A _2086_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1555__B _1555_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3133__227 vssd1 vssd1 vccd1 vccd1 _3133__227/HI la_data_out[52] sky130_fd_sc_hd__conb_1
XFILLER_47_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_47_86 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3027__121 vssd1 vssd1 vccd1 vccd1 _3027__121/HI io_oeb[24] sky130_fd_sc_hd__conb_1
XFILLER_63_30 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_293 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2320_ _2189_/A _2321_/A _2255_/A vssd1 vssd1 vccd1 vccd1 _2461_/A sky130_fd_sc_hd__o21a_1
X_2251_ _2310_/A vssd1 vssd1 vccd1 vccd1 _2454_/B sky130_fd_sc_hd__dlymetal6s2s_1
XANTENNA__2577__A _2577_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_19_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2182_ _2380_/A vssd1 vssd1 vccd1 vccd1 _2469_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_53_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_230 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1966_ _2138_/A vssd1 vssd1 vccd1 vccd1 _2137_/A sky130_fd_sc_hd__clkbuf_2
X_1897_ _1897_/A _1944_/A vssd1 vssd1 vccd1 vccd1 _1898_/A sky130_fd_sc_hd__xor2_1
X_2518_ _2518_/A _2518_/B _2518_/C vssd1 vssd1 vccd1 vccd1 _2519_/B sky130_fd_sc_hd__and3_1
XFILLER_0_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2449_ _2449_/A _2449_/B vssd1 vssd1 vccd1 vccd1 _2449_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_29_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_29_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_506 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input43_A la_data_in[48] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_325 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1820_ _1979_/A vssd1 vssd1 vccd1 vccd1 _2034_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_30_244 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1751_ _1749_/A _1750_/A _1749_/B _1746_/A vssd1 vssd1 vccd1 vccd1 _1764_/A sky130_fd_sc_hd__o31a_1
XFILLER_30_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1682_ _1711_/B _1682_/B vssd1 vssd1 vccd1 vccd1 _1685_/A sky130_fd_sc_hd__nor2_1
XFILLER_7_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_701 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_734 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_723 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_712 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2303_ _2299_/X _2302_/B _2300_/A vssd1 vssd1 vccd1 vccd1 _2371_/A sky130_fd_sc_hd__a21o_1
XANTENNA__1923__B _1972_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_767 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_756 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_745 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_789 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_778 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2234_ _2234_/A _2296_/A vssd1 vssd1 vccd1 vccd1 _2238_/A sky130_fd_sc_hd__nor2_1
X_2165_ _2111_/A _2111_/B _2164_/X vssd1 vssd1 vccd1 vccd1 _2176_/B sky130_fd_sc_hd__a21o_1
XFILLER_38_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2096_ _2096_/A vssd1 vssd1 vccd1 vccd1 _2411_/A sky130_fd_sc_hd__clkbuf_2
X_2998_ _2998_/A _2998_/B vssd1 vssd1 vccd1 vccd1 _2999_/B sky130_fd_sc_hd__nor2_1
X_1949_ _2501_/A _2417_/A vssd1 vssd1 vccd1 vccd1 _1949_/Y sky130_fd_sc_hd__nor2_1
XFILLER_0_159 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_32_509 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_65 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2204__B1 _2026_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3139__233 vssd1 vssd1 vccd1 vccd1 _3139__233/HI la_data_out[58] sky130_fd_sc_hd__conb_1
XFILLER_5_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_39_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2691__B1 _2766_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_196 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_62_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2921_ _2921_/A _2921_/B vssd1 vssd1 vccd1 vccd1 _2921_/X sky130_fd_sc_hd__or2_2
XFILLER_31_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2852_ _2852_/A _2852_/B vssd1 vssd1 vccd1 vccd1 _2901_/B sky130_fd_sc_hd__xnor2_4
X_1803_ _1807_/A _1884_/A vssd1 vssd1 vccd1 vccd1 _1839_/B sky130_fd_sc_hd__nand2_1
X_2783_ _2783_/A _2783_/B _2783_/C vssd1 vssd1 vccd1 vccd1 _2785_/A sky130_fd_sc_hd__or3_1
X_1734_ _2920_/A _1700_/B _1731_/B _1704_/B vssd1 vssd1 vccd1 vccd1 _1756_/B sky130_fd_sc_hd__a31o_1
X_1665_ _1666_/B _1666_/C _1666_/A vssd1 vssd1 vccd1 vccd1 _1726_/A sky130_fd_sc_hd__o21ai_4
X_1596_ _1597_/A _1597_/B vssd1 vssd1 vccd1 vccd1 _1641_/A sky130_fd_sc_hd__nand2_1
XFILLER_58_406 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_520 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_531 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_542 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_553 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_564 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_575 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2217_ _2218_/B _2217_/B vssd1 vssd1 vccd1 vccd1 _2219_/A sky130_fd_sc_hd__and2b_1
XTAP_586 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_597 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_26_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_53_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2148_ _2044_/A _2148_/B vssd1 vssd1 vccd1 vccd1 _2149_/B sky130_fd_sc_hd__and2b_1
XFILLER_53_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2079_ _2079_/A _2137_/A vssd1 vssd1 vccd1 vccd1 _2187_/B sky130_fd_sc_hd__nor2_1
XFILLER_22_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_49_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_262 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_472 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2002_ _2002_/A _2002_/B vssd1 vssd1 vccd1 vccd1 _2002_/X sky130_fd_sc_hd__or2_1
XFILLER_63_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2904_ _2904_/A _3000_/A vssd1 vssd1 vccd1 vccd1 _2905_/B sky130_fd_sc_hd__or2_1
X_2835_ _2884_/B _2835_/B vssd1 vssd1 vccd1 vccd1 _2836_/B sky130_fd_sc_hd__nand2_1
X_2766_ _2766_/A _2766_/B vssd1 vssd1 vccd1 vccd1 _2766_/Y sky130_fd_sc_hd__nor2_1
X_1717_ _1648_/B _1688_/B _1716_/Y _1651_/B _1689_/A vssd1 vssd1 vccd1 vccd1 _1718_/B
+ sky130_fd_sc_hd__a221oi_4
X_2697_ _2697_/A vssd1 vssd1 vccd1 vccd1 _2810_/A sky130_fd_sc_hd__buf_2
X_1648_ _1716_/A _1648_/B vssd1 vssd1 vccd1 vccd1 _1651_/A sky130_fd_sc_hd__nor2_2
X_1579_ _2818_/A _2976_/A vssd1 vssd1 vccd1 vccd1 _1623_/A sky130_fd_sc_hd__nor2_2
XTAP_350 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_361 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_372 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_383 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_394 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_12 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_14_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_34 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XPHY_89 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3060__154 vssd1 vssd1 vccd1 vccd1 _3060__154/HI io_out[20] sky130_fd_sc_hd__conb_1
XFILLER_6_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3101__195 vssd1 vssd1 vccd1 vccd1 _3101__195/HI la_data_out[20] sky130_fd_sc_hd__conb_1
XFILLER_1_210 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_239 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_228 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_100 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2620_ _2620_/A _2620_/B _2620_/C vssd1 vssd1 vccd1 vccd1 _2624_/B sky130_fd_sc_hd__nand3_1
X_2551_ _2747_/A _2549_/X _2550_/X _2608_/A vssd1 vssd1 vccd1 vccd1 _2554_/A sky130_fd_sc_hd__a22o_1
X_2482_ _2577_/A _2577_/B vssd1 vssd1 vccd1 vccd1 _2488_/A sky130_fd_sc_hd__xor2_1
X_1502_ _2773_/X vssd1 vssd1 vccd1 vccd1 _1502_/X sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_49_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_291 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_464 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_36_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_3044__138 vssd1 vssd1 vccd1 vccd1 _3044__138/HI io_out[4] sky130_fd_sc_hd__conb_1
XANTENNA__2762__B _2762_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2818_ _2818_/A _2818_/B _2818_/C vssd1 vssd1 vccd1 vccd1 _2825_/B sky130_fd_sc_hd__and3_1
XFILLER_3_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2749_ _2749_/A vssd1 vssd1 vccd1 vccd1 _2749_/X sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_191 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_180 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2953__A _2954_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_42_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_14_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_87 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xinput19 la_data_in[26] vssd1 vssd1 vccd1 vccd1 _2322_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_22_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_60_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1982_ _2009_/A _1982_/B vssd1 vssd1 vccd1 vccd1 _2049_/B sky130_fd_sc_hd__xor2_1
X_2603_ _2603_/A vssd1 vssd1 vccd1 vccd1 _2603_/Y sky130_fd_sc_hd__inv_2
X_2534_ _2534_/A _2629_/A vssd1 vssd1 vccd1 vccd1 _2535_/B sky130_fd_sc_hd__or2_1
X_2465_ _2532_/A _2465_/B vssd1 vssd1 vccd1 vccd1 _2467_/C sky130_fd_sc_hd__nand2_1
X_2396_ _2393_/A _2394_/X _2919_/A vssd1 vssd1 vccd1 vccd1 _2396_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_56_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_64_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3172__266 vssd1 vssd1 vccd1 vccd1 _3172__266/HI la_data_out[123] sky130_fd_sc_hd__conb_1
XFILLER_0_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3066__160 vssd1 vssd1 vccd1 vccd1 _3066__160/HI io_out[26] sky130_fd_sc_hd__conb_1
XFILLER_63_42 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_8_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2250_ _2454_/A _2310_/A _2385_/A vssd1 vssd1 vccd1 vccd1 _2250_/X sky130_fd_sc_hd__and3_1
X_2181_ _2181_/A _2181_/B _2380_/A vssd1 vssd1 vccd1 vccd1 _2181_/X sky130_fd_sc_hd__and3_1
XFILLER_61_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1965_ _1965_/A _1933_/B vssd1 vssd1 vccd1 vccd1 _2049_/A sky130_fd_sc_hd__or2b_1
X_1896_ _1895_/B _1895_/C _1895_/A vssd1 vssd1 vccd1 vccd1 _1901_/B sky130_fd_sc_hd__a21o_1
XFILLER_0_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2517_ _2518_/B _2518_/C _2518_/A vssd1 vssd1 vccd1 vccd1 _2600_/A sky130_fd_sc_hd__a21oi_1
X_2448_ _2446_/X _2521_/A vssd1 vssd1 vccd1 vccd1 _2449_/B sky130_fd_sc_hd__and2b_1
X_2379_ _2380_/A _2464_/A vssd1 vssd1 vccd1 vccd1 _2462_/B sky130_fd_sc_hd__nand2_1
XFILLER_44_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_408 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_78 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input36_A la_data_in[41] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_345 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_367 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1750_ _1750_/A _1750_/B vssd1 vssd1 vccd1 vccd1 _1750_/Y sky130_fd_sc_hd__xnor2_1
X_1681_ _1681_/A _1681_/B vssd1 vssd1 vccd1 vccd1 _1682_/B sky130_fd_sc_hd__and2_1
XTAP_724 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_713 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_702 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2302_ _2302_/A _2302_/B vssd1 vssd1 vccd1 vccd1 _2302_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_31_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_768 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_757 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_746 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_735 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_779 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2233_ _2305_/A _2230_/C _2233_/C _2233_/D vssd1 vssd1 vccd1 vccd1 _2296_/A sky130_fd_sc_hd__and4bb_1
X_2164_ _2110_/B _2164_/B vssd1 vssd1 vccd1 vccd1 _2164_/X sky130_fd_sc_hd__and2b_1
XANTENNA__1834__A_N _2501_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_38_356 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_38_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2095_ _2206_/B _2206_/A vssd1 vssd1 vccd1 vccd1 _2096_/A sky130_fd_sc_hd__and2b_1
XFILLER_53_359 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_0_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2997_ _2998_/A _2998_/B vssd1 vssd1 vccd1 vccd1 _2999_/A sky130_fd_sc_hd__and2_1
X_1948_ _2036_/A _2036_/B vssd1 vssd1 vccd1 vccd1 _2417_/A sky130_fd_sc_hd__nand2_1
X_1879_ input1/X _1879_/B _1975_/B vssd1 vssd1 vccd1 vccd1 _1879_/X sky130_fd_sc_hd__and3_1
XFILLER_1_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_116 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_153 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_518 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_56_186 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_56_175 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_44 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_40_510 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3178__272 vssd1 vssd1 vccd1 vccd1 _3178__272/HI wbs_dat_o[0] sky130_fd_sc_hd__conb_1
XANTENNA__2204__A1 _2568_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_40_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_466 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_304 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_164 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_35_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2920_ _2920_/A _2920_/B vssd1 vssd1 vccd1 vccd1 _2941_/A sky130_fd_sc_hd__nand2_1
XFILLER_16_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2851_ _2904_/A _2851_/B vssd1 vssd1 vccd1 vccd1 _2852_/B sky130_fd_sc_hd__or2_2
X_1802_ _1831_/A vssd1 vssd1 vccd1 vccd1 _1884_/A sky130_fd_sc_hd__clkbuf_2
X_2782_ _2808_/B _2780_/X _2732_/X _2733_/Y vssd1 vssd1 vccd1 vccd1 _2783_/C sky130_fd_sc_hd__o211a_1
X_1733_ _1733_/A _1733_/B vssd1 vssd1 vccd1 vccd1 _1756_/A sky130_fd_sc_hd__nor2_1
X_1664_ _1699_/B _1635_/B _1623_/A vssd1 vssd1 vccd1 vccd1 _1666_/A sky130_fd_sc_hd__a21o_1
X_1595_ _2933_/X _1592_/X _1593_/Y _1594_/X vssd1 vssd1 vccd1 vccd1 _1597_/B sky130_fd_sc_hd__a211o_2
XTAP_521 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_510 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_532 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_543 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_554 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_565 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_576 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2216_ _2281_/A _2216_/B vssd1 vssd1 vccd1 vccd1 _2217_/B sky130_fd_sc_hd__xnor2_1
XTAP_587 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_598 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_624 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2147_ _2177_/A _2177_/B vssd1 vssd1 vccd1 vccd1 _2178_/A sky130_fd_sc_hd__xor2_1
XFILLER_26_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2078_ _2079_/A _2138_/A vssd1 vssd1 vccd1 vccd1 _2187_/A sky130_fd_sc_hd__and2_1
XFILLER_41_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_14_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_34_381 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_30_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2956__A _2956_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_429 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3106__200 vssd1 vssd1 vccd1 vccd1 _3106__200/HI la_data_out[25] sky130_fd_sc_hd__conb_1
XFILLER_9_525 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2866__A _2939_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2001_ _2002_/A _2002_/B vssd1 vssd1 vccd1 vccd1 _2003_/A sky130_fd_sc_hd__and2_1
XFILLER_35_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2903_ _2903_/A _2903_/B vssd1 vssd1 vccd1 vccd1 _2903_/X sky130_fd_sc_hd__xor2_2
X_2834_ _2884_/A _2833_/B _2833_/C vssd1 vssd1 vccd1 vccd1 _2835_/B sky130_fd_sc_hd__a21o_1
X_2765_ _2843_/B _2764_/C _2764_/A vssd1 vssd1 vccd1 vccd1 _2768_/B sky130_fd_sc_hd__a21o_1
X_1716_ _1716_/A _1741_/A vssd1 vssd1 vccd1 vccd1 _1716_/Y sky130_fd_sc_hd__nor2_1
X_2696_ _2922_/A _2694_/X _2630_/D _2695_/Y _2538_/A vssd1 vssd1 vccd1 vccd1 _2702_/B
+ sky130_fd_sc_hd__a2111o_2
X_1647_ _1647_/A _1647_/B vssd1 vssd1 vccd1 vccd1 _1648_/B sky130_fd_sc_hd__and2_1
X_1578_ _1532_/A _1576_/Y _1577_/Y _1567_/B vssd1 vssd1 vccd1 vccd1 _1612_/A sky130_fd_sc_hd__a211o_2
XTAP_340 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_351 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1680__A _1681_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_362 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_373 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_384 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_395 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_13 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_46 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_68 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2407__A1 _1888_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XPHY_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_45 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_9_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2546__B_N _2474_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_57_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_17_145 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_17_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_424 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_40_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_6 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2550_ _2550_/A vssd1 vssd1 vccd1 vccd1 _2550_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_1501_ _2984_/A _2984_/B vssd1 vssd1 vccd1 vccd1 _1507_/B sky130_fd_sc_hd__and2b_1
XFILLER_5_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2481_ _2556_/A _2481_/B vssd1 vssd1 vccd1 vccd1 _2577_/B sky130_fd_sc_hd__xnor2_1
XFILLER_36_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_432 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3083__177 vssd1 vssd1 vccd1 vccd1 _3083__177/HI la_data_out[2] sky130_fd_sc_hd__conb_1
XFILLER_23_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_23_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2817_ _2818_/B _2818_/C _2818_/A vssd1 vssd1 vccd1 vccd1 _2825_/A sky130_fd_sc_hd__a21oi_2
X_2748_ _2748_/A vssd1 vssd1 vccd1 vccd1 _2748_/X sky130_fd_sc_hd__dlymetal6s2s_1
X_2679_ _2744_/A _2679_/B vssd1 vssd1 vccd1 vccd1 _2683_/A sky130_fd_sc_hd__xnor2_2
XFILLER_59_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_568 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XTAP_192 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_181 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_170 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2953__B _2954_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_14_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_14_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_30_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2800__A1 _2723_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_542 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_586 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_18_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_21_619 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1981_ _1981_/A _1981_/B vssd1 vssd1 vccd1 vccd1 _1982_/B sky130_fd_sc_hd__xnor2_2
XFILLER_41_490 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2602_ _2602_/A _2602_/B vssd1 vssd1 vccd1 vccd1 _2602_/X sky130_fd_sc_hd__xor2_2
X_2533_ _2534_/A _2629_/A vssd1 vssd1 vccd1 vccd1 _2694_/B sky130_fd_sc_hd__nand2_1
XFILLER_5_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2464_ _2464_/A _2464_/B vssd1 vssd1 vccd1 vccd1 _2465_/B sky130_fd_sc_hd__or2_1
X_2395_ _2454_/B vssd1 vssd1 vccd1 vccd1 _2919_/A sky130_fd_sc_hd__buf_2
X_3011__105 vssd1 vssd1 vccd1 vccd1 _3011__105/HI io_oeb[8] sky130_fd_sc_hd__conb_1
XFILLER_51_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_22_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_11 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_59_376 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_33 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_30_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2180_ _2322_/B vssd1 vssd1 vccd1 vccd1 _2380_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_18_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1964_ _2006_/A _2008_/B vssd1 vssd1 vccd1 vccd1 _1999_/A sky130_fd_sc_hd__nor2_1
XFILLER_21_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1895_ _1895_/A _1895_/B _1895_/C vssd1 vssd1 vccd1 vccd1 _1953_/A sky130_fd_sc_hd__nand3_1
X_3195__289 vssd1 vssd1 vccd1 vccd1 _3195__289/HI wbs_dat_o[17] sky130_fd_sc_hd__conb_1
X_2516_ _2509_/Y _2513_/Y _2445_/A _2450_/X vssd1 vssd1 vccd1 vccd1 _2518_/C sky130_fd_sc_hd__o211ai_2
X_2447_ _2447_/A _2447_/B vssd1 vssd1 vccd1 vccd1 _2521_/A sky130_fd_sc_hd__or2_1
XFILLER_29_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2378_ _2378_/A vssd1 vssd1 vccd1 vccd1 _2931_/A sky130_fd_sc_hd__buf_2
X_3089__183 vssd1 vssd1 vccd1 vccd1 _3089__183/HI la_data_out[8] sky130_fd_sc_hd__conb_1
XFILLER_29_538 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_58_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_58_76 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input29_A la_data_in[35] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_28_571 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_15_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_493 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1680_ _1681_/A _1681_/B vssd1 vssd1 vccd1 vccd1 _1711_/B sky130_fd_sc_hd__nor2_1
XTAP_725 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_714 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_703 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2301_ _2240_/X _2244_/B _2241_/A vssd1 vssd1 vccd1 vccd1 _2302_/B sky130_fd_sc_hd__a21o_1
XTAP_758 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_747 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_736 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_769 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2232_ _2233_/C _2233_/D _2374_/A _2231_/Y vssd1 vssd1 vccd1 vccd1 _2234_/A sky130_fd_sc_hd__a22oi_2
XFILLER_24_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2163_ _2163_/A _2163_/B vssd1 vssd1 vccd1 vccd1 _2176_/A sky130_fd_sc_hd__xor2_2
X_2094_ input2/X _2097_/B vssd1 vssd1 vccd1 vccd1 _2206_/B sky130_fd_sc_hd__xor2_1
XFILLER_19_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3123__217 vssd1 vssd1 vccd1 vccd1 _3123__217/HI la_data_out[42] sky130_fd_sc_hd__conb_1
X_2996_ _2996_/A _2996_/B vssd1 vssd1 vccd1 vccd1 _2998_/B sky130_fd_sc_hd__or2_1
XFILLER_9_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_279 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1947_ _1947_/A vssd1 vssd1 vccd1 vccd1 _2550_/A sky130_fd_sc_hd__clkbuf_2
X_1878_ _2023_/A vssd1 vssd1 vccd1 vccd1 _1975_/B sky130_fd_sc_hd__dlymetal6s2s_1
X_3017__111 vssd1 vssd1 vccd1 vccd1 _3017__111/HI io_oeb[14] sky130_fd_sc_hd__conb_1
XFILLER_0_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_56_165 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_29_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2019__A _2086_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_56 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_110 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_47_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_16_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_371 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2850_ _2850_/A _2896_/A vssd1 vssd1 vccd1 vccd1 _2851_/B sky130_fd_sc_hd__and2_1
X_1801_ _1801_/A _1830_/A vssd1 vssd1 vccd1 vccd1 _1831_/A sky130_fd_sc_hd__xor2_1
X_2781_ _2732_/X _2733_/Y _2808_/B _2780_/X vssd1 vssd1 vccd1 vccd1 _2783_/B sky130_fd_sc_hd__a211oi_2
X_1732_ _2988_/X _1731_/B _1731_/C vssd1 vssd1 vccd1 vccd1 _1733_/B sky130_fd_sc_hd__a21oi_1
X_1663_ _1663_/A vssd1 vssd1 vccd1 vccd1 _1699_/B sky130_fd_sc_hd__clkbuf_2
XFILLER_7_261 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1594_ _1515_/X _1502_/X _2966_/X _2936_/X vssd1 vssd1 vccd1 vccd1 _1594_/X sky130_fd_sc_hd__a22o_1
XTAP_500 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_522 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_511 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_533 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_544 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_555 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_566 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2215_ _2430_/A _2406_/A vssd1 vssd1 vccd1 vccd1 _2216_/B sky130_fd_sc_hd__nand2_1
XTAP_588 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_577 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_599 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2146_ _2179_/A _2146_/B vssd1 vssd1 vccd1 vccd1 _2177_/B sky130_fd_sc_hd__xor2_1
XFILLER_53_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2077_ _2130_/A _2559_/A _2073_/X _2076_/Y vssd1 vssd1 vccd1 vccd1 _2129_/A sky130_fd_sc_hd__a211o_4
XFILLER_26_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_14_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2198__A1 _2197_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2979_ _2979_/A _2979_/B vssd1 vssd1 vccd1 vccd1 _2979_/X sky130_fd_sc_hd__or2_1
XFILLER_30_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_4_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2212__A _2978_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_481 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2000_ _2000_/A _2000_/B vssd1 vssd1 vccd1 vccd1 _2002_/B sky130_fd_sc_hd__xor2_1
XFILLER_35_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2902_ _2856_/A _2856_/B _2901_/X vssd1 vssd1 vccd1 vccd1 _2903_/B sky130_fd_sc_hd__a21o_1
XFILLER_50_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2833_ _2884_/A _2833_/B _2833_/C vssd1 vssd1 vccd1 vccd1 _2884_/B sky130_fd_sc_hd__nand3_1
X_2764_ _2764_/A _2843_/B _2764_/C vssd1 vssd1 vccd1 vccd1 _2768_/A sky130_fd_sc_hd__nand3_1
X_1715_ _1741_/B _1754_/B vssd1 vssd1 vccd1 vccd1 _1718_/A sky130_fd_sc_hd__nor2_2
X_2695_ _2694_/A _2694_/C _2394_/X vssd1 vssd1 vccd1 vccd1 _2695_/Y sky130_fd_sc_hd__a21oi_2
X_1646_ _1646_/A vssd1 vssd1 vccd1 vccd1 _1716_/A sky130_fd_sc_hd__inv_2
X_1577_ _1577_/A _1577_/B vssd1 vssd1 vccd1 vccd1 _1577_/Y sky130_fd_sc_hd__nor2_1
XTAP_330 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_341 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_363 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_352 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_374 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_385 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_396 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_411 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_3129__223 vssd1 vssd1 vccd1 vccd1 _3129__223/HI la_data_out[48] sky130_fd_sc_hd__conb_1
XFILLER_27_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_54_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2129_ _2129_/A _2087_/B vssd1 vssd1 vccd1 vccd1 _2177_/A sky130_fd_sc_hd__or2b_1
XFILLER_54_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_14 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XPHY_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1615__B1 _1616_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_6_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_569 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_1_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_614 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA_input11_A la_data_in[19] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_17_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_414 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_33_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_312 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1500_ _2977_/A _2977_/B vssd1 vssd1 vccd1 vccd1 _1507_/A sky130_fd_sc_hd__and2_1
X_2480_ _2083_/X _2557_/A _2558_/A _2567_/A _2479_/X vssd1 vssd1 vccd1 vccd1 _2481_/B
+ sky130_fd_sc_hd__a221o_1
XANTENNA__2334__A1 _2400_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput90 _1575_/Y vssd1 vssd1 vccd1 vccd1 la_data_out[89] sky130_fd_sc_hd__buf_2
XFILLER_55_219 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_252 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2816_ _2814_/X _2609_/X _2815_/X vssd1 vssd1 vccd1 vccd1 _2818_/C sky130_fd_sc_hd__a21oi_2
XFILLER_11_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2747_ _2747_/A vssd1 vssd1 vccd1 vccd1 _2933_/A sky130_fd_sc_hd__clkbuf_2
X_2678_ _2739_/A _2468_/Y _2677_/Y vssd1 vssd1 vccd1 vccd1 _2679_/B sky130_fd_sc_hd__o21a_1
X_1629_ _1697_/A _1629_/B _1629_/C vssd1 vssd1 vccd1 vccd1 _1630_/B sky130_fd_sc_hd__or3_1
XFILLER_59_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input3_A la_data_in[11] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_160 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_193 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_182 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_171 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_271 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_6_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input59_A la_data_in[62] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_554 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_499 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1980_ _2377_/A _2775_/A _1978_/Y _1979_/Y vssd1 vssd1 vccd1 vccd1 _1981_/B sky130_fd_sc_hd__o211a_1
XFILLER_21_609 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1776__A input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2601_ _2521_/A _2600_/Y _2521_/B _2519_/B vssd1 vssd1 vccd1 vccd1 _2602_/B sky130_fd_sc_hd__a31o_1
XFILLER_54_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2532_ _2532_/A vssd1 vssd1 vccd1 vccd1 _2694_/A sky130_fd_sc_hd__clkbuf_2
X_2463_ _2464_/A _2534_/A vssd1 vssd1 vccd1 vccd1 _2532_/A sky130_fd_sc_hd__nand2_1
XANTENNA__2400__A _2400_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2394_ _2692_/A vssd1 vssd1 vccd1 vccd1 _2394_/X sky130_fd_sc_hd__clkbuf_2
X_3050__144 vssd1 vssd1 vccd1 vccd1 _3050__144/HI io_out[10] sky130_fd_sc_hd__conb_1
XFILLER_56_539 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_241 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_583 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_572 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_11_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_59_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_55_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_263 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_285 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1596__A _1597_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_10_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_178 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3034__128 vssd1 vssd1 vccd1 vccd1 _3034__128/HI io_oeb[31] sky130_fd_sc_hd__conb_1
XFILLER_2_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_61_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1963_ _1963_/A _1963_/B vssd1 vssd1 vccd1 vccd1 _2000_/A sky130_fd_sc_hd__nor2_1
XFILLER_33_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1894_ _1893_/B _1893_/C _1893_/A vssd1 vssd1 vccd1 vccd1 _1895_/C sky130_fd_sc_hd__a21o_1
X_2515_ _2515_/A vssd1 vssd1 vccd1 vccd1 _2518_/B sky130_fd_sc_hd__clkbuf_2
X_2446_ _2447_/A _2447_/B vssd1 vssd1 vccd1 vccd1 _2446_/X sky130_fd_sc_hd__and2_1
XFILLER_29_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2377_ _2377_/A vssd1 vssd1 vccd1 vccd1 _2538_/A sky130_fd_sc_hd__buf_2
XFILLER_17_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_37_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_564 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_36 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_163 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_28_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_520 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_55_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_15_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_30_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_11_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_443 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_715 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_704 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2300_ _2300_/A _2299_/X vssd1 vssd1 vccd1 vccd1 _2302_/A sky130_fd_sc_hd__or2b_1
XTAP_759 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_748 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_737 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_726 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2231_ _2305_/A _2230_/C _2230_/A vssd1 vssd1 vccd1 vccd1 _2231_/Y sky130_fd_sc_hd__o21ai_1
XFILLER_17_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2162_ _2226_/B _2162_/B vssd1 vssd1 vccd1 vccd1 _2163_/B sky130_fd_sc_hd__xnor2_1
X_2093_ _2205_/A _2093_/B vssd1 vssd1 vccd1 vccd1 _2105_/A sky130_fd_sc_hd__xnor2_1
XFILLER_19_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3162__256 vssd1 vssd1 vccd1 vccd1 _3162__256/HI la_data_out[113] sky130_fd_sc_hd__conb_1
XFILLER_21_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2995_ _2995_/A _2995_/B vssd1 vssd1 vccd1 vccd1 _2996_/B sky130_fd_sc_hd__and2_1
X_3203__297 vssd1 vssd1 vccd1 vccd1 _3203__297/HI wbs_dat_o[25] sky130_fd_sc_hd__conb_1
X_1946_ _1946_/A vssd1 vssd1 vccd1 vccd1 _1947_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_1877_ _2043_/A vssd1 vssd1 vccd1 vccd1 _2612_/A sky130_fd_sc_hd__clkbuf_4
X_3056__150 vssd1 vssd1 vccd1 vccd1 _3056__150/HI io_out[16] sky130_fd_sc_hd__conb_1
XFILLER_57_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2429_ _2427_/X _2429_/B vssd1 vssd1 vccd1 vccd1 _2437_/A sky130_fd_sc_hd__and2b_1
XFILLER_56_122 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_24 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1858__B input9/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_25_597 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_44_79 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_207 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_280 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input41_A la_data_in[46] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_133 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_62_158 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1800_ _1800_/A vssd1 vssd1 vccd1 vccd1 _1807_/A sky130_fd_sc_hd__clkbuf_2
X_2780_ _2808_/A _2779_/B _2779_/C vssd1 vssd1 vccd1 vccd1 _2780_/X sky130_fd_sc_hd__o21a_1
X_1731_ _2988_/X _1731_/B _1731_/C vssd1 vssd1 vccd1 vccd1 _1733_/A sky130_fd_sc_hd__and3_1
XFILLER_7_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1662_ _2965_/B _2921_/X _1761_/B _1515_/X vssd1 vssd1 vccd1 vccd1 _1666_/C sky130_fd_sc_hd__a2bb2o_1
X_3004__98 vssd1 vssd1 vccd1 vccd1 _3004__98/HI io_oeb[1] sky130_fd_sc_hd__conb_1
X_1593_ _2979_/X _2965_/B vssd1 vssd1 vccd1 vccd1 _1593_/Y sky130_fd_sc_hd__nor2_1
XTAP_501 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_523 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_512 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_534 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_545 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_556 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_567 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2214_ _2214_/A vssd1 vssd1 vccd1 vccd1 _2406_/A sky130_fd_sc_hd__dlymetal6s2s_1
XTAP_589 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_578 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_604 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2145_ _2254_/A _2145_/B vssd1 vssd1 vccd1 vccd1 _2146_/B sky130_fd_sc_hd__xnor2_1
XFILLER_38_155 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2076_ _2313_/S _2131_/A _2310_/A vssd1 vssd1 vccd1 vccd1 _2076_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_53_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_501 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_14_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2978_ _2978_/A vssd1 vssd1 vccd1 vccd1 _2983_/A sky130_fd_sc_hd__clkbuf_4
XFILLER_22_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1929_ _1929_/A _1929_/B vssd1 vssd1 vccd1 vccd1 _1929_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_39_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_39_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_29_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_57_486 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_55_23 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_615 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_44_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1588__B _1588_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1633__A1 _2684_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_4_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_412 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1498__B _2986_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2901_ _2901_/A _2901_/B vssd1 vssd1 vccd1 vccd1 _2901_/X sky130_fd_sc_hd__and2_1
XFILLER_16_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_50_128 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_353 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_191 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2832_ _2862_/A _2832_/B vssd1 vssd1 vccd1 vccd1 _2833_/C sky130_fd_sc_hd__xnor2_1
X_2763_ _2843_/A _2762_/B _2762_/C vssd1 vssd1 vccd1 vccd1 _2764_/C sky130_fd_sc_hd__a21o_1
X_1714_ _1714_/A _1714_/B vssd1 vssd1 vccd1 vccd1 _1754_/B sky130_fd_sc_hd__and2_1
X_2694_ _2694_/A _2694_/B _2694_/C vssd1 vssd1 vccd1 vccd1 _2694_/X sky130_fd_sc_hd__and3_1
X_1645_ _1647_/A _1647_/B vssd1 vssd1 vccd1 vccd1 _1646_/A sky130_fd_sc_hd__or2_1
X_1576_ _1576_/A _1649_/A vssd1 vssd1 vccd1 vccd1 _1576_/Y sky130_fd_sc_hd__nor2_1
XTAP_320 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_331 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_342 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_364 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_353 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_375 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_386 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_397 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_3168__262 vssd1 vssd1 vccd1 vccd1 _3168__262/HI la_data_out[119] sky130_fd_sc_hd__conb_1
X_2128_ _2107_/A _2163_/A _2106_/B _2090_/B _2090_/A vssd1 vssd1 vccd1 vccd1 _2226_/B
+ sky130_fd_sc_hd__o32ai_4
XFILLER_54_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XPHY_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2059_ _2059_/A _2059_/B vssd1 vssd1 vccd1 vccd1 _2059_/X sky130_fd_sc_hd__or2_1
XPHY_26 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_25_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__1615__A1 _1533_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__1615__B2 _1616_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_41_25 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_519 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_1_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_294 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_17_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_324 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2334__A2 _2333_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput80 _2522_/Y vssd1 vssd1 vccd1 vccd1 la_data_out[79] sky130_fd_sc_hd__buf_2
Xoutput91 _1620_/Y vssd1 vssd1 vccd1 vccd1 la_data_out[90] sky130_fd_sc_hd__buf_2
XFILLER_0_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_456 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_31_194 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2815_ _2697_/A _2549_/X _2550_/X _2394_/X vssd1 vssd1 vccd1 vccd1 _2815_/X sky130_fd_sc_hd__a22o_1
X_2746_ _2824_/A vssd1 vssd1 vccd1 vccd1 _2976_/A sky130_fd_sc_hd__buf_4
XANTENNA__1972__A _1972_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2677_ _2747_/A _2609_/X _2676_/X vssd1 vssd1 vccd1 vccd1 _2677_/Y sky130_fd_sc_hd__a21oi_1
X_1628_ _1697_/A _1629_/B _1629_/C vssd1 vssd1 vccd1 vccd1 _1681_/A sky130_fd_sc_hd__o21ai_4
XANTENNA__1691__B _1723_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1559_ _1558_/B _1559_/B vssd1 vssd1 vccd1 vccd1 _1560_/B sky130_fd_sc_hd__and2b_1
XTAP_150 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_183 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_172 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_161 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_194 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_35 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2978__A _2978_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_2_566 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_242 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_161 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2600_ _2600_/A vssd1 vssd1 vccd1 vccd1 _2600_/Y sky130_fd_sc_hd__inv_2
X_2531_ _2130_/X _2697_/A _2766_/A vssd1 vssd1 vccd1 vccd1 _2544_/A sky130_fd_sc_hd__a21oi_4
X_2462_ _2462_/A _2462_/B _2462_/C vssd1 vssd1 vccd1 vccd1 _2467_/B sky130_fd_sc_hd__and3_1
XFILLER_47_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2400__B _2528_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2393_ _2393_/A _2454_/B _2692_/A vssd1 vssd1 vccd1 vccd1 _2393_/X sky130_fd_sc_hd__and3_1
XFILLER_56_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_56_507 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_28_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_36_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_51_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_51_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_610 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2729_ _2729_/A _2729_/B vssd1 vssd1 vccd1 vccd1 _2730_/A sky130_fd_sc_hd__and2_1
XFILLER_59_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_47_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_27_220 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_42_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_278 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1596__B _1597_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_8_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3073__167 vssd1 vssd1 vccd1 vccd1 _3073__167/HI io_out[33] sky130_fd_sc_hd__conb_1
XANTENNA__2501__A _2501_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_2_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_264 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_18_275 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_33_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1962_ _1962_/A _1962_/B vssd1 vssd1 vccd1 vccd1 _1962_/Y sky130_fd_sc_hd__xnor2_1
X_1893_ _1893_/A _1893_/B _1893_/C vssd1 vssd1 vccd1 vccd1 _1895_/B sky130_fd_sc_hd__nand3_1
X_2514_ _2445_/A _2450_/X _2509_/Y _2513_/Y vssd1 vssd1 vccd1 vccd1 _2515_/A sky130_fd_sc_hd__a211o_1
X_2445_ _2445_/A _2445_/B vssd1 vssd1 vccd1 vccd1 _2447_/B sky130_fd_sc_hd__and2_1
X_2376_ _2354_/B _2354_/C _2354_/A vssd1 vssd1 vccd1 vccd1 _2427_/A sky130_fd_sc_hd__a21bo_1
XFILLER_56_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_3208__302 vssd1 vssd1 vccd1 vccd1 _3208__302/HI wbs_dat_o[30] sky130_fd_sc_hd__conb_1
XFILLER_37_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_576 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_407 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_598 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_48 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_473 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_47_315 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_62_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_15_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_716 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_705 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_749 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_738 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_727 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2230_ _2230_/A _2305_/A _2230_/C vssd1 vssd1 vccd1 vccd1 _2374_/A sky130_fd_sc_hd__or3_2
X_2161_ _2178_/A _2178_/B vssd1 vssd1 vccd1 vccd1 _2162_/B sky130_fd_sc_hd__xnor2_1
XFILLER_38_326 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2092_ _1929_/Y _2037_/A _1988_/A _2404_/A _2091_/X vssd1 vssd1 vccd1 vccd1 _2093_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_0_74 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_595 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_61_395 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2994_ _2995_/A _2995_/B vssd1 vssd1 vccd1 vccd1 _2996_/A sky130_fd_sc_hd__nor2_1
XFILLER_21_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_34_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1945_ _2036_/A _1985_/B vssd1 vssd1 vccd1 vccd1 _1946_/A sky130_fd_sc_hd__nor2_1
X_1876_ _1876_/A _1876_/B vssd1 vssd1 vccd1 vccd1 _1908_/A sky130_fd_sc_hd__nor2_1
XFILLER_0_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2428_ _2427_/B _2427_/C _2427_/A vssd1 vssd1 vccd1 vccd1 _2429_/B sky130_fd_sc_hd__a21o_1
XFILLER_57_613 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2359_ _2438_/A _2357_/X _2272_/A _2284_/B vssd1 vssd1 vccd1 vccd1 _2360_/B sky130_fd_sc_hd__o211a_1
XFILLER_28_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_29_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_56_134 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_59 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_25_543 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_351 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2986__A _2986_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input34_A la_data_in[3] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3185__279 vssd1 vssd1 vccd1 vccd1 _3185__279/HI wbs_dat_o[7] sky130_fd_sc_hd__conb_1
XFILLER_35_329 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_81 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1730_ _1730_/A _1730_/B vssd1 vssd1 vccd1 vccd1 _1731_/C sky130_fd_sc_hd__xor2_1
XFILLER_11_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1661_ _1550_/X _1502_/X _1592_/X _1514_/X vssd1 vssd1 vccd1 vccd1 _1666_/B sky130_fd_sc_hd__a22o_1
X_3079__173 vssd1 vssd1 vccd1 vccd1 _3079__173/HI irq[1] sky130_fd_sc_hd__conb_1
X_1592_ _2772_/X vssd1 vssd1 vccd1 vccd1 _1592_/X sky130_fd_sc_hd__clkbuf_2
XTAP_502 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_524 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_513 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_535 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_546 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_557 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2213_ input2/X input3/X vssd1 vssd1 vccd1 vccd1 _2214_/A sky130_fd_sc_hd__xor2_1
XTAP_568 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_579 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2144_ _2410_/A _2194_/A _2141_/Y _2027_/X _2143_/X vssd1 vssd1 vccd1 vccd1 _2145_/B
+ sky130_fd_sc_hd__a221o_2
XFILLER_54_616 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_26_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_53_115 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2075_ _2181_/B vssd1 vssd1 vccd1 vccd1 _2310_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_61_181 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2977_ _2977_/A _2977_/B vssd1 vssd1 vccd1 vccd1 _2984_/A sky130_fd_sc_hd__xnor2_4
X_1928_ _1928_/A _1928_/B vssd1 vssd1 vccd1 vccd1 _1929_/B sky130_fd_sc_hd__nor2_2
X_1859_ _1924_/A _1859_/B vssd1 vssd1 vccd1 vccd1 _1859_/Y sky130_fd_sc_hd__xnor2_4
XFILLER_1_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_39_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_605 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_44_148 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_13_502 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XANTENNA__1633__A2 _2871_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_9_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_4_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3113__207 vssd1 vssd1 vccd1 vccd1 _3113__207/HI la_data_out[32] sky130_fd_sc_hd__conb_1
XFILLER_20_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_0_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_410 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_48_421 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_104 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_35_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3007__101 vssd1 vssd1 vccd1 vccd1 _3007__101/HI io_oeb[4] sky130_fd_sc_hd__conb_1
X_2900_ _2956_/A _2958_/B vssd1 vssd1 vccd1 vccd1 _2903_/A sky130_fd_sc_hd__xnor2_2
XFILLER_31_343 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2831_ _2758_/X _2930_/A _2828_/Y _2830_/X vssd1 vssd1 vccd1 vccd1 _2832_/B sky130_fd_sc_hd__a211o_1
X_2762_ _2843_/A _2762_/B _2762_/C vssd1 vssd1 vccd1 vccd1 _2843_/B sky130_fd_sc_hd__nand3_1
X_1713_ _1714_/A _1714_/B vssd1 vssd1 vccd1 vccd1 _1741_/B sky130_fd_sc_hd__nor2_1
XFILLER_8_594 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2693_ _2467_/A _2467_/B _2467_/C _2536_/C vssd1 vssd1 vccd1 vccd1 _2694_/C sky130_fd_sc_hd__a211o_1
X_1644_ _1688_/A _1644_/B vssd1 vssd1 vccd1 vccd1 _1647_/B sky130_fd_sc_hd__nor2_1
X_1575_ _1614_/B _1575_/B vssd1 vssd1 vccd1 vccd1 _1575_/Y sky130_fd_sc_hd__xnor2_1
XTAP_310 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_321 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_332 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_343 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_365 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_354 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_376 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_387 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_398 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_402 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
X_2127_ _2127_/A _2235_/A vssd1 vssd1 vccd1 vccd1 _2233_/C sky130_fd_sc_hd__nor2_1
XPHY_16 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2058_ _2059_/A _2059_/B vssd1 vssd1 vccd1 vccd1 _2060_/A sky130_fd_sc_hd__and2_1
XPHY_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_41_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1615__A2 _1533_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_22_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_41_37 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_1_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_273 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_60_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_13_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
Xoutput70 _1915_/Y vssd1 vssd1 vccd1 vccd1 la_data_out[69] sky130_fd_sc_hd__buf_2
Xoutput81 _2602_/X vssd1 vssd1 vccd1 vccd1 la_data_out[80] sky130_fd_sc_hd__buf_2
Xoutput92 _1654_/Y vssd1 vssd1 vccd1 vccd1 la_data_out[91] sky130_fd_sc_hd__buf_2
XFILLER_48_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_51_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2814_ _2814_/A vssd1 vssd1 vccd1 vccd1 _2814_/X sky130_fd_sc_hd__clkbuf_2
X_2745_ _2972_/A _2745_/B _2745_/C vssd1 vssd1 vccd1 vccd1 _2755_/C sky130_fd_sc_hd__nand3_1
X_2676_ _2391_/A _2549_/X _2550_/A _2385_/A vssd1 vssd1 vccd1 vccd1 _2676_/X sky130_fd_sc_hd__a22o_1
X_1627_ _1515_/X _1592_/X _1624_/Y _1626_/X vssd1 vssd1 vccd1 vccd1 _1629_/C sky130_fd_sc_hd__a211o_1
XANTENNA__1972__B _1974_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1558_ _1559_/B _1558_/B vssd1 vssd1 vccd1 vccd1 _1560_/A sky130_fd_sc_hd__and2b_1
XFILLER_59_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XTAP_140 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1489_ _2960_/A _2960_/B _2955_/A vssd1 vssd1 vccd1 vccd1 _1490_/B sky130_fd_sc_hd__a21o_1
XTAP_184 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_173 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_162 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_151 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_195 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_15_608 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_54_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_14_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_58 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_379 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_2_578 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_18_435 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_45_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_33_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3119__213 vssd1 vssd1 vccd1 vccd1 _3119__213/HI la_data_out[38] sky130_fd_sc_hd__conb_1
X_2530_ _2530_/A vssd1 vssd1 vccd1 vccd1 _2766_/A sky130_fd_sc_hd__clkbuf_4
X_2461_ _2461_/A _2461_/B vssd1 vssd1 vccd1 vccd1 _2462_/C sky130_fd_sc_hd__nand2_1
XANTENNA__2400__C _2400_/C vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2392_ _2629_/A vssd1 vssd1 vccd1 vccd1 _2692_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_3_63 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_96 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2409__A _2978_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_64_596 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_24_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_24_438 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_298 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_51_257 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_600 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_622 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2728_ _2728_/A _2728_/B vssd1 vssd1 vccd1 vccd1 _2729_/B sky130_fd_sc_hd__or2_1
X_2659_ _2589_/B _2589_/Y _2657_/Y _2658_/X vssd1 vssd1 vccd1 vccd1 _2718_/A sky130_fd_sc_hd__o211ai_1
XFILLER_59_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_15_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_6_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input64_A la_data_in[9] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_397 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_46_552 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_563 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_287 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1961_ _1911_/X _1915_/B _1912_/A vssd1 vssd1 vccd1 vccd1 _1962_/B sky130_fd_sc_hd__a21o_1
X_1892_ _1981_/A _1892_/B _1892_/C _1892_/D vssd1 vssd1 vccd1 vccd1 _1893_/C sky130_fd_sc_hd__or4_1
X_2513_ _2595_/A _2512_/Y _2523_/A vssd1 vssd1 vccd1 vccd1 _2513_/Y sky130_fd_sc_hd__a21boi_1
X_2444_ _2444_/A _2444_/B _2444_/C _2444_/D vssd1 vssd1 vccd1 vccd1 _2445_/B sky130_fd_sc_hd__nand4_1
X_2375_ _2296_/A _2296_/B _2306_/Y _2364_/X _2374_/Y vssd1 vssd1 vccd1 vccd1 _2444_/C
+ sky130_fd_sc_hd__o221ai_2
XFILLER_56_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_419 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_607 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_57 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_47_305 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_55_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_43_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3040__134 vssd1 vssd1 vccd1 vccd1 _3040__134/HI io_oeb[37] sky130_fd_sc_hd__conb_1
XFILLER_7_401 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_11_485 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_23_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_706 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_739 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_728 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_717 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2160_ _2160_/A _2160_/B vssd1 vssd1 vccd1 vccd1 _2178_/B sky130_fd_sc_hd__and2_1
XFILLER_0_20 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2091_ _2021_/A _1943_/A _1947_/A _2034_/A vssd1 vssd1 vccd1 vccd1 _2091_/X sky130_fd_sc_hd__a22o_1
XFILLER_38_338 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_574 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_46_360 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_19_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2993_ _2944_/A _2944_/B _2943_/B _2943_/A vssd1 vssd1 vccd1 vccd1 _2995_/B sky130_fd_sc_hd__o2bb2a_1
XFILLER_21_216 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1944_ _1944_/A _1944_/B vssd1 vssd1 vccd1 vccd1 _1985_/B sky130_fd_sc_hd__xnor2_1
XFILLER_21_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1875_ _1875_/A _1913_/B vssd1 vssd1 vccd1 vccd1 _1875_/Y sky130_fd_sc_hd__xnor2_1
XANTENNA__2422__A _2818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2427_ _2427_/A _2427_/B _2427_/C vssd1 vssd1 vccd1 vccd1 _2427_/X sky130_fd_sc_hd__and3_1
XFILLER_56_102 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2358_ _2272_/A _2284_/B _2438_/A _2357_/X vssd1 vssd1 vccd1 vccd1 _2438_/B sky130_fd_sc_hd__a211oi_1
XFILLER_28_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2289_ _2289_/A _2289_/B vssd1 vssd1 vccd1 vccd1 _2307_/B sky130_fd_sc_hd__and2_1
XFILLER_29_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3024__118 vssd1 vssd1 vccd1 vccd1 _3024__118/HI io_oeb[21] sky130_fd_sc_hd__conb_1
XFILLER_52_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_12_238 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_4_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input27_A la_data_in[33] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_47_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_308 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_319 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_43_330 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_31_503 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1660_ _1611_/A _1647_/B _1659_/Y _1612_/A _1648_/B vssd1 vssd1 vccd1 vccd1 _1690_/A
+ sky130_fd_sc_hd__a221o_2
X_1591_ _2977_/A _1548_/B _1590_/X vssd1 vssd1 vccd1 vccd1 _1597_/A sky130_fd_sc_hd__a21o_2
XFILLER_7_297 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_470 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_503 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_525 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_514 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_536 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_547 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_558 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2212_ _2978_/A vssd1 vssd1 vccd1 vccd1 _2281_/A sky130_fd_sc_hd__inv_2
XTAP_569 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_603 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2143_ _2071_/A _2316_/A _2386_/A _1968_/C vssd1 vssd1 vccd1 vccd1 _2143_/X sky130_fd_sc_hd__a22o_1
XFILLER_53_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_19_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2074_ _2255_/A vssd1 vssd1 vccd1 vccd1 _2131_/A sky130_fd_sc_hd__dlymetal6s2s_1
XFILLER_61_193 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2976_ _2976_/A _2976_/B vssd1 vssd1 vccd1 vccd1 _2977_/B sky130_fd_sc_hd__xnor2_2
X_1927_ _1972_/A _1974_/A vssd1 vssd1 vccd1 vccd1 _1928_/B sky130_fd_sc_hd__and2_1
X_1858_ input8/X input9/X vssd1 vssd1 vccd1 vccd1 _1859_/B sky130_fd_sc_hd__and2b_1
X_1789_ _1813_/B _1789_/B vssd1 vssd1 vccd1 vccd1 _1789_/Y sky130_fd_sc_hd__nor2_1
XFILLER_39_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_57_444 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_29_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_47 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_44_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_322 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_4_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_3152__246 vssd1 vssd1 vccd1 vccd1 _3152__246/HI la_data_out[103] sky130_fd_sc_hd__conb_1
XFILLER_20_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_48_433 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_48_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_35_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3046__140 vssd1 vssd1 vccd1 vccd1 _3046__140/HI io_out[6] sky130_fd_sc_hd__conb_1
XFILLER_16_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_385 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_45_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2830_ _2863_/A _2934_/A _2935_/A _2913_/A vssd1 vssd1 vccd1 vccd1 _2830_/X sky130_fd_sc_hd__a22o_1
XFILLER_31_388 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2761_ _2862_/A _2761_/B vssd1 vssd1 vccd1 vccd1 _2762_/C sky130_fd_sc_hd__xnor2_1
X_1712_ _1753_/A _1712_/B vssd1 vssd1 vccd1 vccd1 _1714_/B sky130_fd_sc_hd__and2_1
XFILLER_8_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2692_ _2692_/A vssd1 vssd1 vccd1 vccd1 _2922_/A sky130_fd_sc_hd__buf_2
X_1643_ _1643_/A _1643_/B _1643_/C vssd1 vssd1 vccd1 vccd1 _1644_/B sky130_fd_sc_hd__nor3_1
XFILLER_8_584 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1574_ _1533_/A _1533_/B _1573_/X vssd1 vssd1 vccd1 vccd1 _1575_/B sky130_fd_sc_hd__a21o_1
XTAP_300 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_311 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_322 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_333 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_344 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_366 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_355 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_377 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_388 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_399 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_27_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_27_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2126_ _2118_/A _2124_/Y _2125_/Y vssd1 vssd1 vccd1 vccd1 _2170_/A sky130_fd_sc_hd__a21oi_2
XFILLER_26_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_17 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2057_ _2057_/A _2057_/B vssd1 vssd1 vccd1 vccd1 _2059_/B sky130_fd_sc_hd__xnor2_1
XPHY_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XPHY_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_34_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2959_ _2856_/A _2856_/B _2903_/A _2957_/X _2958_/Y vssd1 vssd1 vccd1 vccd1 _2960_/B
+ sky130_fd_sc_hd__a32o_1
XFILLER_1_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_17_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_41_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput93 _1692_/Y vssd1 vssd1 vccd1 vccd1 la_data_out[92] sky130_fd_sc_hd__buf_2
Xoutput71 _1962_/Y vssd1 vssd1 vccd1 vccd1 la_data_out[70] sky130_fd_sc_hd__buf_2
Xoutput82 _2668_/Y vssd1 vssd1 vccd1 vccd1 la_data_out[81] sky130_fd_sc_hd__buf_2
XFILLER_63_288 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2813_ _2973_/A _2973_/B _2739_/A vssd1 vssd1 vccd1 vccd1 _2818_/B sky130_fd_sc_hd__a21o_1
X_2744_ _2744_/A vssd1 vssd1 vccd1 vccd1 _2972_/A sky130_fd_sc_hd__buf_2
X_2675_ _2712_/B _2640_/B _2640_/C _2674_/X vssd1 vssd1 vccd1 vccd1 _2732_/A sky130_fd_sc_hd__o31a_1
X_1626_ _1514_/X _1502_/X _1761_/B _2933_/X vssd1 vssd1 vccd1 vccd1 _1626_/X sky130_fd_sc_hd__a22o_1
X_1557_ _1557_/A _1557_/B vssd1 vssd1 vccd1 vccd1 _1558_/B sky130_fd_sc_hd__xor2_2
XFILLER_59_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_130 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_141 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1488_ _1488_/A _1488_/B vssd1 vssd1 vccd1 vccd1 _1490_/A sky130_fd_sc_hd__xor2_2
XTAP_174 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_152 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_163 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_196 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_185 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_54_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_27_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_36_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2109_ _2048_/A _2048_/B _2108_/Y vssd1 vssd1 vccd1 vccd1 _2110_/B sky130_fd_sc_hd__a21oi_1
XFILLER_27_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_36_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_54_277 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_303 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_10_336 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_58_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_233 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_26_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_33_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_60_247 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_26_491 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_258 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_185 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_41_461 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3158__252 vssd1 vssd1 vccd1 vccd1 _3158__252/HI la_data_out[109] sky130_fd_sc_hd__conb_1
X_2460_ _2192_/B _2192_/C _2258_/A _2459_/Y _2192_/A vssd1 vssd1 vccd1 vccd1 _2467_/A
+ sky130_fd_sc_hd__a2111o_1
X_2391_ _2391_/A vssd1 vssd1 vccd1 vccd1 _2814_/A sky130_fd_sc_hd__buf_2
XFILLER_51_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2727_ _2728_/A _2728_/B vssd1 vssd1 vccd1 vccd1 _2729_/A sky130_fd_sc_hd__nand2_1
X_2658_ _2657_/B _2657_/C _2657_/A vssd1 vssd1 vccd1 vccd1 _2658_/X sky130_fd_sc_hd__a21o_1
X_1609_ _1610_/A _1610_/B vssd1 vssd1 vccd1 vccd1 _1611_/A sky130_fd_sc_hd__and2_1
X_2589_ _2589_/A _2589_/B _2589_/C vssd1 vssd1 vccd1 vccd1 _2589_/Y sky130_fd_sc_hd__nor3_2
XANTENNA_input1_A la_data_in[0] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_55_553 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_15_428 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_42_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_63_69 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_166 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_6_137 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_12_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_95 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_2_332 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input57_A la_data_in[60] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_58_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_33_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_299 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_21_409 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1960_ _1960_/A _1959_/X vssd1 vssd1 vccd1 vccd1 _1962_/A sky130_fd_sc_hd__or2b_1
X_1891_ _1892_/B _1892_/C _1892_/D _2329_/A vssd1 vssd1 vccd1 vccd1 _1893_/B sky130_fd_sc_hd__o31ai_2
XFILLER_52_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2512_ _2512_/A _2523_/B vssd1 vssd1 vccd1 vccd1 _2512_/Y sky130_fd_sc_hd__nand2_1
X_2443_ _2444_/A _2444_/B _2444_/C _2444_/D vssd1 vssd1 vccd1 vccd1 _2445_/A sky130_fd_sc_hd__a31o_1
X_2374_ _2374_/A _2374_/B vssd1 vssd1 vccd1 vccd1 _2374_/Y sky130_fd_sc_hd__nand2_1
XFILLER_56_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_52_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_203 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_28 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_59_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_55_383 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__1888__B _1888_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_15_225 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_11_442 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_413 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_23_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__2915__A1 _2141_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_707 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_729 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_718 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_2_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_38_317 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2090_ _2090_/A _2090_/B vssd1 vssd1 vccd1 vccd1 _2107_/A sky130_fd_sc_hd__xnor2_2
XFILLER_0_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_54 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_34_545 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_567 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2992_ _2992_/A _2992_/B vssd1 vssd1 vccd1 vccd1 _2995_/A sky130_fd_sc_hd__xnor2_1
XFILLER_34_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1943_ _1943_/A vssd1 vssd1 vccd1 vccd1 _2549_/A sky130_fd_sc_hd__clkbuf_2
XANTENNA__2703__A _2703_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1874_ _1843_/A _1843_/B _1844_/X vssd1 vssd1 vccd1 vccd1 _1913_/B sky130_fd_sc_hd__a21o_1
XANTENNA__2382__A2 _2931_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2426_ _2425_/A _2425_/B _2425_/C vssd1 vssd1 vccd1 vccd1 _2427_/C sky130_fd_sc_hd__a21o_1
X_2357_ _2354_/X _2355_/Y _2308_/X _2309_/X vssd1 vssd1 vccd1 vccd1 _2357_/X sky130_fd_sc_hd__o211a_1
XFILLER_29_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_114 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2288_ _2288_/A _2288_/B vssd1 vssd1 vccd1 vccd1 _2307_/A sky130_fd_sc_hd__xnor2_1
XFILLER_44_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_523 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_372 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_556 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_38 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3063__157 vssd1 vssd1 vccd1 vccd1 _3063__157/HI io_out[23] sky130_fd_sc_hd__conb_1
XFILLER_52_386 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_12_217 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_60_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3104__198 vssd1 vssd1 vccd1 vccd1 _3104__198/HI la_data_out[23] sky130_fd_sc_hd__conb_1
XFILLER_47_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_62_106 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_28_394 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_589 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_31_559 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_265 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_254 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_1590_ _1554_/A _1590_/B vssd1 vssd1 vccd1 vccd1 _1590_/X sky130_fd_sc_hd__and2b_1
XFILLER_7_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_515 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_504 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_526 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_537 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_548 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2211_ input5/X vssd1 vssd1 vccd1 vccd1 _2978_/A sky130_fd_sc_hd__clkbuf_4
XTAP_559 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2142_ _2142_/A vssd1 vssd1 vccd1 vccd1 _2386_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_38_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_38_136 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2073_ _2181_/A _2134_/B _2255_/A vssd1 vssd1 vccd1 vccd1 _2073_/X sky130_fd_sc_hd__and3_1
XFILLER_26_309 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_38_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_19_361 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2975_ _2814_/X _2820_/X _2973_/Y _2557_/X _2974_/X vssd1 vssd1 vccd1 vccd1 _2976_/B
+ sky130_fd_sc_hd__a221o_1
X_1926_ _1926_/A _1975_/A vssd1 vssd1 vccd1 vccd1 _1928_/A sky130_fd_sc_hd__nor2_1
XFILLER_30_570 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1857_ _1884_/A _1884_/B vssd1 vssd1 vccd1 vccd1 _2377_/A sky130_fd_sc_hd__nand2_2
X_1788_ _1788_/A _1788_/B vssd1 vssd1 vccd1 vccd1 _1789_/B sky130_fd_sc_hd__nor2_1
X_2409_ _2978_/A _2409_/B vssd1 vssd1 vccd1 vccd1 _2493_/A sky130_fd_sc_hd__xnor2_2
XFILLER_55_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1512__A _2818_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2608__A _2608_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_180 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_515 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_537 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_334 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_378 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3191__285 vssd1 vssd1 vccd1 vccd1 _3191__285/HI wbs_dat_o[13] sky130_fd_sc_hd__conb_1
XFILLER_0_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_48_445 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_63_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_29_82 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2518__A _2518_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_48_489 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_581 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2760_ _2141_/Y _2684_/X _2930_/A _2686_/X _2759_/X vssd1 vssd1 vccd1 vccd1 _2761_/B
+ sky130_fd_sc_hd__a221o_1
XFILLER_61_91 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1711_ _1711_/A _1711_/B _1711_/C vssd1 vssd1 vccd1 vccd1 _1712_/B sky130_fd_sc_hd__or3_1
X_2691_ _2637_/A _2637_/B _2766_/A vssd1 vssd1 vccd1 vccd1 _2704_/A sky130_fd_sc_hd__a21o_1
X_1642_ _1643_/A _1643_/B _1643_/C vssd1 vssd1 vccd1 vccd1 _1688_/A sky130_fd_sc_hd__o21a_1
XFILLER_6_31 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1573_ _1614_/A _1573_/B vssd1 vssd1 vccd1 vccd1 _1573_/X sky130_fd_sc_hd__and2b_1
XTAP_301 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_312 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_323 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_58_209 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XTAP_334 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_345 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_367 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_356 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_378 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_389 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2125_ _2125_/A _2125_/B vssd1 vssd1 vccd1 vccd1 _2125_/Y sky130_fd_sc_hd__nor2_1
XFILLER_26_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2056_ _2064_/A _2064_/B vssd1 vssd1 vccd1 vccd1 _2057_/B sky130_fd_sc_hd__xnor2_1
XPHY_18 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XPHY_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_26_139 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_22_301 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_50_621 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1986__B _2927_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2958_ _2958_/A _2958_/B vssd1 vssd1 vccd1 vccd1 _2958_/Y sky130_fd_sc_hd__nand2_1
XFILLER_22_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1909_ _2006_/A _1908_/C _1908_/A vssd1 vssd1 vccd1 vccd1 _1910_/C sky130_fd_sc_hd__a21o_1
X_2889_ _2846_/A _2846_/B _2847_/B _2847_/A vssd1 vssd1 vccd1 vccd1 _2908_/B sky130_fd_sc_hd__a22oi_2
X_3175__269 vssd1 vssd1 vccd1 vccd1 _3175__269/HI la_data_out[126] sky130_fd_sc_hd__conb_1
XFILLER_57_231 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3069__163 vssd1 vssd1 vccd1 vccd1 _3069__163/HI io_out[29] sky130_fd_sc_hd__conb_1
XFILLER_25_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_15_51 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_131 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_40_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_500 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_72 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_5_588 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_5_577 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
Xoutput72 _2005_/Y vssd1 vssd1 vccd1 vccd1 la_data_out[71] sky130_fd_sc_hd__buf_2
Xoutput83 _2730_/X vssd1 vssd1 vccd1 vccd1 la_data_out[82] sky130_fd_sc_hd__buf_2
Xoutput94 _1725_/Y vssd1 vssd1 vccd1 vccd1 la_data_out[93] sky130_fd_sc_hd__buf_2
XFILLER_48_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2248__A _2380_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_36_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_415 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_63_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_172 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2812_ _2877_/A _2812_/B vssd1 vssd1 vccd1 vccd1 _2836_/A sky130_fd_sc_hd__nor2_1
X_2743_ _2745_/B _2745_/C _2744_/A vssd1 vssd1 vccd1 vccd1 _2755_/B sky130_fd_sc_hd__a21o_1
X_2674_ _2674_/A _2548_/B vssd1 vssd1 vccd1 vccd1 _2674_/X sky130_fd_sc_hd__or2b_1
X_1625_ _2966_/X vssd1 vssd1 vccd1 vccd1 _1761_/B sky130_fd_sc_hd__clkbuf_2
X_1556_ _1588_/B _1556_/B vssd1 vssd1 vccd1 vccd1 _1557_/B sky130_fd_sc_hd__xor2_4
XFILLER_59_529 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_131 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_175 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_153 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_142 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_164 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1487_ _2999_/X _1487_/B vssd1 vssd1 vccd1 vccd1 _1488_/B sky130_fd_sc_hd__xnor2_4
XTAP_197 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_186 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_253 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2108_ _2108_/A _2108_/B vssd1 vssd1 vccd1 vccd1 _2108_/Y sky130_fd_sc_hd__nor2_1
XFILLER_27_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_27_459 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_54_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2039_ _2039_/A _2039_/B vssd1 vssd1 vccd1 vccd1 _2040_/B sky130_fd_sc_hd__nor2_1
XFILLER_52_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_50_451 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_50_462 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_348 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_58_573 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_404 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2485__A1 _1929_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_45_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_113 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_13_197 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3197__291 vssd1 vssd1 vccd1 vccd1 _3197__291/HI wbs_dat_o[19] sky130_fd_sc_hd__conb_1
XFILLER_42_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_5_374 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_5_341 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_5_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2390_ _2700_/A _2390_/B _2390_/C vssd1 vssd1 vccd1 vccd1 _2399_/C sky130_fd_sc_hd__nand3_1
XFILLER_3_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_3_32 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_201 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_36_223 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_64_587 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_36_245 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_51_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2726_ _2602_/A _2602_/B _2668_/A _2724_/X _2725_/X vssd1 vssd1 vccd1 vccd1 _2728_/B
+ sky130_fd_sc_hd__a32o_1
X_2657_ _2657_/A _2657_/B _2657_/C vssd1 vssd1 vccd1 vccd1 _2657_/Y sky130_fd_sc_hd__nand3_1
X_1608_ _1621_/B _1608_/B vssd1 vssd1 vccd1 vccd1 _1610_/B sky130_fd_sc_hd__xnor2_1
X_2588_ _2585_/X _2586_/Y _2526_/X _2527_/Y vssd1 vssd1 vccd1 vccd1 _2589_/C sky130_fd_sc_hd__o211a_1
XFILLER_59_337 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_1539_ _1539_/A _1539_/B vssd1 vssd1 vccd1 vccd1 _1544_/B sky130_fd_sc_hd__and2_1
XANTENNA__1520__A _1555_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_42_237 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_10_101 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_123 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_7_606 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_6_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_12_41 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_12_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_2_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XANTENNA__1989__A1_N _1859_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_37_60 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_256 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_513 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_61_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_33_259 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_1890_ _1890_/A _2022_/A vssd1 vssd1 vccd1 vccd1 _1892_/D sky130_fd_sc_hd__and2_1
XFILLER_41_270 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2511_ _2512_/A _2523_/B vssd1 vssd1 vccd1 vccd1 _2595_/A sky130_fd_sc_hd__or2_1
X_2442_ _2451_/B _2442_/B vssd1 vssd1 vccd1 vccd1 _2444_/D sky130_fd_sc_hd__xor2_1
XFILLER_45_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2373_ _2306_/Y _2364_/X _2294_/B vssd1 vssd1 vccd1 vccd1 _2444_/B sky130_fd_sc_hd__o21ai_1
XANTENNA__1605__A _1605_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_56_307 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_521 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_37_532 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_24_215 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2436__A _2525_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_24_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2621__B2 _2567_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_20_465 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2709_ _1929_/Y _2880_/A _2578_/A _2402_/X vssd1 vssd1 vccd1 vccd1 _2710_/B sky130_fd_sc_hd__a22o_1
XFILLER_58_15 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XANTENNA__2688__A1 _2083_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_167 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_59_189 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_3109__203 vssd1 vssd1 vccd1 vccd1 _3109__203/HI la_data_out[28] sky130_fd_sc_hd__conb_1
XFILLER_23_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_447 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_425 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_469 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XTAP_719 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_708 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_70 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_48_92 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_61_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_88 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2991_ _2991_/A _2991_/B vssd1 vssd1 vccd1 vccd1 _2992_/B sky130_fd_sc_hd__xor2_1
XFILLER_34_579 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1942_ _1942_/A vssd1 vssd1 vccd1 vccd1 _1943_/A sky130_fd_sc_hd__dlymetal6s2s_1
X_1873_ _1873_/A _1873_/B vssd1 vssd1 vccd1 vccd1 _1875_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__2703__B _2703_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2425_ _2425_/A _2425_/B _2425_/C vssd1 vssd1 vccd1 vccd1 _2427_/B sky130_fd_sc_hd__nand3_1
XFILLER_29_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2356_ _2308_/X _2309_/X _2354_/X _2355_/Y vssd1 vssd1 vccd1 vccd1 _2438_/A sky130_fd_sc_hd__a211oi_2
XFILLER_56_126 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_2287_ _2210_/A _2210_/B _2219_/B vssd1 vssd1 vccd1 vccd1 _2288_/B sky130_fd_sc_hd__a21oi_2
XFILLER_37_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_398 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_12_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_60_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_20_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_49 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_18_73 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_16_546 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_11_240 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_7_222 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_7_211 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_516 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_505 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_59_80 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2210_ _2210_/A _2210_/B vssd1 vssd1 vccd1 vccd1 _2218_/B sky130_fd_sc_hd__xor2_1
XTAP_527 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_538 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_549 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2141_ _2187_/C _2141_/B vssd1 vssd1 vccd1 vccd1 _2141_/Y sky130_fd_sc_hd__xnor2_4
X_2072_ _2188_/B vssd1 vssd1 vccd1 vccd1 _2255_/A sky130_fd_sc_hd__buf_2
XFILLER_53_107 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_46_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_34_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2974_ _2810_/A _2748_/X _2749_/X _2922_/X vssd1 vssd1 vccd1 vccd1 _2974_/X sky130_fd_sc_hd__a22o_1
X_1925_ _1923_/X _1887_/B _1924_/X vssd1 vssd1 vccd1 vccd1 _1929_/A sky130_fd_sc_hd__a21oi_2
XFILLER_30_582 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
X_1856_ _1856_/A vssd1 vssd1 vccd1 vccd1 _1865_/A sky130_fd_sc_hd__inv_2
X_1787_ _1788_/A _1788_/B vssd1 vssd1 vccd1 vccd1 _1813_/B sky130_fd_sc_hd__and2_1
X_2408_ _2408_/A _2408_/B vssd1 vssd1 vccd1 vccd1 _2409_/B sky130_fd_sc_hd__nor2_1
X_3030__124 vssd1 vssd1 vccd1 vccd1 _3030__124/HI io_oeb[27] sky130_fd_sc_hd__conb_1
X_2339_ _2402_/A _2558_/A _2336_/Y _2338_/X vssd1 vssd1 vccd1 vccd1 _2340_/B sky130_fd_sc_hd__a211o_1
XFILLER_57_479 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_37_192 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_13_505 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_52_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_13_527 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_346 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_21_593 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_20_85 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_0_453 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA_input32_A la_data_in[38] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_0_475 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_497 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_29_50 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_63_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_321 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_16_365 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_43_173 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_8_531 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1710_ _1711_/A _1711_/B _1711_/C vssd1 vssd1 vccd1 vccd1 _1753_/A sky130_fd_sc_hd__o21ai_4
X_2690_ _2690_/A _2770_/B vssd1 vssd1 vccd1 vccd1 _2705_/A sky130_fd_sc_hd__xnor2_2
X_1641_ _1641_/A _1641_/B vssd1 vssd1 vccd1 vccd1 _1643_/C sky130_fd_sc_hd__xnor2_1
XFILLER_6_43 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1572_ _1616_/A _1616_/B vssd1 vssd1 vccd1 vccd1 _1614_/B sky130_fd_sc_hd__xnor2_1
X_3014__108 vssd1 vssd1 vccd1 vccd1 _3014__108/HI io_oeb[11] sky130_fd_sc_hd__conb_1
XTAP_302 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_313 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_324 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_335 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_346 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_357 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_368 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_379 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_2124_ _2125_/A _2125_/B vssd1 vssd1 vccd1 vccd1 _2124_/Y sky130_fd_sc_hd__nand2_1
XFILLER_39_457 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_39_468 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XPHY_19 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2055_ _2112_/B _2055_/B vssd1 vssd1 vccd1 vccd1 _2064_/B sky130_fd_sc_hd__xor2_1
XFILLER_10_508 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_335 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_22_357 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_195 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_2957_ _2958_/A _2958_/B _2901_/B _2901_/A vssd1 vssd1 vccd1 vccd1 _2957_/X sky130_fd_sc_hd__a2bb2o_1
X_1908_ _1908_/A _2006_/A _1908_/C vssd1 vssd1 vccd1 vccd1 _1963_/A sky130_fd_sc_hd__nand3_2
X_2888_ _2888_/A _2888_/B vssd1 vssd1 vccd1 vccd1 _2908_/A sky130_fd_sc_hd__xnor2_1
X_1839_ _1839_/A _1839_/B vssd1 vssd1 vccd1 vccd1 _1839_/Y sky130_fd_sc_hd__nor2_1
XFILLER_57_243 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_405 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_151 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_313 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_306 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_13_368 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_143 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_9_328 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_31_62 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
Xoutput73 _2062_/Y vssd1 vssd1 vccd1 vccd1 la_data_out[72] sky130_fd_sc_hd__buf_2
Xoutput84 _2801_/Y vssd1 vssd1 vccd1 vccd1 la_data_out[83] sky130_fd_sc_hd__buf_2
Xoutput95 _1750_/Y vssd1 vssd1 vccd1 vccd1 la_data_out[94] sky130_fd_sc_hd__buf_2
XFILLER_16_184 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_121 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2811_ _2919_/A _2927_/A _2811_/C vssd1 vssd1 vccd1 vccd1 _2812_/B sky130_fd_sc_hd__and3_1
XFILLER_12_390 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2742_ _2740_/X _2609_/X _2741_/X vssd1 vssd1 vccd1 vccd1 _2745_/C sky130_fd_sc_hd__a21oi_1
X_2673_ _2672_/X _2652_/X _2653_/A vssd1 vssd1 vccd1 vccd1 _2715_/A sky130_fd_sc_hd__a21oi_2
X_1624_ _2468_/Y _2965_/B vssd1 vssd1 vccd1 vccd1 _1624_/Y sky130_fd_sc_hd__nor2_1
X_1555_ _2920_/A _1555_/B vssd1 vssd1 vccd1 vccd1 _1556_/B sky130_fd_sc_hd__nand2_1
XTAP_132 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_154 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_143 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_165 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
X_1486_ _2898_/A _3001_/B _3001_/X _1485_/X vssd1 vssd1 vccd1 vccd1 _1487_/B sky130_fd_sc_hd__o211ai_4
XTAP_198 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_187 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_176 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__2350__A1_N _1859_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_39_276 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2107_ _2107_/A _2107_/B vssd1 vssd1 vccd1 vccd1 _2164_/B sky130_fd_sc_hd__xnor2_1
XFILLER_27_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
X_2038_ _1888_/B _2037_/X _1988_/A _2273_/A vssd1 vssd1 vccd1 vccd1 _2039_/B sky130_fd_sc_hd__a22o_1
X_3142__236 vssd1 vssd1 vccd1 vccd1 _3142__236/HI la_data_out[61] sky130_fd_sc_hd__conb_1
XFILLER_50_474 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_10_316 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_10_327 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__1518__A _2939_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_3036__130 vssd1 vssd1 vccd1 vccd1 _3036__130/HI io_oeb[33] sky130_fd_sc_hd__conb_1
XFILLER_58_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_58_585 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_18_416 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_449 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_268 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_60_205 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_9_125 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_9_147 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_9_169 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_364 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_3_55 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_3_77 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_1_592 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_49_541 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_64_555 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_441 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_290 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_32_463 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2725_ _2725_/A _2725_/B vssd1 vssd1 vccd1 vccd1 _2725_/X sky130_fd_sc_hd__or2_1
X_2656_ _2653_/X _2654_/Y _2605_/X _2585_/X vssd1 vssd1 vccd1 vccd1 _2657_/C sky130_fd_sc_hd__a211o_1
X_1607_ _1561_/A _1561_/B _1560_/A vssd1 vssd1 vccd1 vccd1 _1608_/B sky130_fd_sc_hd__a21oi_1
X_2587_ _2526_/X _2527_/Y _2585_/X _2586_/Y vssd1 vssd1 vccd1 vccd1 _2589_/B sky130_fd_sc_hd__a211oi_4
X_1538_ _2977_/A _1538_/B vssd1 vssd1 vccd1 vccd1 _1544_/A sky130_fd_sc_hd__and2_1
XFILLER_59_349 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_47_39 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_27_202 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_23_430 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_42_249 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_10_146 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_117 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_2_389 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_18_213 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_46_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_46_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_18_235 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_53_71 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2261__B _2261_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2510_ _2510_/A _2439_/B vssd1 vssd1 vccd1 vccd1 _2512_/A sky130_fd_sc_hd__or2b_1
X_2441_ _2450_/A _2450_/B _2451_/A vssd1 vssd1 vccd1 vccd1 _2442_/B sky130_fd_sc_hd__o21ba_1
XFILLER_5_183 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2372_ _2371_/A _2369_/X _2370_/A vssd1 vssd1 vccd1 vccd1 _2449_/A sky130_fd_sc_hd__a21oi_1
XFILLER_38_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_49_393 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_37_544 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_24_227 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_64_396 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_20_477 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2708_ _2568_/X _2496_/A _2774_/A _2404_/X vssd1 vssd1 vccd1 vccd1 _2710_/A sky130_fd_sc_hd__a22o_1
X_2639_ _2674_/A _2639_/B vssd1 vssd1 vccd1 vccd1 _2640_/C sky130_fd_sc_hd__xor2_1
XFILLER_58_27 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__2688__A2 _2684_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_59_135 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_28_533 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_3148__242 vssd1 vssd1 vccd1 vccd1 _3148__242/HI la_data_out[99] sky130_fd_sc_hd__conb_1
XFILLER_7_437 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA_input62_A la_data_in[7] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_709 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_511 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_67 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2990_ _2988_/X _2920_/B _2985_/B _2989_/X vssd1 vssd1 vccd1 vccd1 _2991_/B sky130_fd_sc_hd__o31a_1
X_1941_ _2036_/B _2036_/A vssd1 vssd1 vccd1 vccd1 _1942_/A sky130_fd_sc_hd__and2b_1
XFILLER_42_580 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1872_ _1876_/A _1876_/B vssd1 vssd1 vccd1 vccd1 _1873_/B sky130_fd_sc_hd__xor2_2
XFILLER_9_98 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XANTENNA__1616__A _1616_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2424_ _2493_/A _2494_/B vssd1 vssd1 vccd1 vccd1 _2425_/C sky130_fd_sc_hd__xnor2_2
X_2355_ _2354_/A _2354_/B _2354_/C vssd1 vssd1 vccd1 vccd1 _2355_/Y sky130_fd_sc_hd__a21oi_1
XFILLER_57_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2286_ _2361_/A _2361_/B vssd1 vssd1 vccd1 vccd1 _2288_/A sky130_fd_sc_hd__xnor2_1
XANTENNA__2447__A _2447_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_49_190 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_52_300 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_547 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_44_29 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XFILLER_40_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_55_160 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_28_363 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_558 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_43_344 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_31_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_43_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_399 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_7_234 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_7_289 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_50_83 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XTAP_506 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_517 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_528 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_539 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_617 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2140_ _2083_/A _2083_/B _2187_/A vssd1 vssd1 vccd1 vccd1 _2141_/B sky130_fd_sc_hd__a21o_1
XFILLER_38_105 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2071_ _2071_/A vssd1 vssd1 vccd1 vccd1 _2559_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_38_149 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_34_311 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_46_171 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_22_517 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_22_528 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2973_ _2973_/A _2973_/B vssd1 vssd1 vccd1 vccd1 _2973_/Y sky130_fd_sc_hd__nand2_2
X_1924_ _1924_/A _1926_/A vssd1 vssd1 vccd1 vccd1 _1924_/X sky130_fd_sc_hd__and2_1
X_1855_ _1791_/A _1979_/A _1852_/X _1854_/Y vssd1 vssd1 vccd1 vccd1 _1856_/A sky130_fd_sc_hd__a211o_1
X_1786_ _1786_/A vssd1 vssd1 vccd1 vccd1 _1788_/B sky130_fd_sc_hd__inv_2
XANTENNA__2760__A1 _2141_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2407_ _1888_/B _2684_/A _2483_/A _2273_/X vssd1 vssd1 vccd1 vccd1 _2408_/B sky130_fd_sc_hd__a22o_1
X_2338_ _2567_/A _2411_/A _2560_/A _2021_/A vssd1 vssd1 vccd1 vccd1 _2338_/X sky130_fd_sc_hd__a22o_1
XFILLER_29_127 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2269_ _2269_/A _2269_/B vssd1 vssd1 vccd1 vccd1 _2271_/B sky130_fd_sc_hd__xnor2_2
XFILLER_29_138 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_52_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_25_355 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_25_366 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_40_358 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_21_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_4_248 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2751__A1 _2557_/X vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA_input25_A la_data_in[31] vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XANTENNA__2087__A _2129_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_63_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_35_119 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_16_333 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_28_182 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_44_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_43_152 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_45_61 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_16_377 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XANTENNA__2534__B _2629_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_12_561 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
X_1640_ _1640_/A _1640_/B vssd1 vssd1 vccd1 vccd1 _1641_/B sky130_fd_sc_hd__xor2_1
XFILLER_8_565 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1571_ _1571_/A _1571_/B vssd1 vssd1 vccd1 vccd1 _1616_/B sky130_fd_sc_hd__xnor2_4
XFILLER_6_66 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_6_99 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_3053__147 vssd1 vssd1 vccd1 vccd1 _3053__147/HI io_out[13] sky130_fd_sc_hd__conb_1
XFILLER_3_281 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XTAP_303 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_314 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_325 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_336 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_347 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_358 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_20_3 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XTAP_369 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__1613__B _1613_/B vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_2123_ _2123_/A _2123_/B vssd1 vssd1 vccd1 vccd1 _2123_/Y sky130_fd_sc_hd__xnor2_1
XFILLER_39_436 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2054_ _2112_/A _2066_/B vssd1 vssd1 vccd1 vccd1 _2055_/B sky130_fd_sc_hd__nand2_1
XFILLER_35_620 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XANTENNA__2725__A _2725_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XFILLER_34_174 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_22_347 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_2956_ _2956_/A vssd1 vssd1 vccd1 vccd1 _2958_/A sky130_fd_sc_hd__inv_2
X_2887_ _2945_/B _2887_/B vssd1 vssd1 vccd1 vccd1 _2888_/B sky130_fd_sc_hd__xnor2_1
X_1907_ _2008_/A _1905_/B _1905_/C vssd1 vssd1 vccd1 vccd1 _1908_/C sky130_fd_sc_hd__a21o_1
XFILLER_30_391 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
X_1838_ _1981_/A vssd1 vssd1 vccd1 vccd1 _2329_/A sky130_fd_sc_hd__buf_2
XANTENNA__2580__A1_N _1859_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
X_1769_ _1821_/A vssd1 vssd1 vccd1 vccd1 _2313_/S sky130_fd_sc_hd__clkbuf_2
XFILLER_1_218 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_1_229 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_57_255 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_17_108 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_45_417 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_45_439 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_25_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_8
XFILLER_41_612 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_40_111 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_9_318 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_21_380 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_5_557 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_3
XANTENNA__2724__A1 _2725_/A vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
Xoutput74 _2123_/Y vssd1 vssd1 vccd1 vccd1 la_data_out[73] sky130_fd_sc_hd__buf_2
Xoutput85 _2856_/X vssd1 vssd1 vccd1 vccd1 la_data_out[84] sky130_fd_sc_hd__buf_2
Xoutput96 _1764_/Y vssd1 vssd1 vccd1 vccd1 la_data_out[95] sky130_fd_sc_hd__buf_2
XFILLER_0_251 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_1
XFILLER_0_284 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_56_93 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__fill_2
XFILLER_16_141 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_6
XFILLER_32_601 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
XFILLER_31_177 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2810_ _2810_/A vssd1 vssd1 vccd1 vccd1 _2927_/A sky130_fd_sc_hd__clkbuf_2
XFILLER_31_188 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
X_2741_ _2394_/X _2549_/X _2550_/X _2814_/A vssd1 vssd1 vccd1 vccd1 _2741_/X sky130_fd_sc_hd__a22o_1
XFILLER_8_373 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_340 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_4
XFILLER_8_384 vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__decap_12
X_2672_ _2642_/B _2642_/C _2642_/A vssd1 vssd1 vccd1 vccd1 _2672_/X sky130_fd_sc_hd__a21o_1
X_1623_ _1623_/A vssd1 vssd1 vccd1 vccd1 _1697_/A sky130_fd_sc_hd__clkbuf_2
X_1554_ _1554_/A _1590_/B vssd1 vssd1 vccd1 vccd1 _1588_/B sky130_fd_sc_hd__xnor2_4
X_1485_ _2950_/A _2892_/Y _2950_/B vssd1 vssd1 vccd1 vccd1 _1485_/X sky130_fd_sc_hd__a21o_1
XANTENNA__1624__A _2468_/Y vssd1 vssd1 vccd1 vccd1 sky130_fd_sc_hd__diode_2
XTAP_133 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_155 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_144 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_166 vssd1 vccd1 sky130_fd_sc_hd__tapvpwrvgnd_1
.ends

